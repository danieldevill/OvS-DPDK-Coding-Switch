// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:04 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Tbp2twWWBCe+ClQOwuhbJuNOyJXbAEJjErbLnEqKs9ww8NWpOWKUxyh13Um/gkXL
e6zgl3EA1hJPWVcI6W06XYCJLpN76X7FOhppxUb5zt6nKp8UpT7bmNzMeT8SoyKf
D4ewQw5HRrZiSyJIJHix+S5HROARdaw6wsXIFaaMXcE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18000)
7bnFe2+YsoXilDSC+7tJSNZ6uuCHgl3TjuP1FIKo/wXILqtnDi9fI2Sr+c77P0Jo
zaoKQjXDaBy3kJYXX43mh+/9rx5dOnZq9fYtbZvzVUjKCOjv4R0KuYPoPLIIOZPy
+3kpyTwmaJcDuh3XI5SiZ4PDeQOWYsYkInBxyF/IhFn5ZICE0iwrt2gbupeVPfBt
jqKCoVqKlcsxedCDRFwHSxt0lzc9WZRD7tAnSKdYik7LppdeZwextVVe9SmDBJRA
BUEnK50v0e7ZO+B7AGMbAJcKS09yfCyhjN7NqulAdya+rqFs6tBVsnNA9J1/BmV0
sePSWkZ3KJ4MYB+taUuU0OB+gq99/6IXu48LUnGqTRq0E5/K8MniiTcpKxQEyGCr
yiUS/Hg1YnHrw7ak5cF/SW16X7ojAhO8PfyvVb2xInnQ2AOHyzmomYux2Mn+r7rB
rZP9mvBRqUtpcJoiQW+9056IKqG3r94centnz4I9tdRUY4RLuZfHeAXciGS7MBbZ
iuiwbyYUDrrODUg0c6A7eMdZXPoVMItnAg/GrQHlbEwmlMtx3kXlrwVi7BHq1EGo
3Y4EUWXuvRzGwe8/Qu2NqrUN6hAtiZ+1xslmuOd64bAjNaHmcVy5LxaRXkhXMhA1
hy0kmdH6XBsKAX4MKApfWcf3l3zCHnkLxpQ4/obiAEwt9AuDxG4w/Jk+eSExjbV6
bEMJL1GaSurKzHlSfUVQFjawljfMQsiNvBg6605qs+7k1MiAHOvps8w60ekBkjfq
yW9TGdNPYS0cdEyiBy0WFGKTypoFjbsVvPTfQ4lazDlr6XqJjSpcRG1GKvWSSnf9
+xjTbZq+aeHyh2lEmnV+Volv2xs3tvpY9SV9FhMauouPuwh3fBUcV0TnQ5K7kgBk
JWk5IsosTIbg+ZwEYlesapXxnxMz2NUgPIUWe0ixk3tgSSJE0YJjvZkZYhuY5Avo
T/ccoKKElyxZXHuL4+/UsJk32kf0ncvW8hgGiqvT1ey9pwOsAzzKn3FLDJRkb3HL
/d4+JLjlMY/SBUPisQDkDjovufNbFgPV31Wgh6a5uJCTjgSyYLUUdy0pKINR41zQ
F9O5xQURZvLnr4PPgiDBII5aWvULXOUr+8X/BQnqh4o7wegTEMgrXI6PU53Au4sm
WXpmMBvkGEuiee7NLsczOLu3QKv6OS4wtBsbEEENmrrNo4pEc2pPkmHpz8F0Sc6s
4cF4h1lGOJ3v2gizpbARuF4zjqmenHK/JV2y2x6uYJtYTSsxjGuFkMd9xv4ss3H/
hSjVvoZR//NMq5ksRjuv0459obIKhmNeeNFXynaH74yRJcv9vhiNKG/XuMcslHmm
gY0pl2VrEK49ZJPoL8JZ82B6eBcI19PXt4gq3NbOqaktygCNzsSPkesiKs3hNkaT
wQRv5P5BvpT7LJ+7cg9rMfGOg0DDlZ0xSbwbKWkGWws/RW1ojpsBp8x1ipGlZhru
EyO+xabj2xu8wsvDi69/l6mEIQCgR25f+5Coya6bzTayBPzUDGHGx2m8P/LUv6R4
6uxX9q7d1pa5sziiQMAF0pPGb/Pj/VbnRpFE1GSvY8ql0wCypvcCPHohSUJ3xQjB
Gj5zrb13d1dqYuBrZGgWMQdWY9RS56BTK0ey72O8CfEoJ7xfzLlESlcgLc2ng7GL
plPPEEZNyS3cRDWQtsejUBHPRhtrfcLzSnUosupmBkF9mF0TCtk5aa3eNdhOFxB5
tURnvJwgcJ4avCAtpPHT3yZqL0txSMmQJ1guxAqecvag6M5yxRhuBH7AjnR2jhIM
Fddw245ndp4kIS0NrI7JJW1/bsypM1BCSB+Iz/Nh40aLNE4+GA/u3t+iSFV+imQR
T6ZMQCCFfoAQSBn9TeGfz1nz298WK+FAqXAhtbfwLwykSczr4J63rEqQj/ZDhOyb
G3qmXLK6AdkvCgdUjz43hswGhWlQsK2qMcERQlJ0v3WF7z+Shss+cHjTeBr2Y16X
SXrgJIlWIDDBkoICt6ZOEm8HezJS8Jy3cfcRUiPzJpieWBYqbDcET4OhOcETx8kj
JlD3Jyvt43RxvLOqSXItqbFq42FlqvGZp29O5qCfz8JrRDEpiNq4yRPNLDw0onOa
DBThyU8SaLLj/rH+vD+RsYioDP1/a5cLxC5w72i+YMNWtSSvf06da6aiOT5Hpxcd
BolFEXZw/pkO6ewdz6IEiGAtYwv0s8OBzFyGBmDYmXo6uZW2Y5rkWty/OIUIALOD
EXg40YKviVfRvkOA00+HJWbeyZBS9Xbax3jTVSjYO/xIgSJyD16H6O0uU5ZBO72E
5HkaP0c+cJgKsGZWg4VrMz8iM+JQqTMbILhi8KDaX728otCxP2asfbas5QNMUpic
gbCZX8r8R2oFEtne3P2eKfHFWevaWQ9mzNJMx2/g8D0cbxkFl5CB1iLzTCmI3gLT
0CInjAPRMyWqicVIZBNskcs/fRAR8u5FcWZ4EZdfeFVL3LeqTDiWUY9eYhIOmnL4
Fx87ayVPQV8hx0BgvJsBCjLLVwBsaYP1pueJz87vyQ9VzSZli/etrb3Tapelw8/5
ijm5qM+1WsGwSU8DksG2yEMfpqKfC365Q/BzEAs4AcVNrUXOx30XDQGAwoNkchrt
UGhdryaKjWVvxG3tV1+Id+GwZQcajZ0b53XrDlq/5kFscizNjgq60rod80abNsej
Npp8rJQfFWYQWW7lz+LKWVLP1SYq8h6WQVkMe8rSV01dn+kHJd4+cRhn/RIpapay
xRvNwwMHsobZrVocqDWePxSTkg+v1yGpbnvLfU51bgqOlAl93h1BeQVhWZGy7N9S
j476D5u2yf5Xa9nsvT0qzkiaUW/Bs258+8/Ie551JD3NZZAsVQ8c10ImEFy4LVQ0
EFzBqAdBRzalb7HpYaMDkqt6VACXYmbg3pqUPGWoBynTiq+VDssPsFrm/qga2b2Q
F9+/17z3sNJYm2/hxsMsDqlYZ0hshMK29jkPa4zmA2cI2izci4iZA1JT0oZZfixD
Z1h1/LjCfw/eTVsEg3bD49vC1sPg8ZJHMSk5k93dHE161sfoJ+FyAF6n9llZIlbA
pMKLE6FuMMGxBDBHJlgKu7UTYNxqEO+r4+c+i18W2nkl68ce8vyA8P3+bRrucF5T
1ovRby9tPyK+RTftHBFw+9HLhvtb1EJ40egN+cDBJd//R+kVY6XfX3G+claTnSoM
/L5au0ldNufXDu0Uwrr2Mg5+L0N9gUEpftoYMD4bH6PArZsUt6MZL2zYmrGpRb74
qJzJ581YSOhyu2U+UxqCajI9Vxu5QddpDs3TrnexOoywAfnhPf6WztZn9r2y6KB2
0wiC/XfhZyyn2UKXkMAW7VPb9DmxCqhizukpYcUU1vOpDMDA/o1yA8htms0QJOeM
ZILpC6fcKYWJNv4kjRXARlmou9x0GCzhAi66mxyfDLZNHHrmVFkCJ9JmT+O99dut
kbVg8lUaHe6ot+SgsmjKG2qvNjEd0V2DhPIHaCdd5bz3m7GJZhQh7ftt0qYz/LEU
YvbP9rfwzofrYlCqxG1MFxrgEx+KtA5Y+3jRfIJrGYbcOXetU0HaAvhIKg2xPBEa
l8p6V90dI2OMxQKwejO0CqaZFBeCvDV0Qca35lBu6tfBkCjDh07Pi9HJasux51HB
+FzpMv4KzA42lRdwD9zv4H0O6PRzjMtx377wcAQliwVz7d+9vAQ8qpLY5PVOmemI
iq/8/Nq+HnWiwdD/vZ+B3caBnrMR0GndA+n+hu1C/AzJ8QF6eA4oqmfaMWBP9rUX
uO5t3ukuiqewTtJG3kA9CthaCd5pE1BqDy3hJ1LMX3ST1Jf81ZGwhZtSMCuVn+av
Mnuv4bNrbFDBK68cG86IAKn65k67UtW23dJoIVfK1m4ZFC3HPHBvV6l7pjbPJTWP
HwHvC3buutv/bHSQLUFC9VxsPAeaUlZxy5SFVbZitYEYfS5EiCrzCyQ7jaG4ChUi
oKaSXsZNgVapDIsbAqDMnuKTm3Xs3zbByqTmmi7fdU3DYkAXkEiWgkf87wb3XnL/
lypnzYT88kpLTnlWQfYL1476pqqzFhvwx45CIH9X8cRK1B3tQSr277siPtDga6qp
576TLWSJXFzQrSVM7ky6BnczeauMsGfcDrY1uDOHZuLsmcNJEFemhoPELShoa9pk
F1d4rthLA5nYqmwAItElujm56H988GWaEoWYeJOPdZ/oI0R1mT31IwwPrQrVWA8a
VvTqvxLt79YHoWiAtLzFoNGf4I+DgQjVod8dVucrtOp2/CoNA5dc0yKmj0G1n7rm
ocQXRnyXNuTSHrruamt+1Edwj5pZVxpIaHLVAQSEPtms70DsPalAGTd28X++z/zN
hfXFspsOgzeM5fXM8aZMN+AFuhe8nqNcHWKdjY/O+zoOnsCNRJh2abljWuLPK5SJ
OAQsvJUYrRZXAKoULFxldVlC9wz/0xwTvXQ8FWOUhBkj0+nV9em819K0oht4Eeka
YFzv8Q1bdkPUoH7IGaXRCObsqwMIyPiNm5ubKr53QOYJ7mLlluNXrVu2OcZiSXU8
lSoF3XKVIEzwUknUT2R8VC99EGkGJMndVJytLu550vexCQGiseNBIzi95WA2ffmw
MhJLjv6z8hy8tVYeVFsk6XFBgzGiVfjnxr0BIKgtvj+eSjX1BHvEd+HhZsSCIeSU
RTU37jVJN64Q8UvwE6uFhZYQedjwfBGW8FgJh08nJqOSM7rOQTiWy3VjogeuemMa
yyh+ZhuCx2/kuPOOPOKKIvxgYHahyjt9ijnkAnYBCrvbNErnwlpGoKMkeJkhmLvb
Nf4jYTp/WMpRpZYhTGzZp7T/4oX3PPbJLHO4M+BW0H3p3RC0pRX/prhfR5iK5fXC
5jZKMGHVB+XdQ3Il6kcJ7rhuMbeiT9J5znDHpvO+SzT/AtMR2Qh0wJNoAx9BT2B2
L27SjOb4Cij5BdiUEn44G9FZctnMTME+C1iq67Cv5HQ3K8C5ZXHoL0YWESaGqcJH
3xw3qp4NEhOgXarhngZRBMLhH3PTseTwLPJA6L95GY37x5lfvoJ8oOWTJG4C8xXa
oPfDH6oUOs38dXHhhBbiMPtJS+tAPAb94g/Ra4Gl/jncUpsfs9/Tm6wd683WrBNU
QdWJQymVjGZR4uI0GylT8DTc1Fu+drSo2GwvxJzalGvrGTyUdM2B+vC68lDMuvfN
HV0OP3DIN6hWbFHmSIS/ErMWDzJl7Bfnzal0ajdW3M0XmKuTlx+OagSP98A1wKIW
Aq35HwmaEGelPWliVgj74mvOXa3IBO67oBQ+O1Lm+hCXwIpXTz3bD6xn/JhFe7Rb
rTmFsF69aWBZYaf/4N+M9qD+fVMTd2fJzK35YDHyiqu2J+msnfZbrqSr0dqbqdmB
nIHj5cwrQ/znYjQ4wBAkboftxFvsb1E296xe68jdUXu3MdPWDJP1qC5DVp2yf9M5
2w2+hT4At6lU7qs2xEeL/uCR1v6vJlsqY0ALZcBBy3hLQmsNl8Rx2oBdqNBo0x8G
qvh2YUtYgRkqczOwGa43fHrdWSZ3e/LD0QnSNxeL1RZhU4IclUc4wWA1feZ438sX
9J8U0Z6bXKcaOOVP9hm83RgTd9wwAMwgwR9FK+FmlEGtJUvQ7DMH1ThcFfTcUuMt
za7a8WW17f8Dw6f5Vtzcq2gvZDN776kgyBzlMFTAtUqVAHSMvy+E6m+WGfkR3kmI
EBTR1oTFASMqH4K1AFH+lvho4QKy82ytaADYAI/Ms68hPsgpjTlEudKK7zdfvR8G
Dk7l+yn95YzNzbiArS4JvaY5JWQw8vpMS0DKPgU3ic+loaJ5UT8PHLDmEoRUHxIm
5QC6GtL+N+yOu850BWfIEEat3ra+c3WpRZmo0gIlIaGcWJ1iYhKgFq6hQ8AFx0gO
B8nFLidN6stT+45tEzLN+iqTCr8nSpFJddChuPVPJKDd5L14FUClEIO69rh10cc0
IOGAvIRo5f3I44JmuiRkp/7JNpl93mmA0Rr8uGpa8ADUG08ZNobBFqXMbc6c+fNA
x8Bp8CUMKugDPog3EhBCZpTkNHV3XxlYsv3avvmfrb8mP8EWDtk4aF+YFM0gU0kd
0pjiw5NGt22LEQYU88VrKRSHAlkueiVKLf2P+X2O3iBtG/EGMFvztSTZGc9LUZ+z
NF+XrmsKy9xbC/um22sZWtDTii8HCqTgaGkeSo+U9hoooyoo5Ak8KuaVZ1WVV6wO
vv4s8tRelugRfWb8RVdnhKzzu+aLGYg39fzi6851zWnjxhbXvuJm2NG03G3KHGYo
xkxytu//HhrHndywjVvKEAO9C2ctxUgcTah+ttVnbKwDyBBxuimYnVHbDKeJ8+YJ
e1WAmWWBmEVDfOFFrr+ikTw8trVDADdI1CVdci2KyE7oDyUPUwmcNqE7C8vy8Pah
7+lsML/ciWatnRlU0TTfquFimfKkE744iK6r4bzKzv0hJSiI9acvo1WaBTKCKC8W
RklAz3lvdhJcgCz19PujLL2RK67lt6i6Bs3PWd2PRy55KW4Pfm+fSzVOnBMVNa7A
wKPNJq6t/QH3q7EJ2K3C6YgM7LTf+sgLiDz4wCn5/dNRbRRDjlq/PQGhJxdWLw8d
CZba/XIiGOwh3IX61BvtBnJ7YIjtXBm7ZLieo4EAfHX6M+a9sT5EJ9NooMp+VPrs
nZpFyA3/pyYDnS9rhG+Sa+fyYt2iiK+rL7Stv9986+izOeqNPAGYGcN7udpZFL9C
nRbDlaPHQKqG4FE0GuOsvZ2valD0dZwsZBRsoNgEkvxCOTmFlwXzlqTTjqOue6FP
f5CkG5QPDEDMES3FuOFUFCxK3v+0IeWq/e2kW4dicrAcjqm+4EnamfDpxm+tZJbe
GGbnW5ydpP0ZTNTY03fXKFR1qHAVm+++gWNh0XOJNRzH6DA7peoV5ZCeb1jJEx6s
tU1EOxp9ushl+UOH++iSqm0Gt1WvkwLe9PSqUlCSLlaDfAThfvpfMo3KAI3wRBkJ
hpuBecQs0jJpdcdL7n5EN5hRuArxWwRxo5CO2GW63b5BSj1Tz/YP+HVFSNIXbu40
K7kkFTdJdj77opJR7DU78gvL0TCPW1K8UJeD6nkrQAd5rXXEqaeAzSOXIWeEHEMj
AaAWnDMvYs/ChXaAD57lqC1USWyCh8A2cqfP7NmMEJMg+8GWdcmIANyqDupPBA0E
12lAzsnyY6w+S1lb1wRYrQ/YkSHLEH+x5MlaBuJtSkCrGClpoZVnSCzIV2YIsRkb
oVnFWAMLI7oMWxLRL5rzn71qaV5PWC/4Vgy+SQ2AZOwEnMekxlMHQBh542EDmDxz
A9BvEWPAupTztJf6OXWEIrSt0TYmo284FsJf65dxQv1xIXdID4gGeXwlBs54QoqD
LGBBOg2AYuEhRvdCbMUMM2TwuumQ9xpI1Kyaif2QBwPUlywNfmeHNzEjFtgSpws1
Q92Tt+Q6MgOOnbZaCeiwV7n3Myn4+1nHmamnm2Yqny+dEffdENcmfb+ewovoqwZ+
GQmts8Ilq+3xdvpdV7jLfPM1N2FK33C0zZYTklRtEHNqxoSnW7P1gM6h525mALRj
owoJW3880gtYbh9sjjsmsxEFBRHId53V0Ua4SEIMFjIzUNStjPSlKbv2gAGh8uum
PhAPPr2MBtyUe20zcy+JhORy/1COnEdn8Y2Xd/Nu+kFDVlGLavgK7JztkpomYA9j
Gzkw0PvCEqGC/yZZxxz1p+/DR2LY2EeO9GCpkGf7FJ+5bBdfzkxNhTt261S+hM9J
hu3eC0vh7QHZXoMHAEHJczDGZDGPE+HfCMHenvo3mGY8Tkrfs10i6mXfphxyQTyB
q2YfZAJNsyajzFQbqgSYrUDHx3J39uBEHdKXG/KJclptD1BY7X2BdsqcxxsPraSS
RWXm0//LMvO3hXh2Z2sgDjIL1yYLyRPSAWZyI1DgcZiRN3YCrGeh5FbLLKyCRtu9
HhMmDv1QBO1s9RyZysTHRL6TIcn5budcJbrwm5hXXJWCpPX4XTFpdWHFI7h1xWI+
OaYuwfNtiOrCZ/0A1SsVSSofon9bB3A95z5DUUgKA4q6B+AucMi26neAW+8OFXyz
5rYcTZAIe4otdQTxpFxQgsVgiwDjshP99o4Z6eXoItJt+IMT7jyQIa8mfxov8Khr
lm8U3GZ2ufuW4vZEnCE24TnoFKP+yIu0gg0+oSDABMxuEN4H4StRsriQ0m3ZIWWz
rqS6tDRDaJPW/DCaQE6GHkb9rFng6W7MhnoL4KwG1Js2N4Rxc4mp4SbRW9wY2+6H
qXDqb0DhP7u52xCZ/+/AoZdZFZkaPNLMxnV9pzLkUoHhYGIIvoZ4X/AQ8awbv0O0
NdmxM4zPJshmwIR0kJR9QRRKgFOZ7BFG/RoKw9BOvDzi7hYfUmW6sW/xM+tWnPVj
a4BQTEjSMfQRmnAJmF68Agdqv0AlComY//5I05ebdxrLG+mML02ZuRxUzPy3lAtG
LL8/zD2+E+yvDrrgPKrEyj0IsXfwEooOXXOAyFDsLJ08cW32JX5SAdUN2HV0VVVw
OXhNu6SU+8fh2v+py+vbrue/i6NwuN8qlGvoSJzSykLDsw3cpbSXhWAVckOr4/mX
nF7u8osieRsJ+Wc5y7zUSo4EYp2b+e/wPeFS+OAVTwzsxSzYLcu800ZSIY6e9Z8t
Bw3c+GHNxKIiOLo88nLbJcCQoS8wbh4DN0f1uqTLsdtTfDVIH9UfWRftQkK90B78
m9kgQx2LHYpryT3Klbk5kj0RvBIzOasC8pJt5A1EiUSGk2glUOSxpZstPswN0yNX
+1hUbyX9f+7rvqX52PtaThgJ0xX5/RuxnDk4G6EAQqHR1Rcs6m5u3VrjauiNuCFG
1XKx/dWmzAcNR+qI2SbV5+rbsnWrfahkdRQWBzzJXbWNI3Nl7HQt5rzHYVYzMlRo
0fHIPx8U3yfkZ2zx6nVsyQNQiyltZF33VYhzeaytuQ099Y0WQR119jZmOzUcm91t
GIq19iYaLYbJoQiEHWQxzG+YX0foi/fCfWeO7kdR6yBUlkSdYpQUv9GQTMNmLgbC
tb0wXyw0xFm2L7r8Oq5Yv5lwl1ifOu9xdk8AJjeI5QLHLxsBXGIreKfHsLH7CI+G
1r2oWhnq0r4by7Yzi7DsxJXta7V/1oBylghs2wLkC09VuxHGAsBOWrQTRHiIERCn
ssw62+Ry8xMZGO2QKZJUU0qShinnfJIbY9LUFXpxEQZsAjop2HxYMkn+0FNrswij
omDsJWzFu6vAespbOhCArolg46zmLz04wcj13HYfxAvn9uKMtqN0qdvbD5otjWlO
ezYKxkGyywW5sZh9LRWC7rcTj5rtc3mkQ8cy1RSGcscS+dlCtEv2aVNVMS/M6vHO
3NrhxmksHqhJrPBUAhZg2nM9Vq7g1M+zzIV+9nxAGK/G0ufhIvFvNza7UFj7WR2Z
MwryVE075mqBJB1ikncS7YHBvUe1jCttdwRS/QuvC/Yph5jcNFqhC1tViLl/P1V6
DUT0Fbv9vcJnjx2/tjvYkPjthmYmxB0SsNmPbseIxu2vjtBjU86c4YDr066tTSx6
8O6LUbC4ExzKhCgtENUYk11PZPPIST1w4gKVKS6uTCEqoZ4bwXDWhJwVTfTZlJS+
8n+xoi/crhmqyhosu1lT4d/vE4kdShTUkCFdKNw7WZcbLRP3dE1z+Xj0aqgthTPJ
vUMmLvKU53rXVGEsydF2YTFPSVkKBrLmO3QG47H95+zWXB+TtMEi2SzyaG8Cnayy
Fm9lJRdKC0PoI8PSeuxOpNee89MAL8IRoP5yJ/OSctY2d1dWaBvVPMrynBadUPBo
v0fV3KTbSKirP0x0jIuO3OZa59t9DtGWW3CSoKYgUCwvgBo66dW+8gRAI1TpXJG4
9EmR51i2iempihF3PXitQ8mnC5UedfVd3JoJsc3s6CvjGDwBpuFjpBN3zgQGcC5w
XmhcWDyhwyzFEY3zOA6aqfaCHsJphMbk/tr8AclIewG/J89Hey7TV9rzZ0/HDc3t
9RHkEC/60vgOhWmFW5YwtCuZBS5/O4d9KAf9+SDvVauQek2Iv8RIAO+5zX4cL1qZ
+PmtWUu32h30biY6WjhSt70P/w7R3Lc3IBnDYvOp6gYcAeTySYySDPfAcstz6Vs+
usLx2j0yGROsSHTV6spLiqqI9YjVwqkbTMUzg9VJe91gbGHzUEg2vHNNJCRanMeZ
wdchnv9bI5AwmN0eeAsoSOMZqQobVDSvzKJ8lrAfdie+yIb8EWaCy9E3zj6bemvv
lPw7qtkIwG11bSeJvFzTDOhUTlfgFagQbMz7HvVSyPa9Pc1XOg9hrvrw5jfdGKb4
Ch+6FcrYkM6CYapIGAlaWplGxOo49cqB+Zhz1V9Iilf+5/91FHdI0EuzxNI43pof
ZraySXmZkUXtmE7RLR5Y8a0wmFIKlqgFOAegGFgYsCmBwAot7Rf/eN3p4mRtQ0ko
v7C9UbP7uHbDIQqn6NYfQ8qBqQClRF3ltE7AzLj9bjMKIlcWAUcpTW4N8htJiqUw
ap8oDBdsZupO9E/GudbU5xEvrLfWVO9wAPqlIbqKkYo3zwxZ+6wn9Z8Ih25DyhWh
VOfhXAj/rwzvnIBkYDWr/GYCWjJLB8rm2gwgS+YPD2Br6c8a7w21O6lhN/ZIcJ8O
TDr2pQVdY2t2xxby/0F6MozA9iiVehqxrZNSp48FkgfIqEg2eRO/EIpbZ6z9svYk
ixwyrRHC5kATK1YgareoZHSK/tZ6+XdOiD6hs8GBR2YBZaS7DDpn98aqO2yv/q3Q
mjvejkyPQel+aaWtvjL+MPInJKX2sq1hSi2kGwsw+eXIB+rh5p69oNR6le7eOZ6l
Txj0YWdqz6Vop04dPi1MOQ+jeloOOydvpacT6y4XmHQ6zplS/aA4XEdTZhcdd8jA
dZwtf8AhTeAemKBhTUOAilbH5QcJdSzOM+xyp7RMEnFKsrXA0/GozpIe/UngBfUb
GsgJ6wU3ZFCowvJjiNG7MgyhjL+nBsYOYPJplz98RJiLa5Pzm9erGAk6IVZEuYwX
iZMkvpw0lleTn6NjTqLslq06r5RwL3CK2tVEXXaZHhochZ2g/jQ0WmVA3BTIGPKy
cUmQ51hQPr+rcLETaxayG/vg6FiMfxu7/HK3pPZOdgFTmH/j5s628ZrGygVibjEi
IF06+LAzyVQeGUKfD+6nAbiUnHoKDE34V726V8h4RgJ7kd7W5RUB3IQbn6Z86QnA
xi12dlIwevpw9ZyomP1pG38aRbAejWao9WA7gQZg/K2oxpgjti9ZIE7HWDrETo/I
8vWuwe8pfFJARc3NWFWb9Z2oFVOHqScXB1n9FxHyN3Hi8cSP6jzIyl3lPdjx2gsZ
cihkQQN//1GAt1Wmw03DlaMyG7le3JC51aBeOA4MO+df0SX8twD6BEiX/B3eVLBL
sI0pls7RI520CkUOGQIv+DJYHgVSRj9veTxLswsgtV5Fmi1bLug9X1VmFrBRWwRW
4UQAkuz1wWup6p1jXxNzDYy9wTLYvokoMv6xAnS6ZIUsTjqEQZNFLHKYCqHFMOua
/xa1OhLBkiwvzIaZQsfOnoeYgbMPGqqfV0BPo/5CS+sAqgLNiihuXsEQ8sNR95O8
EsdsS0JbVREaCjfZVxTze0IhbJp/Ujokl+uUodoHYQone1VFKf4M3fwjU53QjVTw
8e1/4yVXxItqvuHXZcQyg6jjuVRSAg0EMR/X3z+PmLfjQk5PLPBKSHzOQt3ETI9l
t2OX8ICI1FAmEeu/XiSdjm0Mowc8rOvjWSoWaBVBEMD5c9CSFRwow0EKTS1irSST
DguclQL3LhTMRHMEJoKl/dxrr69ZysRB9xxZfBjUYYSMArT22m7ENYC7wMo4NZFt
wOQtnUF3kzhf62JdlyRCOEbzEpCAmx149RwFJQdstv16AjUjlZhdkZKPgMccvQEM
SgGMeTrsZG6G6Xtt1Zr6tYBJi3FFvMnbxarsu0vM6eezXtlzQGhMhWqwhhQWHoG9
Wo6qGsvv/bW5N3xxkbx44zRH/9CL6EaMznSmLAAZgNpk0eCHnsBk7niKO2j7l3pf
x0P4JB1GPcANURSOOhg5bC5Ceh959aUvUZr5Syzjws6VVA0shv/s5+0mkjhEJYPK
AJR6qj50Za3XyhHdZI8W4MR9PWdELtbHAMuK9ddV5y7vW0gbmZLlqhzJodM2BFu+
L/XeNM+je0BesQdHBmfyGBHmcVdiX1UC6cbiNG4c429MLhXaMvkUyM9eTW+4KUfK
G5SWKJzC4PgJ5dnW0UK40wcyrP4OozkCnasbtl2KFQP/ZKjEbVujoe6n4RapPFWp
b0qGPBdsKcjNMJ17XwpBZ6ubj3KedizeNRFlwYp1rgH4SEga08jjjrC49th5Orkc
DFTMel0Pem6e1Gk9DsWZ4MB4iu5kg6EMQU/3iVufbdaqPUHgl/S/2/XlnISW6/Jl
VqEwcfl+y8I8Mq0mz5iJ/QXtgeDJvNtsajaEI+FXEB/P3cVvnzusj0MHVUtImEZJ
C/z8eGQLGh5kxX8Z5JLw3ci+T+AYOuklSjSMkGKTMk3QskrDXX/ZEwHUzcGNqdL5
oriShvdF/pzBg+64oF2V6nwbp/1gvR/zPuhjIz2RkfqIpS28UlC2Y327UcUCDL4+
0kJ+MbQR1motxze/DYHKcWextES1WZv6d1+8ONa01+dZ1yBzSDteYO4DYtdCQJGW
92nGkUOWd+IdV2GMCf5wkXtCU2tK3VFySTH+4p9pid19tuXO26TxuN0ji1mroFjy
D2GOh7RKmu0yXJRjUKXxIWse5/TbZjnFdPeZwKCRtKNjwiNXFjOuCNvrqCsPKbDU
cGLFV/V19VDG7BJ5Jv0L4aSK4G4kvoh5OM39m9JXpQcp4y5zcl3964Cmj1rFKvTL
S46PArGdyluoH+KjfvWZgQo+bs1JQnUnEA44OsMyyDTpJGWd2qSlTbo/6TaCzSGi
JBAbj+iFIbkrlo5u9EgyUQ7N4vmrsUz1GlROJVKk9TQkm/mdyGvGhxv4aCVKKOvs
VF00kVyEbHjeihreEBgy/Mf8uhwDCX2yPGlBnXaoJdhX+ESrHQUszvbzpo5aniPF
G2ABwzf23fa+wBtelufhHKi9IZGwHCpw3L9VfUJvXr4qWb/rNaRykzCLCJqwnY3C
o9clWcHuovv2s4szOcV2CHQueYl10T6HRJKy44T8znR6K3tG5a8tfT4Rw1gQ28dd
oshTbmbMo5G7phzgamrOJ+DQX5ix+qTBoVMIxsaEQ6p4hf09f5/JBQmXQY1Qcd1E
pCl2ooQQqvOCoh8eje+93IG1Iug1EUBH/fT703QtVDF7MJKVyxdCUSXmwyjMmJoW
FNYxWBsEhw6/a7d2u7hCKkWRcUbJrWmASOAO2LYSxORxEoXqykJIx1cE5aVWoVIF
Jip23vCQxvfOHXM3hpt/q6HlKYsb4oM29yjC4hjTLfyRc3DbTDYXSTEj66zhYk77
XxSc+k2lB2T3fvt+yKUPfeZZxgL7uZeQQSFdP9EnaEMQu2d1+JLvM1Q4IsoNXR7S
I2f3P/M02B/c1ibopGwIlvi1hPm399MSvXD3WoCTfWiyNGqQ9Z3OOa3tFBpkm6BD
pVafgvCdlDLi8w8riF+5MymAWju/tzEGCf+MJuF/nxw7QyPYyQgj3xz0jrbNQ4Z2
XJoQiM0KZEBoJBOdAsnizdsDjwhVfp9L8+EerlQWvXI//xNOkpabu4xLr8yCxVid
1WXWUAbFosrcgWrMVynnLB5tWH8EL2Wq4XeuPMdJ32UTFrjrwe+uSBG9l8Wj2f1G
YF1/ZE45VpqPoYOrm4skSQkO6UJ7mwgEAwb3J4WUEiMXn+l/JB3VUMBNUPwqEPIo
cyrVjU0tGWE8G7Cji7rXNDWqDbF12OLomO7rXUFA3DuGCnkL9fYa8aUtQsxbdeX9
tJMKNl0TUsSiwdgtoGASZdjP3gjUkyfqcrSB9DBGLJVSmdpvhfnJiyTjp12/dNUO
12EvO1va7RCDk+0CVi3Ui71FmUwcigB03uFaDEZAyoaOqubfULs+dqwg6pzXDRDq
dbavigLwKfIW0eQzggbAeQU478bFn9VXOQWv4bfthQg69BUL1+IbbuW/MQvm+FKq
evnJ9+pqnu/H86YdNtOLnkqypgDqoeb9NjGJCvSo9r6gIS6EhZK3RLsEcy/4esz2
Qk1vA/0W/VR58OqMOeDSlc4sZJCQyXvR9d+avtGt86yTGGvoDBRuPMejSO+pOJF4
Mfs3KM5nnupC3W1Qa0E2PgySKGQRN2yLGhuIAKXMhoPsOsn+OMWC2p5gIt9dlOSH
z7p+mnp172Mn5Te7mEq4mPAaENsAwX8B/mK6nrHwCA4mAp4zb12T1BCV4NFLHK1A
AoSePOEp0Hgf1qNbVMbLMzbvtC6Dw6hsjmcY///9Lqz34ulLgLAgFCMZnBnCpA18
0R4eLXQ4gGYbyyH9BTSBqGJw7ZLXmATKelbmiGArQ7xN562tKkpyIAAyJ6ztbSwY
HkwkcPIfNjJjLG72N4FR10wGIbDRmSc82aer40PLtoaTFJ6l3YJA7wpLHOTW8BUG
nzSf3XqHXuR5gKUmXofm8xHR8SaLEmqwUszSsm15ulcV/m5hOq3igZ+5y6R+eDlX
6SB75pDeOtFWKJtqfhgey4ZzJP/FV8dEA6qPe4wBTTDFwRs76g6A8r0F9/I6QQkE
EGU+uMjyRwhP1cjeo6uFboIML3P3YG0S8VMENMNVZlS4hOho6ggcYM39Cma+M/aA
19S3frf0v6ZWz8O24xR1KsTw4WzpJru+DuM4lvH2gSrxpevp8SmW1JF1sDYH7ze+
LR1zUjhega5ifwebXpfrxd+4DRQbLfer6ZbRHOw2A7T8WwegxVGfy+ngXk8ouQG2
PR5R/AvJZQo+XN2QWhF4EJ/IF/PboIOhLdveEZ9a/9AiI2mdVyYNi0rQVXSoyx5y
evTNY11tUDG7x6n1ONdlCcZ+P4dhv6mGgAI1oAiwvv/ux2qwKi/8qtBbwrVcIQ9f
95aZ16ebcy4UFq5Ti3olbS2FyJYRQOZK/7mfWea1OxSIJfgPIefxnTVTzh9BAqrD
OwfH12Ha+SQyaPEVIE/X1jdLz5f3GdpYFLMiMYzaYkZjRiaI2BMgle1WrQlDLIKs
P+rjDXaxL+orEFmel9RwPGYOATytcWu/iuZ2pgdVBhWPjw1jWk2hOL+TmpLPSWPv
+FbRsRzrrBs3sm5gxRdp965Yzf2p2rd6oWcYFTjRY37NXEkVUvubp1i8WVGqDvQR
/bPkdsiT2lH9L4FGb2xpr99vf5nZsqsna9OSr075teHX9HEb/+ZZWy1qB5f9pDqB
e6qjgng0oyjkLMh3jPUjRkMF9cDHXvLVK1uPcmLiR7oyAWd8xEVZH/weq3N9TNxE
7Dbt8Fyfd3p8EQh1MmC0DCXAo9fF5D8zh7sZk4nowHiog/r0IdnvWf67sRNcE5Jk
Ueqd/ibgl5+TwiIgrAG5qjpi7mni1jnN+Cp4b03riLpqySm3do7sCvTBMutUvhP0
JK3suJfkOUWs1cns8lB4F3khgbUYx/JfAF/GDQHU1Z6n9PVw8X/h/aKG+5GRtiz/
B2sMc4OTxKoS8tpkLIcUwpkhvRsn4DodGMlMMZhz142UBcVvCTE3JP7oYKYVUNKw
CesoRUiwo2V/y2bOpiT7bJE76pVqmTQqrw4cKoVnui4AvdPuCg2/u/PLbpYmWlRt
ysl24xJjin86P6oPYan2zBSS+o3sJ5ptpkre58FB2XNoMlks0FqVER0ospkjjyQx
XT+S17LVf/rM/ceH7qwmlLdWvhigks5Xpl4XNbD83cHCktOPqRXxIJHAPlrMepVD
mzZg/zbK1S5n13iLaAOBnvYvfhjOw3n03TDYioRP1MjWAGeaT6k2jEWFPzP6Ede9
6jQzfi6HuujBJFvwQtKwIVvcHN7yHRGGsKR4uSjk5LGMFbCXow0rCLW1SCE/Nanx
PQnCdmQIyGPJq+Y2VoM/e74mL43qEAz0APj43vjky6bNLnXMat+yvyixiXxAeEYO
2BC8z9Hzdnxhi+9J6OmVvtbJqr0vdXIUaIfAOlVZLiagzqXGXlJrnDmF+4b11wu4
HwmldfBEmqsq2L2k6dqFWFhMbbwtwEuTSnyXKZ6WQEapcIkxPnZFeELDYAguPg6a
7ZZ4EUJ7IzbeM7vtdPwxHQi0GgP6+yaVvtqbNl2eHGnf4yi9+st2j1rfW6n8zWA+
xbE5KRu1kMEe4LtHW0AjLWc+/8mEJ2NkzCGWe+NphknxEaeo+ZMi/55dJJPDwX1D
K8fSqmV4NxC/xyBRwPFBw/UdorDC8l4bZgZv0tBAzTnK09QsmIBb0abuS5LBOHYm
BKi9xonflgrFpqm1gOmu5ScZiibI6F4nsSjGntx47+x0nGPvRjeuUQ84brwbH/T2
F9Ly32Lwe/KAaBzISQ0zyTBU05z27bTAZYJEZkt7MayQ97kUi/H+vm9RUR012wrZ
FgF9cGHezFmSRjowOh9rcxODU6UxPDyKAsesV3l8pB6n7i8FkbgVeYnIDAaa8Evm
NESklxPjYnwqe97bKMQdZ1xrfGBUaRg0RKrciu/RwQ5eCqUE3JJWHRqs4fHwvTaE
obzxBPAFQyXluUaI4b2vkyjL7wAO89VS4ZOIrnaioTlTg3amIT2nrUANXB9fBUyC
3ql0vinMOpguybsb0WUH1nrP5u6as/bh6D7Jx6dcQb/0MreW1KHmNbccGYjx1bX0
QTEvhVc3FUi9LacN/pVGw7JZnnb7eOEiF4b6Veei4Ju632uC4SKFcYmHcKyzkcc9
hdjOsAAiyI1g7B+EuT2I+ZNLFxLB50ezeE150eJSOfHfUMU34NvdyBYpr8sE90T9
vxrfil89jB+OnDQYT3Iri2Gzzk/CFfeQPMQjLaF2h+8nvwI8GaJ5SwoKL4cpeTnX
QKZyGtgXPPBh6hAsRtZceSoOJfFvySSn2AnFzsnijwf91DMb7i954QgeSet46qoX
ziSz95BLlXesoGlmM2C5qeZ5h+OiQ0QJLN1L4YWCVceiZpbERQPoa0xrsQU+yTFs
Nc2Su/6hz9jiWU0MTtnDDCsFTs78X0H98wjG7AlGMFyKgraw09RGsAiXfYFbd4ou
bl7C+s1aaGWUDSy6VEwa52q5AJ0zZuBULXdn4O//LgeAP3UNYCz47tqzqWBp6QaX
Y+elXkyUlnTiU8dxqzBYZM1WkBsl5TYW+XIQpeY3NA5VFxz4e/39T0wbmXH1yFnx
ydaIbn3WFtllue+jwHgeQOX1l6bYcOovOJxyBPzUhE4sGiugRtI7HNWzjAnc3L/G
//4apQaFBEok+Lc/gZnodA88ud37Y8aQnzYnUE3TnBj7y+Nk7swn6dez3Ibmf6Xx
bj3OtkVZe3ACOcVn3KvLn4SmZ/WkFDNooBuF4XnPj7mZuDxljWY/hdikQpbGSiFa
NlVOEY3Od0fp+gk3neo4leJ3I+H9OSmsQmvu51LaTq7CPLXn+Kc8/pIx5qZ9gUga
BxT/+tkMCRN47vIMcdalau/i5JovMoG64ztdgG5CaedDnztX9knvYW+WNR3MIFs/
Sk/6GyC6ZqCbffhd9wW2xsPscmqsFWmURRQvLxan1W8tHsqsJ4vvV76RR0sjp8CK
qL2aVrc/wEEAdHWORtmN/cqmk/jbCjelH2QzAZdLPRyOlad3OS3KEtFiXIlryx1Z
Bx/d7GjQ9/WA/qkPxRJaowaqqRwEoN8UA1rPrizwsBh6wnFjkdeAdb8Q+7UF8We4
bm8CMZ7i6dimMaiTY/y5ro3jvV+ZFk72rP0Ae7s2yMwXcu7dObbo+DZDiRY14lsL
dBr+WWDlMqSrLMqMIAr3jKKOZQQL4y8kF21YG41KJnN5ndnX5x1XwEdxuCj+YVW4
UZu7mu9FBhSIM20Ytv5dRFeSyQwwASlC3giX/IN+9YOo3QiM3ENvp2kOUJBvp/zx
58b7UkueLso02rinLyCEX1qQdPgp8tsDdw/lQc+AtdXy37hC9CIZP2EgZ8JeVHif
wtpltJptPlnLFMzXtYwLzDhjH0ZoovW6pN/3K2uW9K40/QlLetolbwIZnSNyrp1b
XWBUOeshHbSY85O5KWJj8A+bjApNTx7h2uuikYWU5tZQhpGCP/VuCLaj4yzypreX
yCVAmJxQLwi86XBmPpR2AXTBmSPQW6o1LakuZd9x8F+WrNSKqZemy56oSYiXa4m9
NGW7IaoO14XKkeAKlJQPUrKMxrzDbq0m24lsSOmnKnHbw9XeFNPCyR3+YDuV59hj
1Lw2RsNEBuP2VLGFtrO8IO/GfJcM/B1PMMdfhbOHkAbMqsIg95R0KPbMS0j6de3b
RW3iXykXYhaqh7S86aR/6gBodxlaepkwaSrXzlFQK6UV8rT2BndTJDS/iPJBFD2M
hXzh9cN7CkQXiGGCzYxsJIfTigxceCOMaMaEzuzY2bN3StkrEGZhetGFACwvoZOr
Nj22Hl5/N0a/j0u9KceeqAw5fJu8ukPharu6XFjUFABLw6nW0J/DsbmbVp5z865f
agYDMgWuYslDo6WIj9OcYTTdCmNLfeH8Zpmv5gesgxrPJZMPz+fui9HuVJSl6HE3
4/ooIYp6YMla7o6OeeBuxRxo+mDzO/pvSvzerf31gIEu+h+a5mIuRBi+zfI10gwF
FTIJd4S0dS1aT2DEuY7jqe/rZRW0TyZ3qqh5Juo8W8YS3GyIFuZKWBIKDA2REA/k
dm/GXd3UHN8nTMnB8uQhrdEo0xqqR0EIJLrUN/Cn8hjztUJYuncN88cERSxahXe9
dI3JiJJ5sVqph17K0EnZVDntQMNYvRtG8/ERPSkUV5XE0S+p7oenla4n3AZq4FFB
Y3GGmT7d4w3PlGJdYTe0NqxNq0KT5jMueLAkrTJbbAUVSrWC82ozLdF3DT0zH29c
E/xXqpPXIdQ8C3LnE4EyN1NbTnp1FlNdhFrWQpE/oHku5kZqYQmplD2W8qGLkIkm
2iFT1strOr7s4NwRKRWJ9juuOEtsZ6i2GGq4zGl1fFnfxgVLlaoTlHClJiki4V0P
4I3vLccxbUmZCkfGdnibBUVS6CP9orhj8GibeMIjR+/IiV1Ugbu8Glv9m+iiPyUO
WdJErdeIHmah2b4Xc2VdvorX6cAHIsLsfxBHgV1A6H5oyfSo002XwvFp01gIT6rr
FoVV6ks0PdHO5h4/dnNZ1ZBVln/J8rtKmCrXN4aIRNI8thgX4PXizH3Ajg72tBTg
lo4hfKGB95dfWofENMuLYhUmDaMM8oqEPuJFtOF/l6QPBrVjypwralkQc9xHu9Ls
RyVuMgjFUJBh4YtxkoN/ASrv6/xsmHhj6a2nNZIbfyAdUDr0YEpZ8Ea+0hPh5jDZ
++cNvxnGLSY7Ek0hJFUb9APZsxrbrMnJZ6GwxyjLBf9BSteLn21fZ68RbPtZP3LJ
YJcs9Za9trLKxbD0ml91dZNXbqhxtbhCemvqB1CaByL/+VycEZ6hK0QhAcGC+8aE
VNaA2zEgzUY3ZpnP314KrdtjUpisfHz+Xw4WtAjCAH9GZ4FlzqCZlKp5y+IfJ4lC
ikYZPHaqoUyZ/Gs9s6SVdod5Vk5iPLR4aO1itCd9NEfXx3ha/qJPWVJcfYzBFRtj
IoFRUmL32OY2J7K0Yd96UMxcVNF/qkFnY4TzunDCUW4Ug8QU5eoxAwOaq1MyjoWt
KCZtgM1VzRwAsqx7VGjzZFKrHPfNk/R5QZrTB3Jo/H+B8Pe4QigEHDkWktEEK9mZ
EsU9BrQkrFZpocP4OAEM6ch+BKOx1L4M4ZQ77xXZb80uhaOll/Pye4Hfqtr2LuH4
QC1OHgb//VjHYJtZC3MDWbtN6ZGcfGpougs+KIsWgFFmbfOCsdj/WILYVWYenaQ9
/rhzu7xWZIdANQeH7kLCyj+fmZfAljgt4UuV3L3ih8krOyPt5MjIwhKMdxfhho9u
jrEIPcU3pmrj3Jr4ta+zjJ96PRCxQgz+s5THoOF1Y8vDA8fkc3Tc2OLgYcFssZFD
dHqwCGSpXGiyZ+UpRdSe279uElJ8RoBJOCvQbK4sG4l+Fr08DFPuPnMGEiYOnO9D
6raj9FW7y2+VE6+fAPFRAiTUAQMT0EEnJWCXo4H7DpkgzE6kUHo9DJB8WQvLIkU4
PBPyNjRoHaX7tWz8SmZchi95oayunoF3thT4QCIYKNtkAbSdt8ioph5/9ZdVFCVl
bDr/RK2zefmUU0jqeD0uOhUSlu18/qpdprIzymS6bWWBV3qIJgeoLVFNhVqAgrMK
he7gjRMAZ0RHr4XDU2M3h4xJCiFg4ELuHlwGsGEU+pmjLn+8StATwA1isAjeN/Wd
rhCSQyqDMeoRI5twZXhxFWUoQxk1LUPn02VZxOJsQb9tlXkomvwtuDP2cVXmFJ/R
SGLbF5BnAw26mMHNDGx/sxMULbX/MxFC0dC/HYibbOvtAPxquoK9DM5Y4+RWc9Xf
eszvN5hjT4imY6slbFKsoH9/UF1Cs6KHUOJnMzMZPB55cA+LS6NfS1xR/SjV9hQV
jdHan9b7ha6pqeNhv7Ffi9xmqrFPobKeLUouf7qUxrxmteiDhILA8SpL28m/4drj
9yV9x9JVFwZWEGRjxJHAw5bG4bMHgcVtoH5o4be1b1NYg6zOAAidllH/1RnDCx9g
ph2mNmfiC4poQJNCWqXCYnzeHHgUYvjh60pXGHmOXZTFeoFHetH+28tQBYtfgb/s
y0iFIVp43RivB70bYj/A94Af5yx4MR+kpU/G2GbIHCbuRPQ6q/hSB7iYbxlKfTuw
24UOX/sfCVrw1yvtsoG8mA2CRGI1E76NXKe9nfUPAHn+3cFIOZsT41p7yLJJ/J2k
6+Mpvq4sjRjvmTmfG+YvEAn7sE+fKxOVPY7AoTnL/CcnEA1a8Jwiuw84To6Bgw86
uz1Ncaag7bxaBltTy297wJ+ZZK2OunqRRJXmQd7i91YB8z77mSShH7y9zM00JgWi
QT95UFh4isKLYrPVPADbg5hRxKWJOKLK15DwPQJHw8yjhhkKXPbdLFS3KBS7IEWx
CMsUYDihMxjWWdfPd9jkzDzFqrquLwWYjZEV+k+nU5uHZMQkMLbgeogllIo2EuB9
ZXKQf93Hb/675SCwF9CYayIuNIlIWfD7makytoRIRNyELPVfwvgDKjhoEmhUTEF8
TED8wqPQHr1ktUbjTxYxqBsyKjAtH9T6lC5bYMmOAO0WoCmLlfbSkoV8pdAEz+N1
IL/jeBBYLVWBoSumHUqbOkqthN6MZHPnQVWPSnJaVVA8v66Enim8m338DgN/+9WS
MiEfBbOA/YfvokONNHEqAbqc8alqm9POcGNzFtXv7mFZmvP/ShY2cKmHi4OOsd85
NdkCLcFqCh1gzR8p4cJlRj7h9iCTVfTJdDAmgZNGf5d3ghYlYi0/8GtfesbaZgn/
iwSXUaYkt5sIvySbr+SzYT1ZHHnbGn3ZTUyGTovyL5RLeQY46JmXL+dah1Ig3D4f
whuNZYsyDVm4uWJdVwR8l2dkSbL/xviGg/fBmxkDlE2UaXx/W0OyApjI4dglWAcG
DcjDfHDdyko8rqohz5+hnrzKEoSLQHJbfBacMIkQY0S0nj9vZWgDuMhRL/C6uNd1
8zXhEd3CeDjqJ/R62o//p9dnsnjXZgtkyvTKq6zunLIiuyL0wcnDSpBVI0wmLauM
g5nVvf0n8YJNZ9eWJAmFendPxUoON2Zgf7tVmAjV8fUltnBDQHzuf4G6omgb8blM
cGL/EG56jn7jgefksMwCgcG52Stx6SJPbLLXaNtfCni4KVyMtoP2tB70Ep7eRBNO
tbS+Qau0vK6Zv9+RJRbRJjqdH/MdqM7AlUc4oN1QqZotdRcs+xhjHNoF2JZnFmP7
K371qxpoiC9f3BcZnfKkyo31a7uWt1tmR+XcF/+jNysbpeh6Ci2cM6lcaSFwFJ2a
sqyKlP1NLV32a8BiD8fnlHTgjPe8eR7wzQEYeLBLYmMMqBvRmf0Ffwoaww9n6o1G
5wuPZYqwPD6JdCKdT/hVDWr9Vnw1RpsIWii7pXC/BroR2m/tqNzIfjJhDW6J6ME9
6AsgtS8TX87vgff3DHVxpOFleuf4WLMoRPkNzq7U+G2wAyWdghFn75Bl20A9xk+q
I2nA7UcqWNPfqSJmmgEZVH+IZI7/ysLm2/bPKXVwWV081udfG6mmircErAf2K01U
vivD4D6CpKdQIFq9NC7Z/epEcMj/jq21gfi3TQOdYC3/Dbo9LGA91UFzSV9HQP3Q
ei+zRyOU3qwOKM0huP4I52nmgTooeD95HN7/+7cBXv2ZBnycP/RvKuLsZNJb9xFy
PGoVc3DaEKvsib+Xh2TTxG/OZbkC80+s9Y4hs+tHEZ6Mn+joSEkmLbS0T8MO/Bvs
NCB+dfFF0qbVBvq8DYHQdUFaOSoVgzpdinkPHZ3ISRFyHZtLou5fGtVRfYdNfvFL
5va1AY5z10P1E8GOguFkqeDzYrq0vp8VQ+OFfuonatTrgeMjcbM6D/4fz9dFdwgF
lOgQlIAPr/2nizWBKyG7SwuX3gYZY/7oGZQ/Ck+8R5k5qTcb5wSM733WCs16W1Zl
UHrTXXn++/73KkNDYJK8yhjYCQm9nskl896e0q6A8KIKyaulgJX1vKYcYbEn55fs
kiCn2sDfJ2Z255ln21fYnIM6zaCFGIt2SWIkMWX9MjFqkd20Eu5bApcRR9OssC1H
oL09/FT3NfxFmaUJXzPFrD5pbvqbSZ/+UM1GPXp6Z4QcCeZURU62beoWNt4h5LGn
+iZ0D9eJkTbzjbVLaeIn/0EjamX0AL3dFqgVOF2D2xGPgLy+oMiVjS3arxYS7ML+
i1TWXfx5GYx6wpIGw3PiuwYzkqCNZx6de+3PJf0uXOxOqaHp1tJlbfCXSirWyt4t
t3v//dSxr2rOsh0PEJYgz6eAg/4BRbekMhNg00yT+GBHyFVEp5Sx0hLPtyNTgnTw
olePkYNKcqS12b3Sovisbv31ioh/QyCksMwzg9yE7XfuFkFif1Plrx6JB65hZm5M
sInPHXOty6q9bRG2mC1/+4PysjVSTMsS7s3IjXXjMOesv3zA2PrOwgreZBn7P0CS
4/V/PXRSsGzSOYZ+LmzSEDaHdZyILhIUCKf7Ple/F+73vycCZkHDvY16Pte06bL5
dW58dQKvL6c/2czUlkh7Ajv5TkKAzrXeYSqJ2hmlosabMEfFn4lVcBclDnc7dfc1
I8wiClfiB6yUTPZSSs4MLGnoRLNVI3T5nXTVOJ63CwAW3SgkF5UVHMsSm/SEziGM
mrIV9F8PwW5qFBQBsJ92NZHYJQ3QKOhuJZcKQEuvem43xKa/cC9IJLEcBGPfUks4
55eQyewgbt0Ufi8gv4iDf6SO/aqSvXx2pMZVfQyIyoOwNriaRosY6zttUyeMxtAH
d3Zy9H9CId9zTRdNHV85ztweuYz26BuAKNvqqBwguKpGXbLzKXS0imKT05cgO45G
p+KEdFjO2Coe7ijel00q0sFd8hJf0xFmdieJW4U2ZVVC0RNlC2aTafD21V+Wrd+7
eDjSry0eOdsrs+0TfY9Vr3sdlj/q3mEvay0598FETFwdSElXEYkkTyeM9K7aMvRC
MN4dwIK42w432jNRcaytYnPN8mTJ0XYqy4pLfCT3n4D8AfQ+VWoYOwPWxJ+eiLJF
MZkcqFlkM/zbddWYAugrwcq2fRCJzKfGtPKkoZRXOgp2wFyHFwUGnGe9uKUy6bx2
853sE89Ao9Xo2nDaU64LzBaDs0yuAqXp/7QhqK9yF+zwaPxAr6mFH5AVug6EAsX2
o14dJebee5n+Yuld6BVHcro9uGmU5ToDRgo3SNLGSlopDiSWP9wULPH2jHIPpyf3
T0yPItBfDIvV984GW0TzbWOhKkCO0AO0AtaQ+N+Uwhf8Yu6oFyWc8QcIbycusOaJ
HUxzwmAYh02N3Rb1nkH9iHG6Q+fY0H0aQdYGwBtP0sDz9vwKTW/A4gccjG8MAy3V
KfR2gObC2dKPn+1226EmmpdmqjCLfQru/XnkZr6s92CAAP3PwDOdUTrmFrDd2P7t
`pragma protect end_protected
