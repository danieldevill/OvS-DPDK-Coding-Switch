// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:34:48 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Mskuwkyec9LcvU9svyghOw1NW352t7SaRlp8lFZA7gX8Bp2BFZ9ir0EHwNvJhXHL
SSrge0EYc4+an5HZV9EuS8FjQLqjN9Zr0nol+rFhIgYtnW30ikLqJj3lHNlQBogM
ZRQFTnnhj9CypTtsz7Tp68U5P6mVfneBiUZitObnM7o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5456)
2RqcuvXy1+1YnLESCeUAx2KZhwQUZRUt6T4QmR5MJAO1PlMFOFO+QpY3xHKtFF7m
CDWMYmTOyhZGj6hY+v0G1KQZeiRzIJVhtIiHct54v45za6LLzMmhqqKh6NK8Vw8L
HQ4cZnYwqn+gvRtTrZkdD0bTk9XZUte6+Um4CCtd3Hv376G/jt8wGQaCMpAARBtv
+2j3qqaKgZ8BJDCLCJNBUZ6qAh2xioy8tGx0Uf+RESQPqq/0/DgpIzBzcEJlONFi
HBv+dkV78MDbBg3eZOxE0vFg/fyB24z4HWksq3874skY2eIo7aTiQ64W1qxkFt8Y
zUxN2mZxIK0pn9H1jbt2PVOcA6ItJVpG+YtkXa/WXSeQ7JPOs/ElRHnEt6qgicIi
WjF2uwjAjx3fdvd2ZtYBSMpw9YaJHV6Dxc3X75JhxG1AZ0JPsvRL+HVbdt+t722B
HRjFC4CF6hPg8kXSPiBSs4QlGANU/5aGLxuU8wTJ4S6GKWLe48BODgmWKKZ0JEQY
TG0EEXu3idyipkHNMXtpbH3SAqhLxqLr9qNYXVGWiG3W6rupKY68UJv9nbQC0+41
AaRNX7bfKnknETdeSV0mUpaEUJZtPgFdRdoQrcJVk3Hdu0r6CJwOdRTAC8dEn+wQ
yHFw8WBfN1G8I9CoEOPQhMFgnlX7yDJdNCTk4/TOCrEe/4ljuMm5ggP7XHj8EC1E
jQmmRJj3nnKD0z9rwX2YY4zKNfw/jWg9Ej9Au6sgAwW+t9o0sAg72FuABoYKsxBf
qY4sZOVHULqGMJvNlyJpoSGyslhZYTovzWWxTNo9OIerZI6cUNl8LlUfqFtNlzE1
wqcOp/YGgymkkeW9K57n83TDKLMF9hHFM+dhRes26lBxdOo1ur3rfcXUFnBjG5WZ
3/+z3TQoHFDyUufpI2bsDdxPSZly9hnpuKd54V+FpezdRwRqmOxBoErAiXaUlCSV
wWld/9DHjaljBxSWq01EPStTeb8X+jAHRyxO36M6MshipPH/38JsJdv0LOK1CeFB
Ncj89MtYzBTFwAwl79hcV+BfipWQxqkirliGev9m4Hls8UAghMUVH++Ml8JnSXZ0
3ZY8PMt4hEhR6KJqwzIsm5P+CHMuVthaQ0YH50/wq7jpMj3FbUOjT/o2ZwWlzh1E
s0fKNoHRZMHBnJF1ST26r8Lf5HmYGn2mDMDilb2m4D6leLK8YjFPzTgVT8GR95ov
G0RonvogJa29FSPKfnM2cx0gZzmixKHEKaXnjWcW2KEf71U3ECc0LFu2cYSAmGQi
JeA4jY+eznb98OpaHvLEGPOKzldz/FEZekipjSdGLUm+MufGp414coGSITpEYLdc
kIVcAdYDJxx1Q2lu/g2ppaVpL9nytM7x0UHPjXc/hzR3e2LKLllrOT2ueFyCM2Ya
qvjkccbPhyGQALB+yBmLMlLsi52QzNG1gVS7xNMGk3OH6UaVGblWXTAZgBZydqdK
r/ehw9bsrfEhumDPbtvokuPQxV/LMfYpbniG57TS51UwQYkYSyXXk+UHQR8C/MQA
jETKGpe7Po1dwnhTp79bJSyO6ib4RZaWh4g9RA501NJCuHAQ2ALLzbpqq/sJobJK
QJHRySG2afhHi3HH1sVJO8iXyW0M7jWNjPBfzkRKDiMB9H+R3bm9hUteDdVKME2B
FAM4WiGHIwwvEKu0Kg8RlchAMs7+KyaxC6ImKAmMgH1F4xvm0S7Q5u6+x0kLfFwK
1NYVxCPN4gRIFbpV0Y9wxX9AHWl0jA31JZ6d0xonk4Jvi1FeLUpLC4YSV/bndaY7
9WldlxHReeYxjHeVTI3arsPTRBPupE7R0KBmEepoQU8Vi6yuhzpTGUK0XTKGpkl6
gbyZ1lcLHWXT838KrhyIT6pEjupEfF5iSRgnbwvFxFxvknOfQMRvfQqiFSvb+5pw
MLJFJMSBES+8I/Fe4FouVPsAjmMYWq/UipFhQcQ4290eBOROZrM9nmIYsscoOMdF
O1JC8+muP0v4JM8dKSRCPM4Jg/osBaDiBvs5LMCV8GhDVdGgmQcO8NWlIcXiwZFO
jdP+lF/Vgi1JAo5/L7D67j+VDqy3wS6n7aqvkELHondFaESGFxvy4nzpB3ReSPLx
RBpZD5EjcemOn2Sj21NIq8MeHQFDVj7mHHqeJ3uMSZjqcAy8L0XCHjAuK5knjCvE
I5bmYSj+MkrwZWw8W+hQbRco5EYn+3Cqf0JoQxEciywX5tDru+DOUHqzsN/6lQPc
vqycbxlW/o53DcwXSc2R+9AMS69QmPYlMrVRxdKTcmZeiLDfo7FFNCfg6wR7JWJ3
Fo34oYK/J5eUDWa8lTer2S+b4ytzyErnN0ygUw7DGHsR2hfT4huAZ1m8unT5jmV6
prWuaWj5nJRj2zYZTtTDpjJRGhmOgtT9LjDrlclp4ImhTGM2MskcK8pvBwu6TpIS
9Ca2qSF+7DSvfJnjE4y7QW6aTs/Xv0gE/Wwpl2kBljwFRCVafpPPPZ3iNe6nj4+B
Zkn9lQlh01gXsnHRLaH7XlYzcWO3K2SMEzGc4J5Z7TeV0DpRRlB+8XDOFjqXKccj
6+fbyw113XnaVQpPQNkv89dm8jkY7TWlzkXpsKm6v0rBuPVM/gUefY1gfwlb1Z7H
Rt3SXdg7ADvYT+X7dWF9+nGCTyNAwN4sdxrdyNeCspBUeM7jkCUisa/dHfXV/Opb
FB0mga2GAwU5ASB/BE0qt4pS0X2AaYYyrK29mdZa7xci+S6Sh0PphN4yEkvsM1xp
jCNZoj5ingcjt8AT/UiwDiIHbGxFZMg+tja7rkPfOyM/o++biXlyb5AjPQzBaOvD
ROxFRjFhGVZGkV4V5EdKAe/bAi9f/Po5Bmm29PuClsrJGVNVa+x9+zVsgiBIEYAs
vNxv8hernM5tU4c9sQ2J1I13w2Mm/XMGh96G8aHstCQmzmax0FLFDCwJIqA+dUXN
GswcG9h/vUHKA2oINWddv3oac9qn9uTFSTi1sxwLZhgQzmc0MATpKQ3x6hJPOBDc
i+xFZ8qLZ4c5YxNEA9NVsjo1ifrLW6EwDsl4xinpvDKG5sShgKonekFvBV/n+F2q
s0tUwJaM9CeckxjnhTB5GMN+t+AKor81HfWWOEDkPcxbpzS2/CccNXF2jt+X5bAd
pcKCVDYY+i6gBXhC0SDwGMTvyayUqi/Y1wl+M2JigkmH315Ndv7kU+cyhknOAumG
suzY5h8Mf8YLYiz5EpztII2wlklAPO2AwOOQHknMZqXjvXFf0/9v3h6kxMgjHPj4
/RyJlYZqVEpJCYgGoE5bCMGJxfOOXz7UcYjz2fr47sO/lp9lvzzW/Dq0Xdd4eyQO
3rsg9ZIz5KejZ8+HeMDhFAVyM/Iqf5iY5E1VU077bmvcQDF5GSZm++d3U/+kNZsv
w+eeEa4H/jow5iPnhWRAHMuBbGsFfo2xp/ODpw66OBHniWLixFiGDII8blAVYdaS
SeHOm6bLGEYFyQZhaIPKzsMDdL2zRTJk7XNhodhynHnP50xOkWzCxq26Flp+KS4l
9lmFtevxpya2tX5I6jfxkOZpZfVWzqjGGM7l/xRVWATbnEvUn8ZXq7MOjNdbhEi2
ARXq/B+BehLV2PLGXTn/rfvzuWvaniMMR1r43CIPBSIGUgNfphe/DqA5/U5k65Zi
Ki+P33bDi+NCy8qlosGW+U3D6YMxvsPjBhWugHpDcTRWQ4cfOLgTrOwQmf1kbaJH
Ui1kcQEFPCYYvzPD1ELg8rHPbwjCjt3RouvskxoFuqj2Q6c8ovUP+50dF76CFDuO
rWxVJEjIQVerDiJsR140A5cCgxSsZLCwY8ifnLtsk3/Ndj3BFgSIs3pJrXGghcgp
eSzXCHAPKPK9TAdA/sgGyWsBmqTDIlcQCU4S5WYt4jKPojlM34NNrGATF2wzVl6q
LFwXdtnR6vQbaghxwjLD0OHmamLBHLC/CGAFiqzXnViE5SqDGOMjKEkWfvJ8b0hK
Ch6R0dMfc+zpPKF9zAwkXEjbYRFDx2LSn8aif07QhJh1o35JIRp2ixlsOQHGIzW3
24PkwtvX9GXq/KCqcUuumvIfWiNpEz6O74w1ZGy0br0IYigNalIDJwnUl1HfOR2s
+RkzvPNMyCP7+BglPk77UQE/m6MKjSlmMjoATY8peEZNmsBCddkq5zMzh/n4cnlt
r48oafNEuVRds0Lq7ioK0PcDg51l0iIClXoUaMiQSZiWpRu136EjgLbF88ALozGU
dNDr3TIci93NinSV0m+sMKvGnxdcXJaRPPgnfTrTubfhItMOfFk1G+VSb99bYvgX
F7ORLuOohKEZbZemWLOdTcl7rWnbKPPOSjsBXrc5tBfeNzNzcMrtJlNzJyHfQ7fu
tDMgXw1rHICt/nDLQhy1gl4vKZR7fStu6fQefTTMielwn3VaHKdwAm4lU6KUB7gG
waF/UlRv8JIfqvNMokgjqCJz+LoTfT7yklr9/y7u6D375PRVm3u7gwVOffe4PJSM
1QNpSLje+tgonJPZLhnwIfFMfGbXVFEb90LKnE4FeT4YTTdHaY6uaSkfA76icI9J
eoxoJWkWsEEVq+WZ8sNbmNze1NsNojq8tEFWgxc3JUmhv9hIZyTN+KYzW8EvADnj
FyukpeuvXPvnjXFWgRVUNi5RW0F5QPPTWZ/loneEEKBPOV6BKkMfL94ARMhZJnMG
GwXpT8KDWJXyko2p22UMiulbOGme1mK4o7tyjfCgoOSNfv6A4VqQ8wXt8qu0SLeL
IAXnNuUcmkkpZxRAtoK+buVJnfa9uRu0LCTeIwrSBC3cyMrEwq7+4IRQwIn8DN0z
UyVDMviEpwZXg6Q+v/f+TzaE7HB+hwCVhmp/LL3hDxIYYgDB48PiBL3xckkmL3RH
gUD6mTTksEL508Q3cngm9KKvOPC3TL5lSdhou0upJMr5Ngiv77t742S5vBZEkmuC
ff9PBAzVTdVKgbh8K4FwTd1KSI3PkvaH7+u9EeNLDvn5lDUFmgq9OJbqpc+1DOG/
fG4JUnN2Nr9GZGypQP2Vp0ngq4ye+kdHJPQkdcVdDHU9XJCy/wOLI6TmZyIC5Wxw
W4bR1Ypb3Wx5C0fSthPinNyrly3SzI+TO1rX61Iu4qeN1rXN1D1Kby1vae/6aDjU
itqA6EyvCTe0EG4g+Nmlh6o5YeEmtQpH5H11ScHQzppxBsBDSNo43BYciWbWyPeH
GuO1yoE9N6+L2EaUli7zbP8idstiVA7fiAYNN4J7lAyo9bTuca++ZRe/wRtBC8QX
/mzZ4MbkzDPGAtwb6Pxycp1fZk8HZGV/GRI8/MyoNu/ARNn591+o6mTNb2OXhKdP
wg25PcwIGmT1dzn/ULPbehLPifJGIzV8JOhtQkfwO4z0k0enxwOqHH44zNPMcFGA
3MACBMY8dnflr6UuHK27f6WUpYCo70KH9vi/ExxDJzR5XKw7BtwtjUETrIMPL/Rh
L3fVBcELU9gLT2jTFDUNEh8WQ9eCqYQpywrl8yeRTjxw1rIve0dQITCYOPXGhD+4
0E+/P83hCaRQaDuTaorhUyedwsxjDL70ri+PYkeUOgxYiuA9eqmuaEkU3iLcfQXM
fO8G3D5Qsvtogam4Wx7eGDVL9B6iYjJaHDIgkCWv/aUTerRQXUZUrvmcTfU9nnno
R0dbtWu8zIq0SKMFC6poU3hz4DpbWLg++E2CIgnX5tfvK6vxsgA9+tXpPLWdmCAe
ElYDg/BmooHSfyvsHrMLVi+7HJ9Wm+GJnAHu78ru8zE39Llph2rLydFVXqR8Kcmp
XKZK3HsiR+pRTBJtYU7/GhfIqRSMcsX4cfUEqRFLeX0s/47cwSSfd3LKTEtC2POL
qoAZWMNVLyNsbYTyhrdtK5RvvxX3v12U2DXff4EN99W7lbf1tsjDEWN8EtB0pS86
Q1DM1HuGjE3ahDzFgY/HaDZ6VwcXxswFRVKpt5x8IeCbGke/tOq88pulemY/2wmP
BYn3m4W74QmcnKLdx1wpRdM5Qwte+eBjruxBXgOmd8rj2+9iKayymPtzHGH7BPQm
r8m7+XAsufZC+KT3AWuN+KtsxNSiD5b1SGkjQwtznQVGKWMKHuLkdAcETNpR/A4G
aof6OfOWT+i/4WQJsxlR6LMWwkKj2AS6wF+qQiSbeGO0PV5juLoEvbny3shLJPeC
s8+roKgsmCjTTemSD5Fu6XpIykjOuBOPasI08d4St/xSfEsYV3JAR67NrKrSPaAS
ITNv7vAq+W2ghRHjMxMrJbJd8ns05o9xar35vKJ0L/7fna1xbfxRVl88GGXESVWg
6d1KnfuxVMXYg+Hjm78Z5MWUy2fQJdebNsiy8p4ENBImeyA6CD0D6ICwwSoLZ2YN
D+ygtY9IxsQTHlFWxbzMI6P/20A5CqhbuGL9twokpRrT6h4mFGiXxlCH3Pl/GAra
pE7OzC+g7kAEOKO+kvlLQ2p/KhfqWgh/JesHN+QnyjhOHcHzllVftHp4SBNLgd11
C8CZ0PBNQHlOw6YoAljAU5vK0YNuxvELE4uhKScC8vaygbaLhhcNv4O9XN7iqkMP
8pQMoq3IGd/z1iTxYTSiLkv2ntZRK0YmAfKtjTX7ZcZXxVzqpHQTL8+2vcXZy4SF
/1walcbgsXWyLvDaakm3DHyyp5oYYXLA72JvBeM0F8xb0SXLVJpXGWw/zxKdrs72
fuJlCmB7DyF03IHrPENP5RQ/qeBJLBZ4KAQn/6Uzw5EoTf08oKsZ4R1vML4/msSF
37rNNn3BLtbOjB5LybqLSMYMtTQ4BkZP1BkTHg8nFLwTOnPhdsJhen0ynGyQmkEW
qZoDXGGc4TCL8x3F5TJErzClqftTIwGn2dZqjiyTFy5FoCBwYNwpN8qjt/vjt04S
M2hOHAWUtn8M3yloeygvwIGCkIREsTJWXysLycN8VpT0+iA76QYNn9zME5LqY6Oo
GrqSKlLFimy2LSdUouQEeZhY5frOhka/HPCn8dPsNOa17Xct8B8U0TSJBlSyd4b6
0EcbQc2HzLmc279z7WihPLP8gyC+CDcwaUZIwkf/+Y1ZN8sS9CBMLkzSuUC5NFN7
3G0xzuJXcwiSqZmERYD2Y7myr0yxJj3T14+yiOmv0MwOp/8qq1YcG8mzHvLI1e6t
vZj/qHqsN3CQkQ4JUw3Fm6it/J8qRpY/XqjAS9GUvXE18vAzduhEvxsXc4yRBgUe
O/GDBdtQUq8ljnWRloZ9XUotSLznbc59j+F7cuu7e1wVhhwX7XqgFc4CvdC/zEGk
ycSX2izstorRjsX04+ODwdTwtb5I4EabJ7GB8rT3Hjs=
`pragma protect end_protected
