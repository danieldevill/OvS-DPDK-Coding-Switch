// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:04 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hPaa+5gIaAoDctf2uwhuqkVj18hI4JaqDkurf4UOA01TNO1oC5rrfjjnNTvDoKyX
y9iDiCDodiiI3iIx9AhotO8ALmw6WfCo1j5pQy5/PRcc/KJ5y0jWCoviKNIZa6Cx
NZPZmNHUVWrWd/Ribbb/Gaha95o7us8Sg0lbC4vmAho=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9632)
L7KGHuYEsLH0pOj13U/bzHTuATnbOBroynBkw+eZE5mmk9nMUjpxVbnO62Mpe8Vg
A//zqdIqMe0BxnNa2rwIShcXYq61DQJnUefNMKbl56vAB6MahX8GhjQfcdOvwMe4
py3lc18qdbZjPUI3p5CHEGT4Pz0LwnXhk15TE4gPVSmCaFbIjmVqOhRuJSfym4C+
lTWZJHgdR4jqE2Ch/qTVuiwDTdGQLe+Gm1KnhO9W1bUTSFfKETSZcmt2l5kPzJ9x
vwRn3w6Cd9FYVVyxEHLuBbtL1iU27EGSRw/JrEHn9ZTPCwrcFB7tagkKoBnTOn1e
HVSXsOFbapEa/eSTivLt2i0Ckgc8cPHYrL8j1BnZCI13q4vB84IwaL9lli3cZgrZ
bx/CY5W404cPrpHK1wuwMpqt4rN5aR4/zJdT6dGUzLPWkWY7vtg6V8fNhCy/LsCz
nTgSeMIahojMMEQYVdRyOrxWECN+D++/OpaG+svmSQ5N7c+0Ac3/RkIy7pJPjpDc
lZMs+gxOFfKj/gAoQ+75wE5kFAIxdm2mGI8YBJwTOpJ6Vx9zB6OtmHffIGxnzu7v
wnh5jkik6Q24clCx7ZFaRlsAXuK1YBRAUer3AGbu4vtDW18KwDCild2yw0FsJ9e2
0ZqgL8F59IFVVURjltPGuut7pHdGxr7GdgGKSxcylZ/8SvH5bQ6hQ1WYCys8Rmfv
Svvn+8IWwTOTuySpOKT4j3Dzf9kvNNXVFGS56UMbeEneBwAzcdunBy5pqr0C6ohM
8T8+yGf/6yvPAouXfhdvGM9J276PGzNm0ARcXZrJjZSo/y73iRPP46DGrNWPU8YX
U5paDP9En1JXgx6bCBwPHtJs+YgoQdf1hxB588diM37GCpwTP8P2fv61MN08/gD4
YgbVerwyzInKBZG7k8DcpkG2QfLEHXW1vR135kdjuBIHpfF3nAmCg4mcHBVvnXpY
27rs74kx7I4zbtSMxxjZs1nWT0MkCD657pZgTjHpB8Fo4Mi9hZ8/Xsyjhy3M7mEQ
269ERNY1q6ttjcJ57afnLkDFS6qt6vq+Z+tRwoeLV3Uu/hP5nvvEWHbEf25xVDvO
+VwNYrGdQwbijGW8gi7X/Lq9dcOjgYiTQo06Nttuhlx0Xwovjk9XrtWwGcelf3sy
+lVMHtxo6/+eLwfiyF9n0L31igcsg9/R/A94FhA+M9vSFiummpLRmHlCCK/NW/O+
0NiS4JvM+cKm3GPi/2y1zVPAt+WG/U8HEchJbtMN9dw+ti35YdnOwt3NF6EnsrSy
16HiVlCkGmrOzajGvZqSvkf+IJ32rvrWwj07W93JaC3QAqoBLprt1g/638jGeq+A
haJQH5SEtwdo4kY3Ncg6FKsyfPzQDMK61HQ0RSo4v0G2NlAK7TwgiAAyP0N4vq/A
r6v6WtXN+mhU5y26uRBl75IkehmQ1sWpSt9f/8TzyCHuuPcP9PLe4NTNB0W2Ijiq
MESNBX2Lf/Oigo+T8WBJKv3wrlM5ETU2lAPW3H4LH+AggQNF86tpkiE5DfmT7ki8
8liCiNDtq5Bj8vf3X+itBvP+22LTGLb6cH4xIsCCKPuDvxW9iPq4rx1v+5/IeDNJ
ClcNbyL4immMhMD0/v/PZVpyjE4bpLqesqdSbKP7ieIz5IiZ5zQEVL39sLNzim7I
aAU/JlerER8D08q2bAPphLVLYEC0pFD/LViRgy0P3fu2lsHnfMTimTwCbmSmqnEf
/M1EYDBAAUJXUb6MTu8r2hjqknAgU3sqYbK9HKgAx0o50/lZUGp0StdAm3Avpd+z
YX4AxCaAbUn73FogsvPXn343wV3OciPBrAujzvEGErCBjbBhv3GP78ZuRrPVofiC
m44akztBwhSSjXwoGpZvM58+uA3xAmUX12GmVO2GOtmOzu+w6EQzbAKVhY1badF5
pMLL/GANqxQ5rnBVy4xcz4atnQ+aRXOBPkPzvLrAcIsANMszUh5oTV6a5/5kbpmX
XfCwI8ixJ53rphaUSstNR4z31akCiKu47FU1gIM+KIsz8BJsmIhljIJQKJOTQsTu
kfeUdnx8Zg+Xiyz/xaqG2iJpsM5p6OnhGxe2Syd9KX1xISBkFw8aL+EylkuZVU6L
BaXhaCnzuCvpg+64Ad6amsq50fVHbg6mZewOhbW/kLuaokSJM2Mfvr7eDZeEa05K
pECVtXvsffMxsH3OdKBN/0YB83Gd/uUKf8HFvb6WFU95nl04xXPP9SY/ps5HFvr2
gn59Vf5NtLZrwKxFaiNdzPct2C7TXw41I3F/lIpodkoVFxmpZzzR6AylAevzO1tt
0tQJeOmZRJR/vXnLNsoJzsPaNlKcB3KxuAtl7qz5S+XrC4fllKW90IcgRJ4t80Nl
xveURYB3LqleyKbK9VUCkfN0sWXLxoHZSDzushArpF5ZNKSKjG/2h3Nx3EjplcLw
wZUCW28PH6KIVwxaSNs7bETUlGOwfooigVYq3UMsB0//P8ecYh0N9Ebb8sK66W3Y
Pw28ITkYl/dOZ0gaNXuAFZkHqZJg6zuA1ei6uEbh/JPLQwTu4YSJ0WipIx2+6qK0
uTQNKI4be/s9dX6NlvIormOgFB9DEoLNWIBdYuzD46B85qapUs7l6f2GF8CAZkDQ
BiPygsE6D09FY2EKxbtaLLuk/F9HewY9tWUzZ5Yp0qOvJOIH9JSxsMwfWFIkbaCf
6kQZ+du5xIB/jK+OVzK2BmE/ODmyVUn95se1v2r51VsRAhLs5gAeVOxxplMwUTgl
cPJsdoiJ5+rHyqi4R+rv4oL8qaRRzqnpXUNODSGyphkZ2h7gRCjAbbDxuCLNErAz
1g2vqVPUAWFtbGX+iPLvHlyQtCK6Ai+69xq+WC/OudvN7VDcDuUZqwoTziq2vXQe
TKbh6RUJgpTIicMwjK6bnjkK2UhWNOekF2ImSN7P5oMWQyfG7ZWOmUT1GnHj7+J5
V9CgvWFZwjL2RzG+QWvIa11LAHrs0PgUFMJRTBgDHGo6SClpQiNEDP3OVQRYLsg3
+PWblQ671HDRaGuOBgJSBMNvZp0FGaAyBLWRT5GlSAbDBASvFYaPEviATs5/mqH8
HqRUDqOpXepn+N9zhX3xORh/suC22zCyd04nNt9NjNXtX+NvKcVTqj5L33V53S9b
E5IuLaZPM+HE4LyPUz0znugq9Xe6z125TN3P/CmTtxGnC8Vxbs1eHFlpyje6lKic
0voqyqZAaj4YOnG8n+qwa82vBHL4oWJn2xsw23/iwDUcxOiQuLsKprG/iS0Dfrds
SHXTAAs/JmAmxWD84dbowSf97wKx16WOHr5CSd6Hp8pl6XPKtGkL3YNLzOayo46M
MZKjtZ3l2vHJ/b9LVCRtPL8yw4yRRU70CnC2Gw/XHxM+vpLDxfr2pvxr+HedqV5M
5LwjTxZE+1wAerxPKh49wk9N7tbkD4zZhxJoW+GU6jlW9eJtFW9CKuB6umsp+WcI
2oNuiHZkINll0f5km01ms9DW+0R37v/7C/lJgjejBq2V4AsnAgCn5+nNGH1Uffc0
jxD9uJYLkNMR2Qz54lvm925ZtzzRt2ZUudtjIdG8xUWMTHQqAxX7N7KzHeQYtw1w
tCi9l1cOg/qChS2NNDTQLehBj4j+I0krauPW/dHTkK4ePSzR96LSk57+FvYdMAgA
wV/TZsi7Tx8y2XXxqDDwTedBLtwvQ6ugR1lYKirBwVkd6sAvXiaiYtI2aVIsEuIF
jdA7b6kVZ/LuaCDZAN8NucSxkfR0djWiqnQdlsPCqDlryNK2uJqervmcd0ILmOPd
bmXhLg8ENOLy3+hAuTXEx9MmEvXDt3Q3AvG9vFDe5psVeRN1V8QYf5jYq6VNoGn8
JhcTEjgVNkCKVVhmWj6+c3iJvCpV5nu1lCn177Th0NCiIxsyTC/vvZKoAdrTnoDa
DAeo5NHI2He6hQUVhlA2GfkdyLaC4iMiXqQ+WL52ngMD3wDvr7vdiD11cgwdp/mc
fYStPKGSpCElGN7YOsck4EGnfIgSKRi9e2cddax8M4QY1Dc7am7K9zNnKmoS8uNu
yODBkRhz1Rp0sb+Kft8TV2cxbNsVLpqAI4XjgHDDqRPWncRe2B2M/XJVzeBNgJov
1ZvJOTtZF8hJzU4L7iMzSmH3N9CzruqxormNwvn7yrj2Gz8mHQFUU3vLIwGRCdfp
QBjOmZ6/Th3tHxsSkSK6GrWMS8imQcLsCRpdqWjDm8Wua4k2380i+N4CnOATspZ8
POAg9coA1gtr/wQtu3vBsAbiSRQdKbd4UfGqoH1YKeH2nzDf8NSnoaoUb5XE0gyb
TTTW5vgzItZTPhl8KVmAwhp8+GXW/J8iPQyYru9oyPsGxAG7QF37a0BfzVz9TEit
ZwJfn7BzP9Xk30a7+JyYxjSKYHBQQ5gjyFDEFoxtemuA3FZwUw7J/D/4Hn/i/AXZ
n1mk5ihQmeI81OIr4xnoMqYuBnpbz2HzyE5U2iB5iRSZl51sk9u9KIWzhPKkA5cj
yM4w+z3w7vpbtiQKpSnct4NrV7pQHDqyuVlqBFkPsn5ITepmv6MD6eACCM/+6VKZ
OtgxAjDF06ljFTJrfZpFQBzTwD03ldMmjIjnEY6PI30njHg/XnQ3SQ4fzlR7R1W/
4c8RR+OhTgdAPbEQDAAJxKXHXekU2HSfNCQy/NEvWlOaC4Je4HgW7sANe4tNG2BZ
VbYx/Ym3eUlTE6sqz/eBW6MtH7541Rf7tfYyQK4BzOxkMwjEmiPH8AcPaIXeEpCz
RlnVMPoqti9qd3ykbbzQ269V0WXP06L5JwwNfezl+oobRSMwP/zcdNDLo1uITdmp
8Re5YN6VPRIkeksclXF/8rVwTMpwYI4HaPWly/87iSELJBWn3bo8U52wGQck31ip
dymuigjwAdemJzPWaq1AIguKCqEH7ABQOC7BzSINz5p8wl2SZYRkZAZ7n9DAZmqu
QPTVcs2P5/aLmmtCxy4i6EA2Arxpfm76CKLXGbucbRDu6ORyID6vDqIkasJN85PW
LNLdU5aLAPl3XlyKFY+iyDq4KWyST8iRfmyQl9H/Ezb0e08xPkDM9D5oYOBOrwW5
SOj/5pzDo/8YUc13OPIJsie+h1Bi8yHy8KX8mKKtI8r8E3GQ1cH81P6lnmGei4sZ
mbO0wfxwYUcWMTMocCeXPGectUHG6WCNT9dZE5/I9PlCHnhggtaweOjJ29zoHAFA
0kfSTTBhbZoIlhnDnZxBFAbva2d6Fj1Otg+ENKI8Uz/aYA71RkjiEd7vwTWaPBzf
JhWtFi/ecdqgem7JuLN9i/L3ik1vUIMaT/SIJQ7o8mwQCkmKmLwF3s93DOsXm7VR
yXRtmjPNy6p8sy/8+/PVWMKZTbPU2SSAEUJKE5nLGzV1Pd8/ajv5ouVYopmK7816
I8RFESmIQ3H+FdyKOWeHKnOYkAleI8mwqBGnro6X37R7oqv0nxSDKH4nuHPB+c5/
8k0BvnWI6SaDq98NpWjuaO90vvGQsi//52LIUx7mWo+FZ6tC+ArxFH8enyhqNN3t
bUGHIzRC0CtMaBoNkXcM/TQf3aoVxf0SmqIx6anaSMpMmXIh+3xhvVn4fw4WuGDh
0+H6NzzWTn6PZAQ+bZk/qhxOLNr5eGhBIdEcojd7JhK82vMWXENoaL2gcqi0Z+64
Lmhe4MBskuGZKKotS5wZtEWkmVStu8Cgt4i8Y950Asoa9bL4ulsjyz7gHrwPQuGF
rjqMRr780S2qLXMZ2Du9RoIY2dypr0bPHAQd97fA3+G6kjWL9SS5rLd+EO3FdYIA
Z5cd8brVoWK19EtnnDMKJt0xRe6THUmkaR8VlaSeC5A4q5afTy+AdHHXG/R2OiO8
jum9ULfUaoAt2QqJAVvvC4eeCUI3iDbzfwXI6QjDzzVmuF5Omlle/a7wYM7gIMqL
UOZD3XHfxxXqyACnR8GIEWhGVOby75x6VQsK3rRREuDXM7X16a6KeRxJs088yBQZ
+ai7Wg/aOUCCat2sVfWs56+1DBcb8q1RJC0Id+LqObSzNoIrU+C9e8IkzUl7wPYn
naDcHj8ZXD4rMuqjIclq+53Fh5zd0prB82y2bVnubsOnYJYMLZs9bwYe8v0TaxhU
QxIUZZQHGw+Bqv+3ybQbZb5fcKaVGpRTWDQ5D+hTWl2iFQzeJhbZbNbhYR/5REin
oXIyMYgcL/3WkEROLKx4svkO9vY7yZrz4ezxVFBoKbddt8QuVfdRo5AupAvkrkeW
NrOCIxd5ngTVwSp6MMWAh/gRORr9e4sMjMvERqllz0ZIMSotfUE2VqNSWO1nI+Su
qOU5mWKsBz/yoq0muWJEhwo7R4Bpthaox/m8zm+q6gjJ1Ze/7NswBmEwLA5KX1XT
Zi9sEsVOgCyZMiLja2cNx01ALKoPhfQwxIdtlDOASRwnWmKi4aBq7OfARvP3UG4y
KxKXr5Sx0Jj/msX+L1OvEFOlcHjo+S2bVXxDQSLqKTAlm+yTeIO7i8tmxRCScbJL
smJbLCETDkiX2qQGy9FhiV4krim3WxpLTdEz5oEmcTi8/7GCx5rXOEl7ebC7tNp3
OMuADyYDMslSv/yhuy8zDAGPXk/cMO2yEV9ydBugUvvlKcZPOm6JR/BEGPpUy0sT
6CofVo/XZJ5YhksNg+ntHVxD2zXA9hTk99EYZCoTdPkc3QDRMAhxIAOPlC2otb4S
tbsRe8aSTXOziCMtD9SNsEkdQet/4P3vA0RdGJ3RK2GnNrtn217vcC4b+Wjbu2Ay
iLOTQLXybrmPouOIZFrIk9JgKiyb5jTQRG8nJcLxDdVromfwkQiH/fReKmcNh1f+
7XfmuzA4+/pkygZ+Vwx24tQKfW0KI38WYaa3Wypjdp3BiEVvAFVQ46BF541paj6F
+erZCZP/sQEF1lCRcrjHmfM+uaxc5Aq7x1zpLDs/fmTLPZEYUlUR5ZZbAzGkwFUG
C+Yf7Ghgoxy697p3jpAQP31m/C5xecNrmmG7rlVRwx+UGDx1+iwrV0to2pSpDY1m
J2WCukNHG+HpDD7i1Hnb0DQszYzSWBbYl0BBiatX0fl4brt119091twmG4Vptlhy
5YAOPIJIBgnV/AcMEqOeHernDOVWwWZ5apkjkrK++QbV+8rN4HWLZ4hvxbiBQS1d
HC8g/JyNqLWkMC3T8FbjQAi4wnIY8hAd1dDb691VMATZEM3FCUkNaONpG2EEP36b
/Pzt/qI/dot2eQyM5THyAy02Q9DsfEIQRNJ9pMjQS4SGRXF6F+M7S9njBkZj0guS
mpBNvwHU19lgADL5hLmjDbcd6vB7BTluH6SJfmjyHixE2cvgqsqojvZ9ROwCXNkj
zWlfCg6PG/X/2fvNa8q1pOmMje/eO0+4gJZ55lkKEwtXH5W3y9jK0wv8eh4kcIyd
2he+q2ijDcazmHbZlB+4Y7MYFbYXEu8yZLt4YGoYI/OpucVZLRrS4I9F9BkPG6M9
fmh3aYewn118edyvOTj994+bslvMm4DpL/4/YcLSyyXTMtjNG1EKicjq4IKiauC2
Vq6FbzJohDH0xrSEMpXlvixW5iGYu6NS/5u634hJFC1HhEv74OexRfb6erEzYJzY
bE80gTuFinN2/GnLZO/0/YkKUwJZROD5OgWNSkmRd64TC1l7Auv30WgqMrRPTFSF
SBKr3+jMvpBLuGn1Uztu0gUcUV6AkQkekRD1smyeSW13oSY0rpMBKDIyIPVxdHKU
MV2nHvXBsuiYsafD4vk/7bIIONx3eER82t/h3Ukh/drAhrv6D5xKFh4a/Q5JeF8H
5Ze3pL8Gf9SzqoO1aji1cPdKJvCud4C6ZQfsZAH60Lp8IB2F84NDgXQyIntIJ7Ew
M44ZDlYQ1H0WCM2wwOJKm9Fn5n1vPaCXog8A372t73TUvFbIanOqb/CL5n8AEete
AIRptUgTEzJXbLV+IT19+aPPH72Cl86C7MjRoLojFxuRQR3KS18cX7exkKXiUahm
v1tGngr/bmXTo/zwP2aKpnd0eVkpjTMaPtO2elr58c0+VuVwQewUFRAdzmJ+kjPQ
rTZNcE3FeF0qhfI71qiXvXwumclHopIf5rmMBvFTRL27XZwUtKqqfEJB8Rz+tfx/
r8j3fzaAGjgoKQaQx2AoATziXUdJLoJ+EKwOtZra68m5dnemwjNlFhObgj92nPhQ
6jIshJ4tneXEX20USScYacO0si0pa4lI2UCEJSqnz9glnD2LYYN6oiEMw+oac+76
dWaNTa6Ok8sxcNgl0Zz0otB7j2BAJ5oalEmyRHR7T/0noSKyP0pbddv5RhSTtJZ2
iRqeEz/oOVS+6dNEgD1ALe+rc8nhBm/y8XpeFaiFwoi7zW98KDZ0I3oSg5ZRjT2B
uOzsC27DSaY/B8n3CEqCvh8lbBdZW+6hK1dAd5Zs6gcgeWVPXs2cCup/jHfGhqFM
K6AnM2HfHkSHq+ad/scvHT7w6s3vCUg+++81OIgY+suCG36aEICE5kAYW1PqNwMk
dlnvvHd4SMycDEKyqILPfROQzmCS7gHpPupGA3SPeLJ25Znh0rMVXvgxsfO4aA2t
Rvjeqy32C36PhoVkBU1uFUzgw1FI1PM/0rXA+uoQQzp04R/PcWCzERgeWwrboxaL
M0matnJYkFNl0k7NEvlc0SDPkqaClvCOPOZJlKh1ZVrIuCKTsUyVJSJOcgmPoTlA
+SyDz4oBgeo/UvVcT3Aaou1jGuU006ronTK0lZ2vYDKYvWA+F8LbMq7FqFmDurPL
yVbYasi1c3Hp3gJFIm/OVZyAwNUtVukq0chMQlwbBJf47RArgMs+Z4aWj+sCJeAZ
ZkrcXZ/ko/NyuvE+xTxolfKCntkGMh19PvPQw2vqsB33zmODg7E1AGybLPQqIZMC
ttvm/kxz51D6quyzHr1Xmnt7CTR40WSA/Gz8ArqsRrCfl5nuXodlseEW5tcwMNul
YUt+BLWoLq+YVsAk8BncQHDX9R2Z37OVObKEUFVCAyStfLLrRpjhVPfVwWH7Mq4u
+4Ns2lgh505MqdFGzlpLIxkLiDH3IMkmITxqOdXAkIp37AAtQBVoFe+5vGJPFwBH
QbfMNSn5KeRqhjSepVfWg6vEIfXxvBTQUhAPIRgPjPNAmx6lZdmk0v1uVwJ3QERB
bqnFVyaHbno1Y8kh/qiN28IidgKfATHjY56ag5Sy1v8cOtK8S3sXCRpTVuKyLHYr
KciBqpAV7UBf3iwEnP/1FqLYEgUw/c9RfRRyInR4ReWnWUxS9qfhBHrwc71nd1RR
2ZwawKcHAXG7dM/yYzz02tyMyyR3Ma/c+woHbv3KDPEYHrg6G6NqHaK4NgM8ygPJ
2zRIAvs1k0xBDUDv6B+XxAqsCKX2t3DNUXGr8tq3f+hzgFqoHcZTwzWTU4J8fUuY
pUeS7xdY/XhcB0qqtbCkzPPbR0IVBPZrEgCb7Unzb61bFv5S7I+vm5AurC5JRrQB
wtY9Vem+FaxgwebYeMPemq35D3y+am8cvz0RuH411iP2vUS/8fCVPIbC07d6H7lF
H55ycSXhI0pCoFB8HvuWpB98nQiFZeCuWbwljdEWYxBiO8oCWyiFeKDVnLnjRFvV
vT+rX4r7hcDPhTQUURhne+grtli6z3PbgfLpyzUxUzPsRoESO5l4741Kp1ZUOAyi
6rb48BSrLkzsUDiEb/6sLNCrcREGMS/JxA8mNBcCk11VnJkly+K7juWDQFqMgtc7
t+OoSN2bOTm8OgpYFf/KfkDqCEZkT/TSpUqtURau3E3m7JBuGF8kFEU1aIw0PnhG
V1OuVeyCFJrYuHHUu4+T/MoR+bVCxYQtecuQYqmbEGzgdTNbHEh0qsg3xVNHLp7W
xB0JmlyC6v00FO1rQ+kVXktp55EVAj88AFjstyx7x/mB7RTjy8sLxrTISJzKMnFf
T9/lSfMSxOg8IHj0/DSvy//yye2I9IncxN5JDIRnjluxwpTtEKBrNpx1MIMPBgtz
gh+Y5HTNVa3POejz/ru8eqVprMBuyF3iYzqERO7P8NOAl6d5BRc2bWPrVRWjEmqo
WixdTjSVn6qqwgvJEvNXG04mnk8lFlOijzAyI9aT/t/1qvyk3GFdw5zlaU5FndaF
EPf6giznYKINOZ85lbWyDC/HAugnomCbAj51EVDgNrhazCPaHP7FWJRE2mGVV1Lr
xdLN96xf7qqhGQ3IfPo0WzJWcEk8OWCvkGU98U89IpVQnF6kcq0UDT8nTuA/nk+k
0XHkq/15u/BbnYuqiHjVBsJLrApz/kezTFY1n79tY3ASBOHyPKkZITG9V49NE67n
hWbbgkB5O+oi06hwwdAQ0eO74pWp28lfE4Klopf5/30oI0KlekabW5KWtCs/31Pi
66f5LNGBlpMjDnZ8Gr2DgMNUOeuC9550VkXGsIebu9+fx0/iCzr0GGSCW2c4llEP
9l4WThNKQBuz41W2iBlfAJh3Z9orB0K1u39JjAQAfbnwRamfS6eC985cyCh6PFBH
GOkG5LQZlkjnR005aE9AsCKyCm7CZijLEWE7fvOSgzFJLnv8oPrF37JMmhJky22u
S6apLzwTs+PGfng5D80S6tbvQtJpf8XadNDW02/KWDJn1UlLFATNUTWjL55p+DXg
eznhSLxQSlcC2EMuRm+LeM+X1BhqKe1zNwrojcbE4bKboOfubOIgl5O4Q59GvudD
Bcc5uAWOhiZRKdK5/oWEKBOS0voeFfWoh6I1ZN6SDoqZMKzqCe5Pg+BhhLikQoO3
d1MsJQBmYvVM++0YpKJEbw0B7+5VlX+e6JPi8IPVGsujSc5aBFcgKMJflip63rvi
mJZ1N+vP7JNAFAMXDQVTlWmnfMmwXAX6XtP5ayDP+o9E9OHgU1E710E0/oic+C91
KeMaZYdXeGapg+RpP86i5Bdk4PBWd6gPTH9Q+x8ChvCh/qoxG+sJKhoaQeJ1jSQI
4eOnytKYSCY2NkJtQKtYoZ1TKKq1Xl1shjoOWC1mR0n3XaUIz6KHmjQePAarnWey
o0Ilq8/ksS5vADTvAWvK8hjvTdl5eWUVb8Qn5c01PWgJF0XAIhloiPKxzo1INAVC
Xq2kqklINdALs6DHlbyF5d9xUIpemtwQfNlFlNPq4UmRxxDaGA6HcgXVFZwkMh09
E3/Ex3F/CgAskW9BjIzqOOFf5Vqr+DLnLyZLQUpAo2u2k0AJTBYSU2xGV0gebAMw
VNp7s4sHPhLzpL0sd/UCZW6PA067GssuNsexNPE582VXSJGcdh4RNKYoSxVnP6jP
uYiO8TWVRr5XGt4TyfWXCnjsImO2C5/PvBaQL0YWxzNIZpJR8mT9Fu/ijXPeZTDW
AcJT1j7AhoXiaQslGhYxbUra46lHVbY+AoNPYwzZTZt1jx265iIdROTiEeRjH+LC
Mz0wetRnDcQ619zsU81FqMfROc5I7ny/UTOrPXu2t1E1xG5NkatrWVhUE9jpLGrH
CQ4GZobgzUGKFMhjuEw87IXraSxIhg8I/4UnHiRDtkOwJGT0DCx3wvebYGO2h9CB
ImrpVJazTKRasc1lNUhEKJMTJFfv53Nr9EchoVc7/0sm9t6u7PeEmWZhqV5J5pjz
wch0udHgW/yipO6SFvQc9/4fyV2PGmKMlOD2u1Cf4A8YaPWaDGgJOpD95qFqkV9O
k0msUSfJ/MiJtgbJo8WHDDdsabkDaM1PsgpDz0IJKqBzRe8MS8g1s/1CDMxillOP
TjDpIebGAMNPboJeHEb6zLmpsBPBQ8FvpcKdsfrAo+qVzQapE4uowmjz0L+kjb7w
SskD5BP0tskVdZmm14JqLYSoZ8ZCHgA2CqW9S0wx3jAC7G6TUTqKQs9nUyor+79x
OQRR1XhEk3VP6dA2WkyWIkmF+3eGtKg93qIQ2hBZ1SqWOyveuguRhoMEbKJdCv+j
nsmrCy4sihmQ/20E1ce/c/ZCiUfVtpMLV0h1GzXhplcsuT/AKjPANHI92omyhC3b
Ebf3lwl1d8GdUkRUxs88VJSrdGMXNsCAjwfvSZYh53u4bp1eu3WL8RgUomkrueMh
uaTR3WcCPg9wJSLqcQ5dvuuDVAKhFpJR1+BbY0aM0E5HU7OcnjSMj6TxXgDSnAN0
Zj4lZk1s8gSyy13bFJFGdiI2wbUmBJj6hE+TrEEJE/8DeX7nzDmWcGkjZxI/vQkc
pI+pgU0lEFVIxrVKaZhiA9D53ei4ZRgniy6AGqux7HMnaVkUryNrast4SRqkIm+A
IJtnZ6oyuM81x7A1X+FiZjTFc8xLIubEzKgTU3tnUI60jBkAWFpSc3PNlS9BfOV+
eo2cdTyKxe4ecb71IcGtqp2VLbaaWYSVxSCTRJPnEsgeRlH6FTEqP/1h4Uv6BP7v
8AOoS31kvU311IteNh98aljxEV3XTU9YKo1fzr/EVrGrtlInrA8xi+LI3UmvEtO0
WbRUg1YygBFuvTUjmqtnc2C+IvsIPz0peDJNALH5E3ja77j/dcHuLSf6n616KWsa
bKloLIlJLrZBTRK9j70CsF/IuxEDSVZu8skY/HPCM8dD0ifNRAuLbpBPwEuuaRLd
eXLRcssi8ijbEofeGkQsiD7ZRK+ZDqQ1zEqu/5835epeYrRPnOn4rBtlhTaKEFra
P70whM/c1otb9mR2hAvwCT/tNdV0fW+YwOnN4mT1PN42zkSpoNbqualV8jdNYz1Q
xHMhwjV7M5aSYrQR+vu3LMg4BVfUlq7mDwPLp0gcolzoRK3Y2eLSxpohZCPHYsoh
Bqxs2nuLqrTRtKdSB4JkqDHCo6hs3jsgWHHmklD6Kgk+O7KgjXaqEZL2BM1pBxhS
7x813N7rIfFmJClNeNPmu7fLf0ulU+UfdvrRrLCqGIzJpZSqpgaFeVRxFmFU9SBK
rwPulUVA3J0ZKgCo74K/ia0uZ8iQYpwfWsY5EmE7wm8=
`pragma protect end_protected
