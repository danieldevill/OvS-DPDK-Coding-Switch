// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:34:47 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fdznsgHg2IsZn+1eHVjLqmuUsD8G+ZF+TIWZWreNK7xnw3KMSOQ9jWQtK2oDMaJl
JFzqdLr0/IEUNrXyYlIc5244KJJQW2qF5tjNa6dpCIQ1TiuAtfVVwJS0hIViiu8j
IXeAisHV5dYiWC0ZMW4YLG5nae59uA7gsyYEmWMeAMw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11152)
fY0HS4oBlZe0dbc5ICdZ6hHaRKwfQRe6cVtRCq5i31r9y5fVttMipsCnu7WuwdDc
Sj3/N8zVfKo0SZYE6OoBqVrwrJEnnmRbhaJi9qDc3hMCgBSoAET2VVar9hrFtTOk
UXgNa30iAYiK8cC3s1lF2bU3VKUiDeRkA4YsRMmjjuIIgHZOKw8J7Ukq6gFN/t4V
JRIjtWLXnejtSayXdXarXBo2Npyk84PJAWTq2JeXnJpPQkrw5gDAus5KnJg37gLM
zMPpGYFk/vspQL71ulsApFkIK3rX/dcSG4d4UwJB5xGrlkgTgj7Jq0cOQZpbZCqo
YEaqdXOc9zj0qKIKvtHbhuleDlsTAd3RxtTC6guFKcEW4KPTQcEZgegi+zYIJkX4
LpqWDaltkyC3MCBqrxJt6vG+MQmlVcREzt0SIO3FkwlWvLHwPOjiFcB6+wq1vxcE
rgsrHBzcmeRYwMGPzDoLoXNU36htf5mbS2f/tW/+Db98LgEPvBIxl5045oAwpDEQ
P1loRokgeEaHaoc98B6oh0bQ5t1UMWhPiiKR4Dfj8SYkuKZKC2jwNLQ1Q4xIxfnG
igb0FFBDO6wcF3MXYQ6qctWUFlaZ4sCWETg8Y9hwqrhg5m2dc37gSHzoQPme2+cQ
fZvhB6xueCDUAorQUpR7eBHutMcj/XtNNKFe6uWmqhjLkKJlh1/aDBArL+mYFqM2
HmWJomqrV9Xr4Lt4uH2Irr/0ZKsuocBxmC8Wu2Ka7KlUTv457ha5/QRK4EbVPbmb
Lo72DcS5zIurxmtHctY0xMsfhRS5HUtOARwkus45zBQT9V05B5bMgOcFhB5KfLiv
Px4GlGVehWN70UCs6iT1/FHnoRKHRySshSkf6ispMuZAVWZp3NXcMq7BO/LlfOmY
5KswQRDR6pCq7UpEP2WjhVHE81hZFDgZw36dRvgZ2i4guQzXjoBxNTKf3011Erdh
Prm5hRuSOglN4uVkGonxSl6D+cfYFOnLZ6DK5RMwiYFBOKFtCrZd85C+MV2T1eym
TWWAzxlhHe/z7H4i8DkFpalH17RLG2Sbj75fJP0tA2lNKTlW1y6MvbBAz8E08IBj
MvDqj8ZQ+iMMax96iNw2Sxl3tkRCQ6fKn5dYcez4XBBDUS7BYLOXsOkCyBdbLyXH
dMWauwMqbjeUKECImaYBMWZWOtk1u2nz1CGLrzwzKg3GLc0ir6A8SHMZ0recqpMz
uIZwGIqsyVDzWfLkEBov6JJ0loAXaHnfmmhMu0y/dhFipbh66duMgcTDd1YaQaob
SCHiD+ZMAuIt2ivImrrM36fPlxNT6DnhWoFHYwdhb7CKEATxjgTW9InOmPbjQ3eL
d5NsEUK/h+ksRLMYSF9+rEOH2XTHg5e7C4BDF/7jyTWXdxlzGi9UosoWznuohZSV
RQCnSkciFXdv0xPS8JECawFW827HuojIfJk1pyhaT3ATJPJJhVZ7Xi5UE7ujgdPO
Og7+Ay6uPr9pVgNwR1G0Ru+vSDuvmvQz+Q/iEqjn/BbsgwfX/2Qfa/rMEEN2F44V
xJvDK01WVURkDRhlmkNYWfZcDe7t0wGgwnTJM+PR4YmK07DGqcNaOh7yuzF5J0PB
GSB/ZMUoOempFsjvpbwd0C5DCXvfJBqy8ULKNd1m/eHh7V4zw/H6DAj0+5P/mBBo
DH2e84aPqXTs2KDQGembx/Py9fOA202jWdIlnQ/VvvaxjNMR9HBv5R4BupMi1wNZ
moh6ZNyjcNsnPTXhgcyo7YQ5md22d7sMLhrvcaaf6mEUN2wrClMFrua7Xw3QBznM
vHzYxMDw0w1XrB9viH3KlRiYJvy2W8n9WFjbg+W2CZ35uezJsQkytoHFPj8Sa0iF
arBJsjQN8RjQSt5c6/aLpoS0W1rJ1eBCQQhyQv2wtn3hxM/MJbkmg0ONuEl61c7y
mSqZgGf17qv8O6cJY/K9RzL2OPSkSZ4t4qUWHul+FcfGMpnvUmKmpdS8Avkva3Q4
wKfKQH/b9nhL/fbab4eI0aqTbIe6MSsH2m89JdBfols3rVTZ5t/MkEcfSH0X5a+G
3duVtWlu8XRscYhC0kI9J/WLLTrOfVPH09x2r8i4S1vs8I+W9aZXX/Zuf6ld9Slf
Ju5eVsrNM+nr6qhCI6wAOYr0kwvZXc92fGRPB2ca2OdNAwVbRRLyKGQt6Jc6ANie
pM/P7XL4j1sY8viKWcTDYTRbuE1Qyv+5nFSWh+TLuMM1LXke70uAvwh2rhD+GFkX
285wrhx1eCy9m5yZPsOGnFG5tftvLspUR4LvzsVhxeukg1wm69KmWcLYynmWu8n/
Kuo9xaIpKDOYKZPpCX8fMPTT0FZ1R8Z71/kBibUlBcxLKa5N7TVBPZBAOKZadExk
sRh+qRNhO49LMKKazB0PfQazTvlLtio5u9GlmtIcwpWc8e5SRqktUMUUa2RBHwb2
JJq1mDgf7uNjayREwxXZzeXiVmtwwGpxbhWdeTbP6tf+Uqv9b5RBMi9vJgbq1U/G
9Wdin+indbCQKLWII765o2JxFfOw0eLgtb98TkRbyfwH1pYBcyynQ7Ge6ZRrzoFb
RKmBxCA8E966n2L8l1cTyEhFn6ijzurzDoHrH5FqyFr5zx2ocJXmkghVVVdAOpcO
mbRwvDTtwb8oeuCVFZZfS9TfimUYZe9z6oHSPeqKHpWf+HFD0eLfPQgY8akNhWjF
6xf/YadrLvv4IaYbWhzrIm5dOSG4uhf2AfUDaCtHYchcHDOdENL3tALZ9C5Bv/H9
Xiq4+zWwKsC+QVtRw9JHGIGkQI2W4GR1eKzezGcA8y46qJV4+WLTh378iQKWmCCu
dm01OF+dSBN8lmxJgQAwwvJ4xO28JsmX52KqZSFGygXhUNBwqBfoZ8CAAgfcooKU
MQbmOJIjl/QCkv0ew3OmP1KGtGXj/C8Vv7DJb/Xt4p3BKb9bKDKguO4X5Igni10Z
3m6ayfL5VNzezZtBLaPy7qBMthS14Rz4DPWXaCQKoVpeRTv5NzwsSy34KLYStEWY
Ml5QsnmHzWRk1/NG7JCeNzNsmyO140w9ffFybYjWjtc0U0MrR4Xue8XZIoqi8iXs
p07WuuZmSMS2ITpygmrnM69oikw1LAqproa1EbEdfIs6gGB//k2sGmbbiSTXl9b2
8hlCXgvnRxO4etdGMIOSiEnfeLiGjwOCOOiT3AqW+sdWplvBojVF2ksWELgEqBZ4
lZ6o6PBqRRV6eSxCs00Mjr0rrkPw+t3JrE3uf7Zsz/YpHWjjScBrhbbtdcbN9p2M
iTlofU2usj0Ld1qN+H9c4tcllhQ9auzgzRlw6FQo+7En6MqRRzxSe91grtazNHZU
azimc+vYf9NHNuAPkUmL76NV9UGAceKAEyPL3ueXjN24jLzHy3+TbyNXM6DE7qgB
Oo48krs5Viy0h3fUak9kA8insShLQO82AhYRzgPVfnTcbai147lN2Z3/mdCCeY5c
1cjKqO6wLqLFeAR3PhbXpctG0zvMysQDC11weTRtdxOPHllBXOZh8sTAJf8h6kab
SNNCVcDkAeCeJ7Bz8DERWOTdEY2/LFE5v7C6l+NHyOtkpq6m40tCnCkx1w5NJ+qo
1vCK4IoAfeazJJDF2YqwoeGJgGruWnKT7Wh3AhXPrvTxkk8upFE8T0MEK1xnc03a
ZXuP7F1dlrDX2vdInoQhefKtC7KAaAmMqWKRUTgXQTFdFp8qax8whyi82hgs1QX4
yL3qmvFEehDHmj1/QnISE/xcB9jq/zK60mCRo8cWqKtLq3fTuAtcMBRswaFk6ov8
0Oakb2vtYciD5YqPlIPwVXDNmsgWTT7t02XxB20NKECgR2qr7vCjjELJbdMqQxHl
iraBcIl1RQl4WjbGXus8r4amM+CasKuQgg4+Dsk6LTdDYVv6ACaguSGzE/xHFPi6
dGzWQ0vyL3tpmrDSTc/P4KNbqtN4Z2B16/WU41FcdqwGq8HciRHTn8NbHfDkhZso
igj0iSmxu63DHsPrJa26tqben5fr8xIZnm1A8Na9HBD59DLNhHl3gqVzq9HM5C6R
lPgNh+tCuUFHTKt8rFwxhr3GQt/Be7Q1+eDmCudjnY4lsn7bFshFoBd+RPhsvJe+
1qpV0k9Su24f7lD6/YMyIOZW6f74NSp5JAndVAcyfaiROAThiUn7eTLWwx+B9bfU
g/BPw1lEsI+aBOX6K2zfHT/ZhxIFktu1I8UG725yZn4B1RiPeaBJm/pbiAHbKVUS
lnkev/lURvntx1Cc0mrQXFViC0Y5OAcYwcbmvPio+/+2xrLJ40lQ3Xi4II0BSK+W
NbWz6M3e6zc7GscV9OLexGzd0iB/EvaYJS8yg+7JkNmF28Kg5DOW6VD4xrdKh4ZZ
3UYnCMrAWat/ozPhBbwR/ZvMmyamDHiFJdOHrO5ekKyeM7pDyyb9Pjf4wlWWmUrr
Zi2eS6jtswmaSywtI0ESYmtTZ1UDcefNfC6MBQhEbOwvPJBS613QMMzc5u+lJkpq
qUo0qVb6DCriA3guZlGpxnN+7gWIQDkHsaD9+w7KcJguzJQaMlOKzgkgkSqVRP+z
jeNPSLejMRK31DsU2q6j+mxAMKkL57Yshb/PNGVK3cobTOxN2iMYmqH3BuuYrxX0
F4OJ8ACjnf9CiSMpBSkY3vk4hM633qXNovjxUlUKrbJ+TpRtlBm4XNVhkOdVaq90
JO5rOgTADlYWwEQ7mGewLcJGEXl7Oe9kvnasyv1MHPyDepu5vm7bBIa5YrwoaJFd
tmu4iUjp6KA2jm5cFOQtnw8IFzz25Pbd8Kx7cDMEb4zuluYEKcxu2o9i8ZOmvxyL
r1TwVwpxYhfx5zI1zkUkyrntkKGZjah0LkceEMsEEz/cpTpGQbQQBJR2HI/u2v1N
yCC6rXi7/MtSqKeij7/JmNu6eg6+NaG78i/TxiKqi1G86KWn1fOexAjNBp8E6e+c
WG1aAOrlXTSXkm2J7ICK0IHzfkiaQCiFuAGbiK4UnSFr4sN4r4RU3zFoSTHz3w8F
thtv9cXRNKUN7fGx7ie2CxKUYoCR0TQVG0TJKbGThuxStpejrRgJN8kyColFkW7f
Nc1v5gxj5AZMzDRpnwkGFQMaTCB/qSyDOpzUoT2hc8PRZ6nsY5WyI4YIu3o55U38
RWIcgjTmsaclWXzY0OTaJ5QBMvqqgWWybd4FAJlEXjM++KI09tIoE7irvWIEvoTS
DANa0awblbZHwyzvKZJ0xpYmUuRsQvEsWR7VUUKRiXn1kUgHEvVKfscm6vnsJmWg
5uT1F10gr8sRPzodN061bowkgWGEFk+ttJJ8JN0woHYFvOp/ZnHoZfmb7+mFbsBG
QtXlRPxFbXYQPSzECN4sZgVSVNuwzBQOd7zR1ZhNIBwudcXrR+fNpab+Kw9AoCAF
AjbaAVX+JNQXp7D0ouvqlDI+z7d8OLu2UxejGCHcyjkIkw0NKdyjttbatBQK2GwZ
s2xi/fvAqCG6Oisszim/ZU2rtUHsIZg6fggrBkqkZ/isB5kpDTP4sgDGjh/75DGj
EwGl+VfKBzVnyPortXXHk+OAmuN0LX+GOCTEEOVSi1DMhmnqxxY6xg8JaQUUo1HV
81hjpmYngdsBXmA1p5FfiTce3UTMaj1cX74fpwjt8+S4MxuKAXSuM+MGanHFb6Xl
uLM9gz0lG+n1ecHW9phitnZr/DT+r0oJNXc+tHagEyXFJhmiiP/CY+8nm3kWgBn3
iNTkn+bIIEp/dV3V2oB2sJ0GRj2A6eIzCicB8o9m8/ohNUqD0fwVZDkgDCLGTQcN
JXqwSaBQdocCzHfcbfDINFT/w1I3ezNKnbPmsxUrb/Qq97f1eoNI8HG8HYw+I29r
k4n6qJWxNVzZItU5fA0n+tHsC9Pr18vu5RE6a57hLkqjB65Ik4YztqpcmNKRSdnz
iMxNEHXMVjHXfFYAehfVWjsQR4MYvO7if4Go717Z0JqWM2wSzqQiJShUaibrshv4
JSv+FITCiBjIPLL06Lw08zdadH5UzARNfeXWjPvhHRve5waQkt37lYKKgZedew3V
wvw94YhRh491fdSMVWY8B7fpVLrCsbJIsBgQRdNDN3t6hKTQoQiu+Nb/tE3HyOYC
hPulTdHa6Pq2zlD2lnZYgaSbBIWJ2LZL9fIpdafHpAoCP53lcMmbK4eCs+uSl7Ft
KmOAp0AaeJBPX0tMY8voPbTo8AlBliV2m5Bsrd7uyU3l6Bqmpi/+V4ZrmjvcN0Go
CLB49X5mJAzlY24Q2N9kp0u3DJ2sthODeogXetA1FYxjFozO11sEC69y11ePJPy2
5XuWPv0lHsocNwsw8+QdJ17yWurMgGZRXVhXxgpQMf/0k6OSFytmFLJK6NJQf1z9
dgcR9NZ+r2Y38kUQQmHidnJVIqqDJO2IJKyQpnamxVn1OEHMo4714I3Y42tV4KZC
QYqnbgwzxiNN1EDN4E9eZO0t9HqGcJrc/q0s1eprOBDf0+69JYpHn5kaa7EmaG2C
MSkq/lJi68annvoTbSP+0kM7+MnPHSiV0q9WL7JxpOVO/s4dmZasRxViCnqhAock
nqpFpzpaoYhpo1qFYTxDnmA/3vLYQVuZjgREoyCNE5Q3Iyd4yhEryPhQZx1oWNw4
Cm3nYs/yaUMcyTiBDe9tSII32G+hHSxHOqCu4LI+1GftOi/einqJhDx6Agtxq1iw
ZZph5Y4fm/+zMqQpsFcI+t7SJslCBc9nC0iwPP0hw6h/kuQ7cO4OlqMm9AffTLzT
+Ic9ku2k46QkUbWQKcURb/oNGt3n0H1BQJ/KwcXUSxpZG5eeIvBgFUadznMbJ/UF
Fdcg4ImnwhbNyhDf5hR3VMZ0AI/9kXrYjOG2Z5jltHaeS5LgFJFjjuM9cZZM5oHp
eCEtWC9RHUihK5+2BxZa7FEvAAiYW8r567soWzmKx+zcYB3LnAl33+kNBihPIkP+
MoJ6os81IxqnIrBfhtUb63BNchUlLfzOF5UN1Te4KJxsfy37LNfDQm7+NaYDHVUG
/v5Cy4Me6aFovDuavQp+hdz1eiyTFCaAZVI5fu4sXI92T3KqwxvtzoYoZ/qLOZom
pi4+Xlv9gPAa3beP4pAJr6gL/BJx7VQKFU2wJb/ApbQKrTb06mlKoZwH3PGNYCW2
0ek/32Bnkg5Z+NBMCyyus54wStu+l3JpmVrs/cGuj1HaPvn88tyfU+I/0kESEYXT
OQXj3cFzXgY3eaF8RtPDhuvO9QQjay1WutvjgMWIQc3DB1h7eFJKpVkgUWE9dEOA
td18YDOJCMgeWTGuIMaRpEa6d5UtFtDP+V4EsOaOA8p8fDTzhtkdmKzNzBD0Vd09
mZVxwjuoZ5n1Qbq8IJLMGvJrnMIJnUqFGOX5mwb+SzmJO9KWvcIkClmWx5+1DlPu
X8/UugOvMityQFB+vI2ASvV4WHmU3c6UjrN/qg9YRfGuCjsn4yuwKCe+ivYfd6Pz
SyFuImByvOc2BULKgGXcxbk079jEAp/za+IiXfMPQ7oPSNgfnjuVuecWHFm3zMnu
qxrHNOVccx+/sQudV+Y8nsBxx7mBu6A1mljxJ/B2ueKGJD0N2i01jWoZKgElaLIt
LiGSZJvhAmvgU5iWCZ5v0G0RuyduDaI4DeT333c+rgFabM+J0zMw7yhlpkl7IBmC
azeTiu9GWyuWifLY5MCHHFvm3BcXn0bb4QLfhX5NIS7kZeWNbmWJhJ9iHLRZ1TNo
K6IsP0DCcpCRIYGLwkscLUraST0aFyVVWkmquQz4BAXg9I+1vY2OuNJ+TlH4QRk8
s+n+NL8MLG1iU5wu3xLjnVrxRqnJoMeWaBFEzfz4Kq6yhuLyHVMMcnLbTmYJhAZT
AScpl67r0IKmcMtA0nNVDPVgvtDRnklao+Z+mxTx+S9ZXk0VrM+FeBtCEFVAGILO
uJq/u6qkyaqWkxCrD+ercCSWEeyNjKz/hWkKJBp0rj2dEVMjU75PFHdbwbyVMiHN
9UYUe1jH9fz9cgKeDeaO18Xxv4C/pVA9NmFKpyvISHXIiDEPqCUYqNaV3VW6sEEZ
bpx0KwdVJWscODG/RPAWShBgVH8WvMNdks/bzM6rfWvbOJ99bQt9YkeOYDifYjSL
d9XtF2vyLha4Dr1jFDZNU172SoMg8ZiuDLJYC54IN4fX58EzO0ZzH8F5DTMwuZCG
qWmqaxMgrF4aw3W42oVjxmWQha+JuzM3M3LTv7Ck1Ykaz6ChIpZaFnO6TA4FAoPE
OGcAujKQPPiZtdYvH1SqAWhscMk0SUOga4fFv4taEymSdujltlNe2i8lPvu/Y04o
Dmb9s+ui87EHxwqDZjlxjmStiCQNKcY5IpDnE5xjQCEQTAz9Q+qOYIy9S3zu8wnI
YqSwohPg7bkSKITXHayiarobStpo+nFBTjbQGhL2FE4y91kgVcWJ7MJygYnumsyP
egGO8WPKQsCF0MuXkXNrJtvDUzQTDVNiy6XEGZhdKSLMJZaPE/yUwTshHyzIdiFs
3hDVq/TbBx8axD3Nv2PDG2UIxyHy679hnTNkoWpemBqalidO/RcmRU4ImAtGZ17f
ACnsCCEVlZwueJ2OOTT3soGkFRYvRTchW+2S3XmwtttU3dPUAAVzdBkTrsnaARmO
txl16iIvfnrM27xO/NfNMAfBqASyBJjJ1LxZVWNrxZZeJK/7hLjTh92KU2Ro/ill
TuXFJR0aenqM74y4Hp61NzJP+2yoywPkwgWpCbvVCxyWM+CsD+N2aO9uhD/OGmk/
HalHtN8Gg6/qgoxeIgzlPDinetyRWfacDfvNFD2/WsqoWmOAGrxeevr88zHHusQC
4klLNn1z2dv0MNGPF2Ig6PWpMlltH/CVgzopCUPS9sIuAUHrZivscctPliVm5jS+
+1OH4pRen+VesOQzcEQRmuPPDXqgQ0Cl33JvZ8BfV1urMlCK0GwBGgSrAW/9H5tL
BbRENyoz/G+qpdOhuzcQ3Mhuk0hjAZxZTfEUrV+RbXdOSYx6EhD+lXY7Y43SQmPG
wCwnQfV6K1DIeL2swyKUwHrWmGyl/yvHqgD3CJqC2+s2sSQHwQkkhFooyBgt34LN
l+jBBuZ0g/wv/+cCb+fO+JuxqsMWPCk2vog9fnG+w21gygfexpNBCoNz0vVCz8Vb
V8G69W1WakC1YhhO51TLusd3e818F7rWeUyyAOu/nj+ZN7qtQUNVCtBAdVBefSPS
MlUkMMyFgBgSbs8dvmvvHgqQMl/vsG6OlvwAyPUQacGO/iQBKlGv3Rqxpa1erUcv
p4qIEMidgeVJhlkgrpptSFG0tTgEIa5qIHZZc/uJvd9jJNzG3EUxWSksQpoEVnfH
6oJz2EZkYkbFqu0Zb2grbim+/hps3GiPOMje3KvI7vwkuDaHz9lMjM/u8aKXZDMG
Wlku55DXcu5Z0oF1+11UfZ/mnwZ8zv2mYy7OwUNV5oal2pyPAmGay3s20yOZrTMu
W6yXyjOTSE6JIzwxjs7BU9gJRW4Mhduy7bsaPVCCSHfSSxtdhogR6BuGhSWTsIcp
pK1zlhZJ/UZbNqOeNyvdvUgpEyCWnFed3WaFOJnhDT6UgzdoWXCz7A/hggYptVhF
1gRabHDIiY9I/gSDsh9m05c7UHk49HQthK6cFWgwAD8YEoj0z5B4l6IHCcGa1dr2
vB1S5YTx280S1Fd/p8nCXYCIjvooGz1b6gRNRsbX+oeaINXadRnQZvBSR8sEEBpV
sHzNMrgv1p5S5SzdrhnGshjUsSXD6nF1oZtScoE2HhF3FXyqD5d0mRgCySjdKR3I
gR53fASLKJQEdNDpEAkaGeohMUeEjrTRsIkcpv8lN6ONLwem7BGYyT7+kMx14vjT
c1JBpnT4q5AaaavURnZO9Kr0S7n3B51hzBVaY8dc8s5i2j23TUBCzlKckRr+kS6j
0FuWLyQPK+ef2eZDPiEdR+DJHCJw6UhEo/vQtFDqJSL5nYGfSG0oJLBhptdfqXGz
SzcTECCful9+57MYMZbRHejd+B1Y+lahAB5GfnNAMc8GBQ5tzZmDMuG6Qv76eIds
tn+6vrT0nj1Rwk3OFT8oZAtNvvObPmlIG9O6APWLGhAnqtX/dDS5SS7Zz1AEaMJj
m0ubyzBxcD+hTWf7mPToys2dB4J/ltd36d3IWQtx4MbCmreXIgbWA5+M/10ZEJXt
A9Bjh04WyjEDOz2n4NatHkz6AikuAoV9lhHln2at86thn8KeLFbPVaN3smgqFDq/
I/Lb6Qcp3k/9AXP51qOA5o7rhmcluVMu4PtrP3co0L6ifQwRatCPYRdVTCb8tI/S
NcTTRxe28jirNeppgWT15cWpauuy5SDJ9OAwg4F7L8o7RPhdL2UA4u6nWo2sij0W
246srD0HHm2v03IyuZkwtPvcSbjR1lN2KkPU8S2EzswBlD1WI76R/BUl0WbpCYTy
9fPjFTd1Ah/jwKEMptDkB32PBMlIB+FagIJ1r2Tc9p9F3OxqJP1fcYw4bU+kfk3u
lcc4+akho3dMYTtbmDbK+BvlvQZr3ypIVhD7WUJzT/iwxHgEwmbsBobw+b+2NwQO
YXLKJZAmkIIRxzKQpa+2haftyqU78jSKfOXPGbgD0I3xdg4wpbakMPQXe1nK80pm
arOHfQqN5WLb2j/t+GQ3922rsXWRIqJmGcibNwS00pdMbU3+r2yyXgy47FprxQqR
Qnj2u/hOvU8dniOqre4tjPQSZtZ4GEpQvjupztTlBAQsdEt+/X1NDXfZd1bdYAzX
nBu9e1lOsXGykOjmSj2Bw5qaxl2pCrjskmWnk0krxqz7IV1xTxKHiLOnVpcYGOEu
Zm3f3hpmRdTIHgolBg2kxa5nBcRj5t1DSi8o2ZVWT5ga8RtvKj0qNWg7Yn8entMt
yCS6c87gUrspMjPW3KJ6nwqPnzj/XAT+/bpEdK5AHJR6+1xJ8ZdRQNf4H7Cv0UqR
hgfUGEvCrpckhlpk1FOkCXN3gYb7wxSzkRM0tfALhzafieItRd+6hsrG1eOmY5J6
kmsg6/Y8rv4JbTsvytsWGsYWeFU8FTRjb0swJyJKdgmur6H1r/tXcxpAWVB7G8ap
NI/5lGOOr2YtrVE1XE9ivq6L4HjehW8/bqa2gF+HxVRByHgRO0fEksmAP/nsswpB
er5LiL0mg1M9m2uRCXyyxKGsmgyB/h8y6yU70e+jBMSeBJ/z5yUdOa9C09KYsuBY
hr3btLb2OOZdpBucWvXzeXsZ4wDEEbw1uaidpLTeHrGQEQkFdm537okUbNjy3N2w
7X5cOJuXEojTAmtUGkWl/pxZn+y6o8BJzeHBfeO5LDdiiGdZ7vTVq6uJbKXzNja1
oo9+llRhOHVgsWxeO2KZfhi1H541aBdqFrmgsdc5x4IWAgzyLK1D6wtLl0uAt796
gQY2PQBqxXHQjZaOTAzalS/W0/ypOUos3s3j2zj6GHLuX/kssrXhr1766uO3zBWZ
udwwkBpbSPw+rWyCtcKKrl8ywNpCapD7lj5RjCoj+CgfFwRJIzgfWHMLUSAynlTJ
ycu4HXjNhRiVRWWuU5rpsmwbXkyGrzLaDg5FxqOJfgCjN11C2PexT9QTZcyT83oO
TJC/Z33FM+YYlbihA299WWeQH0siEX2fSVvzS4HIsnZabof/dfOh+HYbnBp6mJDa
HmLN2XxcxLPwG1vIEna93Z2BvcxZyfKESaXEt5Z32ByxB8SUG3U3dBXPUiFbYyMW
OVKg4H1pwJE119Eysk+u4oY3LGR499fs+kSeOIyqsry+/WFIQ0GC/kawN/mQy9We
qwnfy6oJrDkJkCADLfuqrJsUAxAZF1BqnSDe7/MVLs0t7slULZkYO81Q9xmQj+oV
CcNRJw5waXjusKCn1ScHamnlD+CqXwQO87GG9aKT5NJPCsoJi2E4MjUjlTfOFVwc
BsPAgroJO/wVeEfdSuR6WcAObxWynp//8l4SMN+55Fdf7eZ5f4eAngxLNgjmISv6
vClyogyXphCIYixatp64jGnZtbIPQsDhSOi/UUO7bGL6tPCuvBM1Q8blLkoSmegY
32OJDKhXM5Fg+j4ps9rZ002ufrQDnJI3NCr0xxJoBcK2thpNMtjRtSG+jOjftvQY
P01O49LgNqlSbGbh3rwiEEVxqZINx133V9K9EGhwVm7mQZWFIw7DGJDUODX0KSwM
TsSXsNsZqcWUfhOwlT22XnBJalur7sJq/l1K9/w//i7b6t8XRkNHEavTBE45Hm0X
pKn6b1N7egO47oDT4SoH7vsrd7ze5G3Aerh0OJQFeSaiDb90XHDNnn078XdD07xf
ltEKjJcWACw6sq2Iig2ppXSa2/u8V8b+2fnVJx5YugfuX5N4IsCI94hiEEaVjnKG
NR2RRHITkPeqNNl5HqiohCfugSZsyB6Y6bpYJCXaaEa9fHQIDKT6Z0n6eTkh2ppc
ebxneE6PcB8dI3NGcYD86W8/+9PSfrpgqHbRlsgHJ2+lEEflsEZc/h7iTQK3Bymy
wI1LamXWbnhqTyOxLrk/9Cp/7eB8O//Y1XdgszvE5JQPAoB+zaOljCCjWzzPbQ16
23oLnIJVIvkr2isQAQt2qSEQ7TVPUS4oVTIrPCFm5qZxKfgU1Qxko583v1xShQYs
TZuPhqTmY0ckGpFSEjxPSO/Wo5wFbDzNJv/3AmN/sXSktL3q35s3ITccFIUKW6MW
Re67RN9uCerGSzsHilgyI5z84zdwKXE6N5Y7z9HHhGtF8eWRBOBSTGrnVaSWlPPP
Bob0Zju00vonrqYQjSIqgvfTPP4L5BMJvJKklZxLPQeVgvSIXFVGGsERx4IoJdo5
Z513YzAZtHCi0jA9T5ZaiDNHTmPgda0G/wVc7cG0NiKPdwbHoDCAClXyXC6M1j19
zWbotoYilbYKhKDNKITVHNMUufSY1jbvOe2UEUbKybLWdoAI1dDpbf49nMLcv6Ha
X7/FLBGc+XcX863qA7l6aayuFtExpxwpO2dl7GDnKFJTaB+GMuLMwaomgVbCqbjM
XyVcaPWfrtWNoOqvs+zZDPhZY/bFUE4DlfK2FKcivzFW9KJJvK3kXMYt/DmCRcMs
7l4XtjiwfwS++2ZHGLpflsGmiVU4Ji8UYVmtiBU3aQXAL/R4zrn72WF1hWPwa2yv
loXakiDFe0T/FR+Ysgv/ib5399ScNEFrHdhq6frgKRUVsZ2PMnbLHu+oSsXaJFFz
TUOt61AizX1zo02zWoxGGzrR5+afzYrX1Jela18AkE2bb3U5aULDhtXaBvZgh+LV
68ktpPwh+zPXL57jopbj/Qgql88YWjCF4eOsavqQlqai8BI8G0rZrP9IBGgvdYxm
niQnSWO+ZkxDuHVcUCjp3NME8IaqRxYpK15dG9Hn9lYgTMmb8ijoAFu9/2vbjLD5
RYIOIQrTKDJGRhqm3pfv6xoc5SP9rh6h+EJWZVgKnr+M0NhjkfY5NgrFV4mkAvyO
rM3QBrr/Jc0GtStImD9FDA7VA7pvZIxr5cxTx8DUTjhwaq74v4cYwL4xwHdepPXz
QqX/9xsmfgM3E4xHmxltrEEdIDbBnaNWD/C+uQqnXvBjs3VDHnC3xLvHex9o3RTn
HO/5SrOJFNMIBt93dq4GmWXS+8vED0QnzwjmW0MQ/eFXtrtKCVflhqFWKvR1zvAi
yjDfht7DVGAX89/THMj+rz/pl10J1VV6QgsHFmAxf4xmVkgRnipUGdr6o6U7JmMf
C3kJn6fiPVpnbIB3eA0Fd1/MBqCishxr6jPPLGZl73SJZZXd+aHPDtiexX62djMH
+Ped80gU5ZjrtY+JGizZ4isffnDGRiOorvcsryItvpKqK10/IBQEg7O3CEDeOLzL
yed6C6Pzz/SfbvdArZu7RLLHKFsIl+ptWCdQ1O3lZNQ3HLUvjwZoYd7bVPYu3nD7
jCXRbqlhuxmXpD8VEyi5DS5pToFNCTS0cNh2oHbDSBR4pSk5ErrxAt0bmVFKmpTu
VK0bchrZD5CHbIYBRIbVb23OjVDq5P3VvUyWJSn307ztvQ3slXF7Fbe34gqXiZ8O
Iei2bu7w556L/ceBQuOonhPrP5TjJnfug9G17oKVIfJj0QZRKyX+97bpUrg/b8Sp
X00rwT+htpADSJDICjizpxASweq8qSSfiyYJR6b5PR2dd+S1hCHih1i8Bt7AA432
hdK0wJGZyAMgiIUln8LC2HVsLKCDK1hHPoZ99b+GhmH+oB9Bt1Y8OeGpEex3G36R
mXJklkkXMxiuuVb7c79VYEM6QoS2G7vq0ecDtn4QY9S7vLDnB02yHkNAaZaMdA1G
bQBS6W4vfTZyGvuif1t0H+1YDDeYn7NsUmBYTG5Nr4UnJJxFV+LgYeBrjrLSl9ea
m6yCYUc4gZoTxaUdHke4y61n6X8upBGQqFbCwNjI4i37fyo81CYh9IHvsz6ZgDl8
MmNbLCV6Km5DGJ8Y55j27QZclLMYG+SLLnaJ+z4YfT4wTsjtflNy+g0MJRgT9JDK
lECVan+WvzFQKQART7dLtCO6tQTeljXzCjCQQlDvzuRzaITXaVEs14rV3bSR0Yt6
NEhvJjAfkxhqAnS3kiuBD2CIYHWiUwpF/HD1Y5NRZej1BWhHI3/EXEkRxO1GawyR
f6tec0RzIDZhYuQKAsgD2JQdoZpgHaY492Qx7UdeLHey7S0B+uyPpML+x6f/FyHN
TjbFlD2RU0or0U2A2gIosPk4/nebC9boXtlD067Scy7EMo09Rcf5WvUw+iD54G4t
RgElmGomUA5KFwGwTxzBIRnhrPUF2bZKjXI853CtT8nSRmiWGG62yw4AhnvWII38
bzWy/WTTJ07r+QvshhZ5HqE8mlKd9ik2bcRf6ErtSiCYefX0VphupKsDEqTbePT1
Q9QwlvbM8dPB9VTzi+lX3IrFlUNEaqD6OJ7NtrHKViqg2M6QdxM55HwXCia1BMdh
vz7OExxH7En2+uaEhhhGyw==
`pragma protect end_protected
