// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hrs+OSiQbCvbG5rqjcyz2iUHzBq8zoZpGLL9gIAsItxLgNUXS8wzDCjSFwshK9fv
WOjxIRtc1FgRRIcX96CPSiaclN5AxJIhaQUKicdhvDV+dQgpdSzXxebtXXlnGCC6
NuiJaIvyEjhJrQ+aRCb9gMM1T2gFE+QjChpsVxpHoHU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8272)
oBqObacan35k1xWelxkR83+25WKeK27L1bk8IVjh7Qxvc9agNunsAavLV201MSHC
l4fTTr/ITdB15poQsRPVd7W55U5dnFZ4jTsr4KILY6vorHn/nh+qrbFq3KypBaS7
XjRqcx+mXLaC5jfGFZ3cdF3BhFkgNEQd30HdbF4nOHQpb5luKZcuwko+ppDBuxLY
KPpGnHCabRCZWQopqVnWxg78tvRRc2sCRzrj41qFmTgqNY40W9kDuVSRz4mrfIm7
VIln9xR5JWA+HkCgFfi04Odey613NSx1L3cLfZ7zM568TzOFVs+PdDe1eUboUgl+
XyAhCNzFBCmSuRdd6AQBcfNhsqTJOfl+lhr5XHgpIohKTFYSVdR4mYjb0KCH2n9x
0ffqts84uIfcmBsUofxOf6imjwcM1wQwri+4m4tS0oUNMWyo1wqbbXAlcRe6ukEy
cs3Ei6p4niCIJ7HxEe1fM3DXNFtvVbMK261qrMkdLbYwQxuDYqJOvUWnpAzS5ygo
uJNfrnIGlPFRTmpZMLj1gHpj+I+sYp729Ewi7JhMvg5B9jFQilnU9Q1z3c9npNO5
Zi4AAtkohanftfJ034OKWEhTv/8SRA2bMReVWOtLjI1gTtYVXZxfp11yVQG0Yu9j
9jwTCzGZ0ulSLa9RoD0guAqp/Ou1jOhfP9ng13DP8TznwEZ6bo3Xd69svZYFF5Tz
FVF4VWHUgKmK7iXRYo6TZbApScUX3NMDbgAaK2cxPCvVh8nVlaFiIotK4BdqV4OA
DVgTBJ2F/nUORYowU7zfpY5h2uCUQSEfXP8Lq5ZiEzqYktZ9nVXL97bogQyYYvm/
8QTQ41x3xTEFQPPJR5S/VSzpsxbF4BPrgzgovz+2kU6TlLmNhcV1GYNUmJFTMnQQ
Zm7ngqI830T3WO7v3R0S6kS9eyDV9PKoPMXekDHuCMYgUGuXXyi0ji/FSxnSZncd
1/b82IZwDEipz3Ga8adYsbZU+XtXN/Zm+SEBpH3xjs6r6+zQkIoJTtaVmqAfQ1Yd
2JFwLduSotLsyWLrgVqBaStKCn/o9aZ7/Gn6zKKuBzgjtLGtCa3wsDee9z3min3F
mgrB6UAoyqqXy3ydTTtgX5wzrt73SdYIrHWmX2pEQgyiIR+iAZc2o5fT/HHhVwQ3
PdqA3UpjzMkRHWjydMXB7jpWH5a/el55fNrXHa7uWG0crURlYDyOPAyzhALPZLAC
kC/o+DPeuRPepeZrS72Sdpi5LZvJ4y01jv1n5eoQ4XFvFbFnPo80/N06SA8a1q/p
S9yr2GNDiMOeNtiHOffbEZgFXQLYzg4C6+GJoNg2raqyFqYia8DI0++h1sh/H0XJ
dASw0KQmP66aHUTdoldwhK24q/+vwJY27M3jDyXih2TjNEyOu9eJcbI+9f6HH3Sr
ZJQGK8oEh8+nFPpyBBHL+v97Srm2hv9ci9gecPwNmE7Gds4/aP6ggWKP+ps+tt7O
hrFfacH7aA1GEShqoaITjqu3v96zN4xr9cxvSgSS5Pja5+zUHKFZJzwkAmU5vwhq
5cMzF++jm8m9b0Iax+iNn4UKL9Ex9OH3/3ba2WkXCd37VWrVPF7NYyJs0dnoCVN8
JhV9VTqi4Hb2Mdn1JbxkSMF6skwnHxuHkEKoIrV/8cWzHwu0VFhupnjIDUtoAB/U
aXPaY/M+Yygp19qZXT/Pf8rjON08sWiHCzgxfEQTIJKCmgomKk9JiH7Ti1PKU2Yd
lCM0ueS7W4atZ5miU46/uXAL23N/DwRaEg5H3cw7U0blBeKVYqyA349zrrLP666g
R3up2K/YSqu0zJJbHwJJbL789bzCRPD7yu/nOYJp68sXB4uYn+AQ5fiQaK/CLK+C
IjWYg8dFL3mI39iQ/CV/1ASTLCpebRpfi/ljFbgTmbQ8EaGylbNJGMgMd7p12z3T
+cOgvVlor1f2/T1aK03drgjTjju2/HBAwQ1FD//LhZg88kv28D+NqAoMFMlBes2G
9cfcSX7LsIQyX3Xvl8TW61SdO1SKHlZOVdxChIteXA9M9oJEtyaj9nnOYjIedAWq
EDYJWxob9jKfngOuJXAz6K84iL7XJNpGOl6bKp+wRNoplY/Ec5r6eGtGpWLB7O/8
9R8B2C+64f3drlWv7+xMM1td+0o8icP5BPy88rbzPyyrwRtwQtaguQ8CYGfG5H1/
VcxoLT/Ts+1zIzaqbogC8A/HWoDkHZH7UIrLGRLgrzvuor5vFUww8+b6S0Y8L+Ln
5/UBonkOtjypjzemGeZ4ulmx4tQCQ/oqNjO3xAcvUAno38bMUBzqLmM+U3p6KA2Q
oYcMJhxTSP4Zm7u7mnEZwrpHSwdbnup7jAAHeIA0U54Z7lGdDPCAhV3lgrIccIZ7
gebdkqjoovcHEAR3gfUqjy1H+QeBjBerdVvsJWiRnFOvdA+4tksV81Rwu1C56/RW
xDD5vvuWWBIYCaQbXv9LFk6enI46cowWF1eovD6mC0+eUa5FkSjWIwxsTs1TtNIp
6Ci73ew3+OYtWYX5EQw4n46oE3AOiZTrBhTsWlx5VXgnn8/gG5crfAj4S08AwQaC
yTkU/p2Wl45sgCSLeK8RmhFU2JSiStSE7YmQdzJQYsIsagwL2AzarMLyufiV3TSQ
NH6lkPaJbxa02fPt1YbFxiyb25PFtQmNvkxoNQR+vTa81Fq0oA6g+pHIGR97tRZM
82G1DscrYZuXX8PdAq0ierJxCvWdnd5LDk7qd9aJV8Lg+VBaXblJSVsTqGkt4UCf
2P7czBs/IYzTgI9uiMfMCwjoaQWZ2MPFGphTHAYH1mmYO7gc9aerdGCRtNfK+GHo
MxaEbdHG/4fVh9dclFm7JK6bmExhZ+Obej3cboszKJGyMcYPNjVUgBkNs/nTvK1Y
HbBZw7a07T4TPFcST7dRqq3MuG1YqxdS6arl0rX8xOnCxAdbhweKFDmpMlY3OWae
Bza/zqbcYPoBC3nVwBWrm7TARTX028QjgSaGFYLLRtDqmxIUZz+tny2hq4sQyVzZ
bdTPrY8qNUxch49oUXcaabR6PSo9HKJ1y/KvPe0eJGCrjRcgtOWCw3F3+7VgnCs9
1dXx+TrF73hR8q30a4iumAuEsg1//EeJqBpMtj89VE+c62wwv3JwBwyvrRZVBz24
GNM7l9QJkUUUtIcQK5M3OY8c3qxYw/f7vwejBEN/pGo59qjU1/ko+2+NdYiKMALo
JCuwdO6t8MCBHohOK140G45Bzr/s1j1smMsB9PBd/4kAI5SIbc42pryI8c+Tqyqq
UVi7j/cyzd8DR7xz9xk9zG9cNOCl+1iIIB76HNGNbWxNwjRw5cbatADNBNz08pOu
zDa39DEfYuaziZl3h5r9ny7w18llO67gJAATtnsRqFLtv2L8qyRqSwfFiL7ASylJ
Ifo5fn4K4wfs/9J+JUuUOTGi8RtPijeY+YdfgOG5UuWOXnaQBIUNV2ef2iRrf8zx
q9ZXDp03TWVy7rJWAMJBD64izt1W5cehiSBKnKdOXKZL9H34Qw0zkT11T4QbeQ4o
/1+m9sMoqMvKua7zz211xDv8fFW5SgVT81s9Qqea9EPaC2+w4yQvdrN3FAkC93hJ
yw5dvgXbmd27nO5l9c2BnWnkYVu5W5AmkiLuj1YFYymRqnMSCSKZxTsYhUwaBaHt
5Efn5RXrqrEgCJ4Q9IPxks0KsxdNin7Da7megdtPSqZw/6fL+jn7p+wFeSr77gDy
Z9+/DgjoVr5pMF/caC9HN6mGfh/A8CpC+EFTxw/2zHLo+/ZX+6K+TZO06MZfUUPm
u4rHSlStU9qOjxCrid/Bxo7nT8VpFOHOBmcTPMsfL/BBOb1EeFA/GmG5UPHGGJH8
Y2bdysH8/1d7+uP/+Qm8v8G9ktCUSQuHoyw+My1ACHbzBh5PiTWWo1SEZlpLq1Xu
S+GuIGqSfF0WVKTn0w6s3/yxrPqpcfHyPLs0PMJNANjCGIpPzZMLYSlWykpJyu5d
h/C76Dr83FxybcFx0Tvrs4B/ZSQX2HEiLvuMpX7+a7nO/RSa3bYWFqSGztEvO+2i
7dqHg1QZy/GpPJ87LayOm50ASlPP1ct2AgbFN6JZGZINfmtUzJ6zW41mx2ti9TVX
xB4GywzejHTRiR5HtaHSbCD0H48J4oBAIS2hS14AHffCVQxxsh1Ll8J6BNg6oGDB
mmSOJLZJanQ4OiBENMQo/AHbbJEKuMW0RFKumTYMLIghaw09IVH7dnFaUu6VP5bY
+kR3BCM5ncFHKsplGQD4hnimjU1FkfxJHPtujiwvq3J5a9YzHyt6EDdhMd8pRCDa
eBZ2JWsbiABlun2f1k9K90TEV0MSECSeqFHkcNylnJ/UGtmuSZ/07T+74Fq1GICS
bZUCu0j7Ibbj7cGLMmuzgUMTRvaoKXre35v8nTHx9s5M0yYAJxdcGPm9EFuQiCqP
uqBcQPJ3o+y+C5OXRTy6BBAZHU9YBDuxtKNGmtjP4xq8yDH6whD7o7b9SIbjTJKZ
4fnpBow7YONr9lAVr+ttCP7p7BD/O4k4ajRJ7Ah9YVNbqnPuFeJ1bNuIzoJMzh1e
Nhu0hNMC3+CxcSiaWR+4wn3qIhZbUZpAiP5/jOVnHwuVfIfdRaflcrQLHWcm4BNE
ZKrKkGk/VmfQ83bOuUIAV5B+UnSyhJmokVvvis8pJor8QBh91lTrhDVGC98VxzAv
i+gzLiEGyNXS7k0obvOFSPCf1TCmI5NxqsCkMC6tDccBePRF+SbOFFa5xSodpuuO
l31/RyojBbmBix4UlFxGnhW9Fcv/MnBWmtj63L2tpLQbltGHfmpXqZko5IAZKszs
B7oE61C6Q+UWk+mEQNX2acgUROA9gYizjJi+YiY/NnG3KF0tTlg/q07v0ZQqglfK
yt6iEdoYVZv35Ubku82TuM4GXPbUGOMeOMFi34yRP4O2Y34WHxHGISxNHmVPYhWB
vojUdfcxXsKqDF+0kGxErEyL+aiSQLKDEZjiY182VioG0Ly45I3ElV/3mZ5G7ExU
G4WDSzNc8tG7GFb3+xCuphj4HDQwqbsqRzGHghe1+6cJM5aIPhQc08U0mAA0tAE1
6TDufMre72ayOUZzuULVRZ2HX9Jc42ZxZOlpRu6C1iSZXJWzL+d/MHciuLHw4TI8
ZTCB7VtXaidZabNy5ThuhsrOkA3mAr6ANUaPSOXEDHv3zkVXTbAHUiDG/KKTB6vE
/FfgHrfBQgg9on380l17Nkh11Zs9bUuSW6SgRdyH4nNyqmFzi23K/QrMUU7+IqG4
y5qI6lajOdb/6CGp1Ia82zDX+aKxBmaka7qho9GT16xkUoNWeGgMpcW7Vhsr2pOD
jofgm4VagR1p1axctqtP6rZGkZZsjSO+hulLyDSLDsH9e83UZe/U1jW2O26UpSuZ
oewb4DoH+kYK8oxOO3xagSDugLSY8zQP4XtBGWPxDgNLJC1SypqJotSDgPHVwpST
o1HMG3s6NKWbFOlBdaw6ds29kupaWbN5s7DKJO5DEGkJSRBy02BO2L9j10qTfsOo
jV5ePvum8M8t+pPaf8N33eoRjAJ2n9lqnft8ek8/8ejBYSyroCUjLU+U+Hhn3rY0
zf2Ij+UtJNCjT8pPy/I+iGo2+h8uiD448Afo6l5VzlTuuc3b9/cRI+M2CMl2/kpz
9WHMS4FiRB7OjeecibCU9ET0vh59/0H1T6oC41bbMDTpfVgSO1bgPtCWKD78fySb
G/hDwIGbiynsc5LIv5w66jd4Sd+yeJ79gwbV8IOpzq3S921T/2xyH9a1TN+UutPu
AFxYYyRNJ8qVsnXUB0PqEz3yuztalNXSqCiwxJEC5vK8oU5+l55a/GS2oan2eLk4
3cRM5MDgQwXj4qDnqEfOWbm7PhYRi4bW2y0UxVg1FUeJXTK9/OgSGfAhB+fy2rRT
hu0vV/ScDq5mXshVukoifAmgI7qwj/kSo+JrG8oiyTXDFMIH3/pIfDAJd+nneLE1
gZjK3tZU1Ub/AjdZGaGdjdZcqkQeyg8VDszleM3BCaYfTwW93Yazf/G5lclYO718
j+4u5EBOvQvvTuNIKG9BRWk5n1dgMMU14iy+HuUeZkDS42PpIUPRoR5QiIA7Q1co
VfKro7s+MzO15pRf93EYn4R3gQaBwQWfdCgNmYxZVurVG4nbB3FqQoCaNjy5yesQ
5G2G6AWYIhBL3ZNzEMmrI9UdY8Nuf80PO+SSkhUjH8k49uPfrN1AjUuoDn3AFfQE
agYMXqkC0tKn2SN4fCcxYmPOeTvZR+7iz/8Uq6XTpQpSTPKU7BvXU9f0rU3DzQxQ
kDsF9/0pQyw9YURZEcs3JbpZd+d94Z2GNV+PpmnYPE42LBiOrkQoWiT9F4/ovIy5
bmrwfkqx+z+UL7glVk4OwwwcZYjFnb99gFcq+y3ezuRLXI/Yemqky5h5pd7TL7o1
K/T8/ttDKGImvfHCwX2yBEbgOOFi6/D5D1bBSJVvdK7nrDebmbqFiyAQ6x2JaDF4
rLoc5wh2H0e0wa4NzWanjGAig81Pzyw0jKqARQjW9SYzilANQ+PltryzjynVMOXv
+qVOXDnWKaNxK+1JJTwCAKDkSXx+j70RuEYmJibpXJpiTca0u6mzRleExdiNQ5us
LpiBmz7iIMrMtpPD4ey0Ofl8UzbNVZHacaWpryT7vQ+SSgk+UmSD6GYv60YNMjUW
6dF+ySW53YuCLSBzmLoEtLhH7bKTMZNGZZUsV1r5Vuam5FEErZ/X1WwaCKlz/hsI
SnS8KZWdHiXFdaNzUd2ipnSIlovXsbngV3YWKNvCjiDxkUAv3d/4qN7Z0eDcCq/U
jwDeNmrkpjjrSDaOcH1VyHD8tx9ADFiqlkyt8GzBdxqZpmyy/4ViWecq4NH3jHwB
dRUNoTwP6K++NPtdw5FQaFPaK7KAV2e3Q8koH6A9+QilWHK2FJPBT4Zlzjgp5cfC
BPHnKjGZQJhCqh9jXoR9BgetsibAlb0dA2yiMDb/kjkcGECQJ7cWwWFoQMF1ZS2N
PQyzq5d2LSS2AORNET6jE5MStgmecmzZc538O866WcXUcXHQmU20wcbFIcubbSgd
K4NqqbcIVKxkxmojuAFYR72nZJLhCPBfd6tCyISUHRxs5rVFmxF9WdsPoIOCac6Q
kg3sN5Ha1Et3pOriKgl11TFQbIXHX1MnmFXzdwiKJ2cgOcANhLKQcSJUWiP3sle6
UGMbAVREc/jaK+wyTJ87LK/YgZW2QIx3yT9juCC6w3arMSnZBKvozsiFqoTwza++
VGtwMMsrIqLz0HzIiQ49leP5UODoNqRLssL+yyvip8GghsLPl71d6tSk/mXRgVUB
46nbxPbeF3BXAyuo+vtSFHJFrbLZRElAlrBeIzQeSHZKRkskgohjRBwAziCzZvqe
LS5nG5K0arQ048shgJl0Xq2MhNnVW3IA2dsb4I5JuB8umqz1taV+IE59Ab7+Dx07
ZqTUWqVo2JSy12+zVLZh8HXhTCif4IZAvuWmEzemCNQkiKl0DHeC6pkNFWnBlNN2
XQl9JAqaabWJUq48fhw+MpxhR6ybS2KnAq6cSFZ/mcN4cFoAKRpmIqVYFvHr/vzw
L1VobqQE9VLnCE4BbL2LQHuYpTIsCsaFJKLdlM7NqwPUaFFHemKv8r0pMw7i8JK5
iEHebB7+b3GCaU1R/Afhj8peC3w6R9/qjFAFTIkJ/nIHv0G84Hk2GNyN9MQvyreW
KYt200/HyyBiEggOIYb59yybxiVEzU0Kj1J/mt1ZurE0KJcgaHXtaIrD3ImnHDtA
dU/IPVFsWmplM2ZvH1eJoq+R4YdBs8xfmKG/RwIj6GIwGWPQi3cBllkno76FMDhz
SvLcB+BSjtK/x7i+eeyqUcvO2Bg9Ho9atC19adlE/f05VMwyL20G69ZOMfMhcXH9
eUDiyUMj1o3fsM7iX2g5f5l/7k32SzF+4Iej+UVnpd27UVKdhuFgHbOfGxjlNdBV
QSBokZDLm8AF9L4ryP6C2SZtajufumHCGq64mbDxp1JqNw1fQT4NQ9ZAgleUX2Mx
QBIXi3E5KiyS4Di5BX3f58UfS5BOttKNdJOfbuBb5KFJIZQGSYWdepil1N2xaOf0
ObOI9Dc9mj+ueXQMcmVygDjZY6taYWgWHPGRjq6naEpCMYSLmUvBsNWYrD4jhCJg
4e3N02X8ldSpx+j2Mlhc3mCoQ3TDMXaVE2Ri7qr0AO9fediu68kz4NUk3bG5uNYB
B2CTJHWyBtuFysHpC6BKD1Lgyg3kf0JuWrD78oWX+bYuB5BpC1hcjmIdaNaNl0+a
pB2YeEmKkPq6cbh9AygzEfdKeHqkQi96E8Pd41FiDsAtB0dLXBkTNkBcUbjuBkSG
jesyqL9y3HaE10tP0cY6MJqA0CGSzunoIGdMivM82FH3GSDqfFODxVxvhtvJTLlm
wD5Q8c9X8yLvvDUgqsVrEOBj/F1HqjBCXF7J4d4jKpeYhorsbgzEH4uEHXFkqrj0
pV+h/yi/5YUQa0XabPJPpXhk0QvgE4D2AUET59DRgjEtxqXwIxLTNHs5ADZpJl0m
e6OoTDfVEvGsh3rk7gI3EjLFcclEwMtA/OzXvXU4B4oocIYJIQj/SquRo53tNSLx
ztVCOj1g4+bc74cNUw6xd2Y2deT0f1I+OM6MwTH0pn8tMWDSH5x/Cb6NcNSn769i
ng29Gx3o9E6x/cLn98RdVDZanY/o81Lt5b2fGZ3aoHCY2JTp8spB5BgAxgwAtaDr
R64CLaiLaW94zunXDnEnWmO7Iy9Z18PyyvAR6ZXP+gaHZtGtoCduvM5nwNwTyb7O
+eUnzYjYFPQVmokaiXw+RyZ5WtQarSIKvzxKCZ4ZuowxgUq1ZbTW3HGvuM4h6g8l
3/F0egSWZVT9wIUxOlfAndlx3dQ/3PeyOajgM3SBnQ16BvXI9eUWhxtXptzkkZmA
duFISW7D22vVD+a3SNYFWicoPmeRYbfxhCUAJPVxraDWS6oX+8y1lIeGuIKCwEeI
O4aTqM+Kq5rMzmX8FiLfYDzIj4XWoKYnfwUEajv45R8iSym5JsJLcMZzFMUO+dRI
IM3wRJTooC+AQmfRyJXpeVNGMEjV3UHMfC/9JieDJc2cvYJfXuhXQCfuHpssZ7Cg
Ezro53NTXAPnu8qne40lXvcqPfyORONlx1FdnVQHS/auhMteMZHTCVMRgrkskPHG
SAS9vswpZeorXoQsM3AZvo9zw2iJWnILN7QLs1Dlznkk6xa1CYUzADtKzObjDO6p
6YXzA8VYibhXwMZCd046dgMfJRu6ejX6CrUZGAnZ0UtwXmSyDNtp56drb0PnmhdP
gAMpGIjkrTQY0TRQmI1xEHsu5RsEd5/bfR/vSOWxNXq8mxEl9a8l+NkT0oWbKISK
jkvQo9G76niZVYJuFW2+q+5XGEB/wfXA9QesB9aAybbFWALme35b6n6jRFocsW95
0fjBY0eofAFffuQikyqDfTmQY9XPOZEh7CSJe47oxe3QBFYHBNHnnNxJD84zZf6z
MMygYKHeUY+YmlMUMbFSQLxmPwnvctstV5IIgWtVV3jL79/Ej1C4J+L99areAhAi
1Ivjo4h/mp+rfA+JsOoNcgy7ryjqTVgLN3gyNZZ9+DiqHKyk4mNXhcT8wWdyWhRf
+qAS2q064H2Azj3P8b5TLXrroGwwi1RbDueBA9cjNA34ZGC4a19eVSyXTQYes5RZ
kjBewuXOV/xHZMxD2s+frBXydJ7dhY/YboEFevEcdtn7UYiBi2CQh3c0y1+lJEQu
5HkmNAxzi1vY0apLWV6Gz7/eVUi5x2Tz8TnofJhFduMU25rB4vgdbnBewCbz8+Pi
Ltm8izmodBqMYa06bdUWyJQjg14gGfqtTJkwBqLaCzTJRQoEerKE0y+YlbE+rwCi
wDjTpQjKx1ikWOm8+ppnrpVK2NNTOTgw2sMuGVcmwWoYI7Ev/SDfpmHze+04vp8x
teuL0XwcNoV811RRxiVLS/Ye/bXJJ9U6pnbRAKsTLbWR5CXAl8EQ37iPqUXDG176
u1YpB84gdMUmPL7dMAipwz3QTZ/aL+2HQuJXNBkrfM6djaEaChPKwgu7rIguL5WG
bHvvc3ou0lRcgbN7lfLPY6vUX++B9p/EPur5fb+LyJvgUd5MAmFcvobRc4C7bP8e
87D16Gg7+1k3d5s9t8Ts+TmNW5jYi8NnCKbcdwyUckmQnbsUxoIt0Y0/ESEg3QQB
VBDT1tbfgPAlFanUdJ+e2OP1G+1LUhalDOtaqssj92sE+7CCxiwgPb3DGTXjsRtc
cyFB4vwE8nLAZuIps64oRjsrh90Mtl6DViW83hdhpirLzpF6VIidfZ//HddD9pur
4ah4BRAQQ2dYg86+YPCIGozPb9h5TgZv0ejL5qX16+HQJNy3dmphsI8ooqhHb6ZH
M1Yc1amXoOVprvuShfjVtol8NjyNT24MmQSvqc8SJpkZxo9jnnazMdwUYDgfewI2
j8Jt4gRrvCkV9isrrrEC08hh6SzK0fYLJZJkFIpD/O4sDHjcJl3b+GbbFDe2CSk6
GlWQyXnjL9rFfVIPyuUDjPh/XimWj4TEwRwZAXbhdE2R9C3vDhbJuDQuMMScA2XZ
KRGoUmJVGZuZwW8omw4fnCD9Zv85zIV/FeTLP94EYAbY86jUsW3IXKw7EZ14tOCw
2iBOjnPaXVKTJgj0fToEdKBRzS/4uW6q06KLnRqeFHT+eUkScuCcoBHWm1kEEHSO
J2FYuV1HOE1/lJSBVXKPKCV0rgyvUM1E1ST31T6x6QfhZumCyuxMgHxFu4P/EC2m
FT6sPpWK9zsNDmPrbT+mvwwDsw75xTbv2GIWitD78e7OBcnBP3U/RS9SDgnNbua4
HLH7+5WbScHamR+ggAw3vc606Y3Q59Gy4HKldb5YPB4aXBPz4rOmXNpakHS3QZFQ
zx1JBYBq9yQTkktmT1DjEnijNdqaWs+r1S+dA47dpGapSPOwvltqRVV1E2OjyG1H
GzDxnVHEA2QgpS9YDJM4g7/aGYU51ETqjz0mWl2kECuIShrpgSNeGkI1xXo0RQ88
9vH1X4aSzpBnUeHPJcVOAA==
`pragma protect end_protected
