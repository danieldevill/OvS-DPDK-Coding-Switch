// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NZJ/K+hsQeMqZ8n5u8kq4hGX9ZIw3WFC2ROVFH4i1gPSWcNfrOb+XAiw+WlgDY0S
wwkTAuU6ka10GAhZo2kS5Fu1C4sKJVKNgAMfWy4F5za/EWWmNLenxFiKyCTz/8KP
7EMD3Fnr/oTMlHGmFHy9OOYKsbovUECtzA7BwPXh9fo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2976)
TTCGtEZuOyMjlrZkwCEJHV6B6O6hyB+d/NjzVkntbva/6a0/PGF6t45gS19Bwz4r
VccP5x6rPWTbpGthLG9LZSr5lrC1LsFS4ibcDES7DtlM2gnuU7ifSz3//e3b9XUK
vcRg+g7GvtELtQrxtP6o2GD975YADtJMqh9EnYWh0cto7nwzBquoLdRbu+XJrKrc
N2eP8sdrlOryou2kyuRGSeDn+Ul+PpUPIoedaXkE3USKKZevZDe9TJE0zOt7mjdb
ByBE1YX6vwFGYMnzu4V6pEiAjd04rt8LDFzhxH7hS7EAALcS5mGTTaWPqZSGmVlv
YGbdY3SV7+qID3quuYqTqLe2/JjCS6oeA6Y2k/003EryTV8BETQWUk9gjNznJzQa
eJvsH4PNVB5SJcP94AUI5E8fACZkyjL5Q1EDCoBu8/q65QEQoCBWxEbTzt986Q+5
3Kp80FPSgtF5UtzoF9TatU9ZAbLjKPblVpBKWz2Y8766gCDNZaoXP7fmEi1YtNoK
5snd9p+nGaKJZsqyR1j+78+UV4ctOL8wAbSebzXCUBn6T57Rx0jUm5FzVATkkSgH
pa3SvRsQSiHVXr0/ZCO89kE49hGCoG5d3E8e/I8GH68U7+NmQViwJvX7ld210dBK
E1iiEuwKSeLGVNmzLlihSmQydL66/9u+V19Zvse1NlfW1tZWYWSR86rrPpGIZoVD
iFRGBFWxDeHnpFUh30OmLrvBA+48xGqJJZtbFtSpjn6xnY6qtrrQxxm//UvQYCqU
l91Zlk/nGRAOaPVXkHX5TaQ4UaGjbKgEoXV9N3SrVytXCbIr8bR7YsiiqWO5wT8e
pek6jNVvG3nVeqCo8f4VBgjSefR5nQ+onMZvYHCWtxXdX7fXpSsLozX9EEGNQsuj
qH7mDbL2pE6nz4QyNL5e7flCoPENrcqujGwKDAi2P/qL4CQXnlyccbxKR5hSBJP/
VtSaTW+7bj4soyoASZPJ3me6lcRNPO+etRK3V2RfPaBIa41o+kkiUffPwqg963lQ
ZfFxYXKBhk0MpUTFuSeujiz3dEXEHot7YFLEg+Nkx1eNwwioS6y8qt39KvRXqXFq
ISi1pYb6JySOR9/PVVxvsArc6YdM0s1SLQ/O92S98ZgmekrOwMc3HIGmv5ONKDdF
JMBGVYr2i8Czum7m1k4T2cV94WZ0aOlbuJkEeeZeDHaQ3CWltlCcaPr10CjSa2Ie
2e1PpAbe9UW/Lb5C0rQ9tkXj4rnM3I4JoCJA3GEJaP/1FmV1nHrHHyC6lftEh1ps
kGyr8Dc9lg4wfgtbqsb88DbAKzER479VxTjN38uuYe5rtVeDmgSnOnqjnYqnqWEu
OhA+FSGc2OiYdiEGZAaUI8cdmY2hZeRF9Mp0edStc7eJV/8e1n5QHUTkRXlCNItg
JwF3wt4nsoFWs3wZqfZP3qfti5XIaM8yKZ+WB+MB8tRqdGvS7hnLT4Sw4omZF/hA
bJVHW20iTelBki/9QIpxpYNBYHoid5HB9N2yIlJ9F1y+3H7U+1Xw+vpgoath9gwL
XPAxvpovquD1xOpl5Zipx5Fy+pTSzDqSWjJZ/3zCeABVBYDtG8yR10gL2GzkBONP
lCS6vpfqdtjFfdksD2jGiQOWnYVmkwvaa9jVGS9ij79gi5XGkeRy3Eyamwn+Bwe4
rKQDWHZa+IkwI4PPm3PGdQdaQrFLigbXCxpfdfdmQ7RQo0zL9AJrT/Cw9wkDPrjJ
HyyoZK+eZUDoEJISNrDRrmfv0IGKPoWqv2r8t9oe3BUavmBeUxzLd91wgs8ZzDiJ
4LETez/BU0jI7bJ8bBYikO1b2VR7Qec7/1zNU0LOutQD5VsuuWfdB9pajUBnprCS
x72g68kRyyeSK6aja8FxEkBn/c/RxEV+U5E8I4Ysf8a/n8JF4eQdFany9cmACnBj
8tVUO6BJexQH9mvbqt99rijXscvSCdkBJh+W4eJU2Wuo/xRB4sz8TOOQ9zDfN0A/
cV4wz8bHVkPMcxQrjRHqMYhB4U0SXW74wL4hmL8aOfhbUQhxyqywDornLoY9FtNi
oT5yrcoIB7ruMQ3zuEH9Wuzm+7Yh/tG7XKA5vGrerMv6DGvNmvytZuz7qONYVvVw
pEl+WO9srEMSqmW/2xf4jXi3cY8CVzZY0+v5iD/wQilJAtHPnL1wD5gQOVQldbo8
QsqIbTzqHgHX93CQ8MRFEIxq+7XuIFGGv4Bc2wRaNknge41+lOg4LyqEVY65tUdx
1ViGknFPYZORP57mT+H07bQXCiSRN2Tz+vS8zLhFpoOhSV6o3H2IR6epNtLUXpgg
pKx/vdeTk3ZzzU95iirfOxb4zB2KgkIrJmp9ptaR3gLrCPDPar69vWohoxVO/V6D
X4VqB4UyJbfjr4v5ojfTCzqADW7i1W8Oa5vFwLLT9nIwy/8cQFJZtdqdHxRQM/VK
4unNu1hDCSrxVOPvSzwMuDmHYD6zxmRhrG8IImKKraGNwBHwmGwauTQHyWaVBfoq
yVGKcKWD2qKdn/jsPELDu+aBsSlZxjGhq+QhedMf182j6Q4Ht4ukn8LS4/i0JqQe
k2MTUvwi5kRsvZPHKkeOymQ6hBOmgtO9Xl2sgxdJecTdz2YNfDSWCBiIfGwJ+SdE
7bBMV0VK3e9ZX7nDLU2asEJw71sSY52ZMWCPnafP4ly0bHhiU8KKHmc7sT7EY4rL
v1I27IfTfUDNXEMNrEIc6xQvXaFXNNOQInrQMOGjb1s8SbBXTel5q79OtxMqravN
D/N4PFSIhXB4lVE2yqmAK1q1v/5enjAEXsGB4Uz4mPhccnAiJT/+qPovacZ2KJZo
GQnE3+oTMHMj6FGekEsW7BaZQp7MGrImnoNRN1Ua6QBS8ACT+N4vFyNK7+Ywtd1v
Cm2rHUluPNRE4Z6bUMwBmW+UU1/S4ba2yaEqpMhftM7ehh30QAqXgJfAz00BWCcP
KxZ/AJGhdDIK1iPX7VOsYjbeLEaxFWa5M52pc/KrhcoJ67bFC4v5xJA/oA+M4/sK
ZHA2U9S1NxuO8vqZZUjuujHbaBMstamQV9JfGCn1UJUKFNjLrCq2O1jRQ1dVtUVP
eCbHLovsKjj7gE2xQtrkMX+7I3yZ2vmwAtQxyugA7r/TTbwy1poTSKdTSXTqx/k9
6hSdBiTv3ne6n8Qh75eXWSPdxYZoZo9IK5zRwQs7Bj4D/C3YAoWq3uhm9MSkcznl
m4/Ei22e9f2H/bf6yNShUSj2tY1ITd5lfBvmvqEsHfvphI6e9hWesG7vXR6V/BNe
rRqSF+yoXhOY0cCoRoHs3kF85W3XOGLT/7EaH9yLUxQ7WPg+I4F52Ar4w+hWVBqY
llLi1l2d/1ouqCYYWZjibxOHcvPAf+WvnNvrxAfc+TvjTSoChmH4n6kdxFAKbKE/
G5hHJ4C7pjao0rL3PNynd1WUrRcAWISzaFJ/NQXyvG7siI5YV5dB189aUU79v8UF
PWCpfZnuZ500dx2rnb4XJ8qlAEN82sjRWwt+A1lK4tk9j1YcHz6FwCC2zGBMw6na
EDG3HEnr45ZHNPY5FA/VM3wQDDPMWSUwPIQ8/4kQZdiAFGg9ldtF12uFi5xX1Q28
PRbdLilgPWNgCvVKRSl32BQViozCU+DF2g1uqaJvr1SW2tZ33sIUOZ1Gggsyylbb
KY30f/XZOQuHsBzGv7WNRpU8LUbQTlkk38hFPIfL85Vj4asBEvTTt72/y0tM4j2d
hW+5UL2tbosL+nj1m6snOsof2DIrydmC9ISdHOkZZkf+F7R6kq2Asbc0Y3ukaorW
NBwqi5c+Rc6RuIOsIvGgPWIdrEq8b6MORRB1DqXOzgOji7/OrTunuQCpd5Mxevwz
U5PPqMhTb2CEhv3+9GwV61F1YXlnAoY7Pcc2SdPZJ6uYOakkCtLwdkXORymXrCvU
DnSR98s4h3+eFzo+MZ9D1YHD861QFkzh5jKVtp+51EKqPVqNoG0PtUwkuDOp5/su
`pragma protect end_protected
