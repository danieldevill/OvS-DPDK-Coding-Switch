// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:04 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WrJTsPCXbGyxeIUpd9DC3jwitTcawRm1E/GFKib8qBMCFMrVkiIBr0A9009MuzWX
4srbaTr7PKENGMF3qwuFMyuYA18hzk+VknB0xHXaJhalheEoym/IKhSZMl/MGMwJ
GC9f4uVdteU3mxeScTOPnyEiPVPBmhrFTauFFmo3/jE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4720)
rEUL8Uvo/q5wL3fItBuLiV+5f/0DGrJKokYCtnng4AveMdLsGLbgNt45NPMfUipl
cRChA6deghrWOnjBKaZxWVypNjOr/zSMS2033+4S8+mPgtOMDCGUd9R6Jw2RzOzA
si97Jox1txVe9O4TK9sHOlvCSW8tWmdCP0oH3ghJwMwsOFS8MIn2RxLsWKrmoB7+
QnvMaMtydsXc3sIRXkw4MzAC/aQZAZ6fiResbnRpQepeoVlz2sfXUt5lZEE3VGca
mLR25c65kJ+CSAnfRJE+wjDonBaTOn5ebmTOnISaA/L6bjr5rnRIjL/NvuE0J8ao
Nf33jeEjRcxE7MrP28hwlhWY3fbmOJ/6veJPFZOj/ZwsJaqz8D4ev1vxPv6abvmE
2VtffyGwwOTk8rKnJvMncK7YcrE9v3kZvs+jcsUWY3RwygqH+NQPZnOuu8UuQT5a
1QsvnfGsN8ny096japYJxIDCp1wfknY+5c7cPhpqQOyuJuJHSvJAfYpQ7sWHEZQr
5ZSu17/VVLJcD6IKDXcG1azNeBeMR2H99/XkuWG3ejQk4Zg0mJOc6teVaf6ymkjB
BwU5zu6PNidha063Km8HvWiqH7oGPUpgWoOL+km1p19DyUHmNPH6kkEJgkPtkPEH
X9fiZCwHgwY5WW8Gbr93GR7TRep8W+qXj55TLSbde5ttMvuW7nb0RHrVstu70/DU
WlGf5CQTIRsTc9HOXmKLXmao20wISChkD0I61fA+d2fFTQofDVsD79suC3MnhTfw
8qJ+tBwxZObVl6NDYShQYJZbrcmXYb8NUDFnBdL7SKsjJ8uElKnWGCWQDj77tdHt
043YZVqjGcl/dGBnySxIyMRetszhIxNHXwSVQ2lTm8LoqSxXfbdupGb3LDWLZQ0p
wdDqOUyr/ME74WGvnai6Sf/dy65Wpadt2F+5+A/kFtrZEAwhNWT3HemWO+qaGjMr
5Wt+4H248mVrbbAuqpZ9o8waG/CdHijXwQj8D6R39I9jeWewDVCM0jpdgy/a7KjS
hGy3dzzUGGjosA5rLdc8JItusyQKLsxbvrd10dceEohGAvtriku0BQGWEkenYHE3
rQm1pL/tABPr1XnXk5cncqHEhYXfUC033sXlU+yDt4saIAt0hzcfWbRVivmNJJ0v
T4rGySZrJY+eCgYwSfKcjZsMBrrDwMWj6AINkoMMIOL7EBUWwZkA3ExEe0FS/qkE
LJrCU5mwFx4CIWBMC4fBk3OpVtH7RkxugoYBRHTB8ufB10hNMZX+Lov1CBA8P4mn
wf8P8oGy1fdXnZpFc+eLO/HtRAj1JQf9rQPEPUTsuthBFHKbb0MOPUkMoqip3Nsu
/2rxCgdHgcmGXdFKCHp6N8Pq1AQvOUjqy0zLaWDOMk556jPG6479WQLbVvf0nQxC
ahkND+XGZdlJCEs9CkSboDxFRmlThc0LxSXkvcNyD1K6dQE7+a3IDSAE5QFLwKuC
YNPSrONEgEssueueYGCxSFpZiakS7ixqxp7dRZDX/QqwEY43Y83PpI8z+VDm6EeE
urGJbGrT16iClp59js+dQ5FwJEFDoQIPaVipMCT3yGEcs3VhZlZgx4uU+SSmypbK
7TeCNsQdywIOHI6lvyV5xdZPFn3bkHQmrcuLzM6aikumhxjP/t0vHCCosKrnSgNs
Ae+i939PFE5eHUeFkL7B6e8A/UIbYOuSnciV6tsRd7M6d9mLICFGB4jb5oMpBrQ2
/LsYApg7IHnwTlME5kAW4tOyQ3tJHA42Jplvh2gWDZJvazhsa8zZoT6aYbWZj0tm
myA4NEkgkKfueHG/VDV/YNCx2WV62FUj4Gqtl/3c9G8uC0QVVijEhaeaeayqnl1d
6I0UHvWFaNd46d0qBdF7hsYamkWKA58OSNc8bOULQ+O89YEIiyfwXVEYBxJczirg
IJM6JePBoYBkx54AneJ7+/RJez/h5ymqVsAYvU9FpvGEHvNKSi9Lwp5F/569ug4u
cEmB3sHnU7vJ4QEK5nGM+dzgfhzzO198+mR83Nz+tDXjJVae0lUy2IlwFyK0dKv8
oANxnkB9OYAXo+rhi+vxTVTHb8aULw6AP8d0587o+g9wBTbpqCMxTpRWNfehxQd2
HdUMQk1efdIxlSqFYJbsQlGg/udC7ROI9Lp/iSrkoH2ZDXWn0YmmfcQJxJxeO0t7
3ojNROd8zqeel02ZDsqbdvwBc762WPPFgiNqwriBrz8lICVqpS30c22aZZ0ybyZ2
1kfjU0+sA/XcDwZQvMe1nFfrQcenNcEgxQ3/S4Aq9F44rTt1Jqd2yoL9IVoDQPVL
zQ54NHILUik6PvhzcsmjZ1DxJQ+LSyOgFUGfIBe9cPAp4yXeEc6ZsEKDh+cNvspl
RvlezFwlaOFZ2cb4zW7yGd7YyUHQd4UNlaGnjd+HfCHxbuy0Vr+uMIBzltw8e7JO
62wpG3I0MCPO1sYbPR3K60Ro4vLrwY4MBDo+zwMtBrM38benz1NjmpY+vrt7ZiPG
1zaPEnZj53AWBmUP6Ig6KeoltCirUTosQ4d4qpAGtolaLhCF4/RrZf+ko7fIZWkn
j/II0PGVvhy03r2LdhJwdAnDi4w57bEuKsDh3Qf9dYaGtb/O2+x3x22synkFO4AW
GGFvQ76Puao1rhG4id84DoIPmggq7U9LBR32eKmvQ26UOaFmkTUJsGK+GAZWjtbd
tR1YEc/GDgMf37lPVi6TGj3S7Kh1stKokku45V7iNAyQGwL3mctQwdTDx0NbM9Ms
/zQcDluS6JlU3AZNVA709Xp5EOd3S0Rk3WDsnuWqaDPCCthdoe6H50E6ut6AiCov
S8NapJvrT7mX3ebjzcdIJHaWCJbZjjImzSQJ9R+6YRurJJGKeqIBPV8FwZLtZvj4
MjOzkpiPjCCXetTP41LRaixTcqYxO48GVZ96sj94YSTibqPgbw5phw9wXyRuuo8G
fKdk330OuauXLE7IqVsScPIu6mY8kVS3vp7diDiuFHdvPlRNNtJoSJCe3ulghaAU
xLHjCyyyR7Fh2DFbVSrwCiOVWHVu6BiWdp7lZ8/Z4fCqr/jD8oeRO4tqYcRpp8Mp
IuRtNTGtKFgWMwt+xAm0b6csreuA6qy/zj0UVxY2O6hVfFXlDlkqBSfl97pJy9Q2
05wMooCSsRJmkZOdxLSl4Gxhcd8iI2/Eh31NznJWzoMELImARLzCqa/YABmnDyQC
jlI9d2OlhDe8abz/JWCq7HwD+EJNpJRJ3u+P1RrN6uKfnbY6p2S8keuPyL7z8wDg
30jt24KcOnuiaIzbpEjG7WSNekY6j0mVqF4J4kwmG3xxWK2ebAzKlGXvJd48YjoI
kMHOc+owfI4MDh9+TLK92tXZAKXgyKYt6iUBxPXCaJQEhtfB/m2yw+5N0cuHYEU8
TcwwPEax//DQfFEZP2Uf7Uy7/w+IJDrxjrGyxnzlZsaEwT4XBs4XzJpvsO4+p3IZ
FYEDN0tS93Bh9Mm8LOv8zu+2tuw0e3udkPJZyogI3QTqSjiZLj+B2FNfz1TRFEwt
KA7tc9br2k+ulwd/BpSIwAKMpCjoWoYNz7AGrKwOvNw/vJzHB3mtLiMltueAR/wR
uFPzB5szk/XCIF8WB9XjiNJahezm5SP2l7PlBKJTftFd0X3E2eXD/OgTpHq3DaPA
azNXfcdjt5QMCmcHTCLoqiBrnQtiS4mCZ2aj6yAGo0BH5tODcDVU2NUqhZlV+3ml
QMiepRtrz8QgfTktoWLlNJ/m+IQ/7w4jJklVDvM8+foCliTLdakDDYOkDC0YLjeo
ZSqnj88yEKTFHddxyJ+ThX4qQIxzV6rrH8CyHfhnWdrbKP+LO/Z6X9t+hVxLpRnQ
cfpNPOQo8bO/DW2KdaSA+TabvVUg/SsUtZ7tKobKba4qv+2KMRu8WcyMTk1Gnikf
kIHAcmWxrmHUeoypUmXWrbof3YHCGcV9tWxw27aPg8a5fV3RH1XzRlovgpRKuNpi
tfBuSRSRJ2211OX0Q7vL+epk7/fzf1Vod80KXfTaMvGNgT5JUP6bzxqzW3wWim0a
/RPhmJqet27wN/xg+qmQSEBI1sbQ0g8XvUMA7r9Axp7JK5mnAsNw7cZe4MGnd8yE
/zxdE/0XlhKziZugQ/CmmvzJZKghT48egxB8YvgaOcUfjIzpmi6I1qd9THXr/ClG
H3K2XxllSWH+I2QQjsXUosH3191LnPlhS8OXtclIkBY/x2Cr8U7TRvzbQf3theFl
xkW4SJcC5481Q/iPYuF4UUoXFXkS3N2kHO0Dr7z8I8al/0GtR+o6PeQ8LoMgaGXc
XWdooiwZM5kfRwb1ivodozKkIQaS76j2UMM7ij9l29vMp7c/JSfV4HdBJDsJjKhD
2vDIeMNAF43JqC9KdwaAhcd3zFNhj5kxZ88vZyhIBRRsvLz7w3Ouk5Sn1xc701cc
+sjdoh6dZBkxla6E1UMUxE7SvgCAKPmSqjr7Wru70YjRLR4vap97vyhJmyBk0dh7
DmUDYcPIli4Se9CZy55WyJVmGyyvcu+B6iIrHVjbZjqGrY6WchRtqixnPGzN8S6h
3tqNlP0YNQ6SvB2wrnVQxjzziuRyxV7LxYDtZq9z14UwqkQ8K0pRTi/+itblMxzs
/fQ84rRzn7cRCfhYMzbJB8pIjMq46LBURIERSSRtyj2bWXnJ4lYSzxC9TPze6CP3
KBCxSlnwiTvBl47rOHY/5nv39K0AGe0Nb2WOkyt5AjWzCvB40646i8SSSB+905z8
qovyhM9up7rykYRmGXmzIlaO8PGk4xoQHB07XcoPOPsbpsX+y//dSgpKNxnhGYIl
qy/pT4ctU/gNuuMDj6QFjzabOr77302cZKZUAMomkU+tpGDchE3WWX1i+E63Ezd2
ZIuEB3/v+sdGNIF/89rcT0MMLb/3xiL0JTCWimV3ZxGsQB9M0cnkv1IgE65nvuyz
hMwbtjxma1UP99U/Rj/49bRD4ZD6yjrMyotRnUKuZxO1Pyr+V6FTUcFPboZJ4w2j
qBLSkT/QVK36pr1/l0MijnO0sY8m3wtBtEP4MdnuX7ubwK4I/EeF/Mfwnci5y2Jn
AJuN8kZp5l0glmR4NrTHq4ZTScoAVJMl4kGGqojpOHgjSCaGCeP68WT/2NC6i6r7
PBIoOze8aGomB7zMyX8Vdw/RJgqdX18OteHQdACYR4w+NWx9DsVeHd8NrZbs+cCu
Y2Ey+KmZ84nN39s9AlKzmts0sfU+EyW+YPa2hOWmo1Pf0vNO5A1LD0dZkVSw5Ecl
1np7ye7QflqErmApH9jJmUYsyX8GDfrboSNX095gxikQ647Ile8BnPi0fXxEQj9o
i7pX+mWOAZu/TkujEyhdiW+T6QHl8mTQL7Tpos2uZ0uwMTPK6WHgBGtTlRFiW12x
f38BJFSOYMajfhYEjtfYJShwjaUpdh2MQD9U8MxLM19DpRwgDs2qDQwCJi29gvPJ
qn+iOj1jipIiQSa6N4DsLGwTIxen3pL6/HE/g+g1kljuANVZyk4gNOxM7FhdYjEe
cvd2CvfeEp5fi1QcZeAiDqhHxr1W8vCIC5HwCUCHIvFivS7/xOY/ivGRX7ghBMDd
Dkk5Vk4a36Tw4XAQduwnW7MekWeP06T/HaJvjgYyNVdUxyUpXNOm4u3eopZkW12+
hEJl1KM0XmAOh2rCfMLoRC6+BR88I++NgOCxC2p+5JSsDdlHixY/dwKm68cHGNex
FfT3VsoVjIIiUvZfK7WDZkuXm5L7M86Ynz7G5ZtH1V0EeftJ2c+jiGfzwItP7IuL
rpyVaql3aX6zsMzYmcGeFSQGcopnLVC5Eh3GwP9pIj373xz/mx7GISPIo/FNFLGu
AMmpIakC+4yQigE2dPWA/4VZeLibsuAk3soEGkHIcLvi2VHeewGa5mCz/20rlKSr
iPtrxJJgaMrMelxeRlV3k1rp6ZbqvA154oeaBj9Ba+yw7r9AtwEvVuANRTDKFNg3
ypH0btS+4sPmp3NdinhSpkeRO+CWoxO2xjN8WK3LalMcW+SN7fiRXdy2NgabkUYA
NGOL5RG071RX7ZL+ejDF4gl2FA3CpKnxQqbdDZNLrajJOZHJZpMlsP2wTVpM3NGa
itZTkptYdmMuLVr3yaE9c0Zs5dleac6YPasEvKtHUBqnzPRmBtn2T5uohsouclBz
7cfsNYQQeooWk/WJweYUVMjX1xz/eAO9ojrY7kF3xxGK00NM81NfX3JNJmix15vm
xl0GqOPQ2xCcsBla94nd/Uh1nr90GrY2wFiz/P+Ei1fGzw6qfg3QEXbFEYXX9mCo
0FMS2Zmj6yZVaPRDP6Eqbw==
`pragma protect end_protected
