// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:04 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XSlXo1imPtBHVX0DmTDMEOGluG2fNQgCiST45ohYF8hAu7ie4b5BKJ3Q6T8RIPKF
SncF7HNt/E0D0bPbGXMa6g2HaSw2zrc/BgOISmviaNOU46dHN1bxcCdu2lDEMy2g
/nn/EukbcfU7JDRk8ebuEEt2O066FQBVjVrpekHoAjY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1728)
2DswDt9s0K7dU+kUwDkvmcNkLYnTZCIAd2kVBf0ayr/nOJvQR/7ykqM32u4odjvh
gMmKE++3GnaNvAGGLd5FmKblibnjcZ+M80q/vys7P+DBzaktS4IKvQBwQeILmGns
q8A2fZy90mwe9m6ZKdihFtX39AmoHWd10swQouJ4J/ROWz4i5k1rt1mli4wU/uWO
B2fcebFU3K7gcmpU8pGq72252iI+qBbAm6rA1keHse+xY3Zyvrvf2iadlLmn7K6a
Z8J1ZnOUu9VKp3tKP3MEBDJdo1tTlAXKh12EwOx7QpNS3mdYRz3qK5P1ALqaIfVL
MPx8xqnvJ4DlFC/Ww8DR1jy1kraI/6RWMxfZ1uNKG56tD2nt0dapCfaZx/heyo0T
VdX9ejI50HakCXwMf2i1DvssIIlXkfyXzSImrWbIR2QcJQLE5C2gM+uyDpm0/+YZ
PQyJy90vXBuxJ55k63Zhpfn54fYNexUwXtOmu6h1eXfvzNVw2giiq1ph5lcgnE7e
7oGnp9IbuILP/el5AZOJMljfZKARCK0hmFYpbxEUW4dX03IsIAtKT43T2WUvXjPl
QgTBUWQ65ycSCe/EMArabpwKiglyvnRQTdjyLVQ4vpTaWjolJ9AT9oeyWXugrDAo
YAHt6eh5aQJ7Qa6A/PLmgrCZIhJ/hqVTZuy0+BI15kAq7zeN2KTSyL8WyHE4y3On
upT6mBgBc+7T7zVY05IdH7RXhZHZzAPDKTf6V0mGTrMhp+fC2gfPB/1L6ZKPleqK
i50WFCUc/ravsh3NBe5xbrisnW9xiCg9fVoPMRQqVTW5UzXhZJin+kX4ubOBzEEH
+i3pOWmQfyiP+enqDpoRJXzX8crXBY6asMULaKLzaJbZACoo0SFzwPbklOtCxQMn
kIPNpC3EG4JuxUxtvkeyMAqb4fdr+9fzhac7PotDDMkTZqd3T93/j+L759oe/sYd
DFXXJdZAxrnj6A++Fh23qkrbFUwdBDjzxVk3VCtHFWxCg+jqgD/+3MWT9LFaEYX0
P/BD2hxYByFJqbDKzrhd//I3V+JSwvLoFO7JeJoZxtw3/v4uJA+72YhTyEIzpbDt
qFzpaBcrVJjNvYkTcQWE2NhvckzNiJBWxQsHC/poc/CGNGVHsmhQ8eJbgM4l82BC
CvZ/0F55YMRH6pGwRq6btq5QApyzjOTGsX/CO9kiwEVuZZURrWAI0ABgceNG/2UO
2sG6PeLOEllJ9/K0JAupJGtVAGMKWDYi3Kn9btoZ4vXcUp+RDGPsN7NVNXHt900C
rnI0ZFQlRrajlenVeIKYwAyR6ckdl7zAdWhV0g3qirp8IgSKM2tr7Vizrhirp27t
it3/cFjFsiDrDDdZn5aYHbeKh0I2IncEUCjv3TeNZLKvAgpTI1hzRepzfeMLFqf4
pegSLahF8QMTmoOl7VqA/O6VovKQvh7FX2XeADceViAtFiseXsWH3sxHDA2aTvgx
t1nXju0lcz1wI0ENzLHzEXr5SK6RBPlweQkuX2ppanNNJxMRBgO/CoeuGtZUaX+i
GKs12sDCNtggpY3msZ+w4CrlEOJiy81tz247J6c7Dr6p9s9/6e22wcrbi9ntoOOr
F1gnzz8f7NxXWwgh1mz2NLjkjL4q637f1g3ZsdNhNFD5YfZ15bJO16GmeYs/yuIS
R80lSGJiJJitPPBrabMffgNS/wyW6Qs/mBu1hSwrA+EC4Gvx5DNllV/PdOlyiDgn
ipYMkyjZCadk6pmYQ+kgXFP1qctGyFtbffFQ0/UtBwb7e2ZPocr69YyItvLeLgJx
z47SPjKstecWdcNjnH0VgBWGEYfS+qq1pe+fGC8KlDNB3pG0VnO3BT7fQ41zvKPP
tmpLg6Id5TQ9/kHc9C9FV09vSEzxwgRKRJR1w0PkGVqZnZlOCjZZrg/0hF83ZV50
z1jtwXunP9KbmFlEhts1bkFshsgCcOlBtC++VLbmPbfezjsj1LWBV3BMHNak52te
4TkkmBtB0+qcleBKZ7YyrPs8nN1uKq0Mp26qCSe5lAxQkaTf4evWxeNSY/RqN399
g14K0kkWj9vwZcxZpj58e4nmbWoSB65Xzzsep1cybqFmZ6FJvpmZq2Nn2GGLU6G7
02UsoPjHJ870bLf7iDKVpjsykjhUeIaaDNApKWOVBidSwA2x0oZyOlxxk7GSdPyj
nFfsfMv0tW+vGlWDwrXXCcJjOetjHrlgqf/P4lJrsaCB2gJDHmmIjGDKFUsoQfxW
eI8voXMHxC4VHflcJozoLj4JLnasLVIczbBgPtVVx6x5cRi6KGcNpxhaIzdsQaod
`pragma protect end_protected
