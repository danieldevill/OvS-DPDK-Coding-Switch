// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NctYu0VpVWSCr9DEHDn2TgVbMwgwPBp4BSSxfkIL2vEkSATzVFmTb2G/WrSHgP56
7BnQspd9gHVHpxN8dQEbW3kIaPkXeTyyqYsa05FoRhzZvazxCm6peEhEGfzmLgna
ZMSO7FtyqUZaPF45Z8RWZC0pv0Fayp5sYBYNkOw2Eho=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11376)
1AoIlmSr6ynDi5wB72q7iVk6ZdZCye49bN2uYLAheN9FmGRA54oBMsAd/eJnbeCh
iGcE7jdenVoEGM9OLFbrug8JN9b+5WHgm9SLPnLRKFZp7Bnckq2q9CtoBnQt+iQI
Y5TMy6UmhERliA/cqQl8V10Q4zWtkpl/+PezTbN2v1q6Ld/bZL5VK132NOLGdmxv
/N5ArIeoeEh10xioyxA5TWtqCm4aORYdnMU83ZmnMzhl0MtDFdgWXQ03CKYEcbeq
pWNpu/W7PGXFrE5tI5iHdcZr70MBEYNj7w2o9G4jR+2LxsV/czM83Ge//3poEkcq
uuaRWI+snHMBfjCefE2LJ9xJYdhX/RNoe/6Pef3h7aovqKfEZRYBVJAapz6pIiqz
gZO3sX68n5zhA+X/c+KXTuLBKk5QlpfPBVc2i4POiIlwm7nHVuJdC8aRPgJi6Kc0
3Rhq7gbMnk/Yq5E8h0loSxP/iTKFBnJ0bvTeGrppVi0DBp9Y9myVy8AXec9kt/Zp
jNKUArvJjFATJb8XJaE1o65thFODDJZ7ySuhSGk4bWnJb3rOGXH7FZokg7G94GjS
mXGdCv5369rn6SzTVYAW6iKgBq+KL+emwmsDV59134SrWwYSHj5I2FLYEpgexZhr
IJvyam5AbDOw2/QSAQzIAO2Rp7zb1uZgjd1DBueO1uy8IG+UGM2Ik7AKXPxxbuOq
RbIyUPER2UFzVh7Ta6BeszWUtF7hYLnC7XUqnV+UJrugoh3ZER5p4VSaU3VT1H9j
cNh3vftasYhJteoK3Vu/ERAeI4rL+2S1NGJ5zkp9HUjS30kEyQ634yvLMjiKgRU5
gM6bTKWAA8sUVdl/fZJ7FyehgXOOx4NfRgqVgA847AHoWEUcaJPu3piiHgvcnu2i
63fI7di/byswPyIvIoi0EKEPr/Js7OvhPW/PcMJbk7E+uPWJF6oGs0+XWzRIl5QY
NLbhSrtgnlH6Zq2jAwTO+A67gdgLfXpdKAQqfrD+wgP7+cKTbg8+6HJtdZOs9vSe
vyRerynz5u4lBtENbIDXZmgZV2i3YFg6aWkv3dVpOq05Rqsvc9iy7g1hAIuvMqcr
/Cjx+phpeaY8R/d+u0R51SuU0LTd3JCUIyLrZ0QRIEfoT71oh+LDpXGbrAz2Vf1B
evCi6kd7Ig0mjJo6w6G0YUitKibYJtoy+cW5hNYW6xO+vAGzQsW7zHFpiAQ7mcaL
p0EsBxtvDDxffMg2SVMQSwrSGDDYb+bKLpzMFYtag040Q6jO9XgF+lMk0xNoUFf3
sMV9J0rLcOr9IVLK3DLPWGQXZjDE9xsuZXSHE5PBEYIIDB5t2p+6MqOttiG4Mvuw
lTErFjIJoe14e7FRiK/xaFPovd6z2D2iM0rf9k/UxsuxZVU/raZON9U64MLEtl8D
CVJy7e/rPKMzwhrgU+oaLr8LndC6ch9AAqH6UT8zKg0gtAZzA2gBRjyMR0ayT1Z8
eLHlfkw/kCC73iZcPol8gfYCeLK9xBqVe/m6FU+LwYC227JVgVdCPWxxfYtZWNO6
Cd8F57VH6oO/kkI1ukpEt0irPGhQA2BA0B5J6MLBFV0sB2EjzPhQ+yOO3EomORbT
dhJJHaYN+G1sQ58mA+QlkBGCtEKxH5mCxkSRdVgm53SU9gQqAWNqpB0EMZfWxP47
jCODGAXOkjhfANBeb2VNjpynSbzN7yThQDDUhjj4LRr8UAwMABo5Z3JZyT+Qo0Dt
9BzkNKOzDLJJlGyLONHhCiHXarZ3847hxF03VPdhmSqyiO7OEbVk1QlKo4rswC3g
UIegmig1PrdnCQKDE4oTly+nBSzIZZDP+y5JGETb/osZsuRPy+5Lvb99hIlxj4hZ
+86KeZZAyXanbytDm8sajH1QTc9lfCss/4n1Uj9BT50BNuqg1ynBkrlTGMKv3XPl
w6B59NgfCuGk5XPkdFTm9gLCwtPneRuDS55L6k6xp+1PFrHlyU2NpimalkcwYtz9
0nteGikCehuvHDvxaIUPisaGCixnTiALWTiFkfjdmOXUudtP0HgPu6ulgQdqMTF3
zOh7aJSPHxY7+433T+iJDMG7nmMuUDuJs2xO/cah3CG5MUF6YyAiPpdvfy5zvzYz
KfZMI8U2TqijxNUxIpj/pzZnpa34u+8WgPec95CK62uy6dM65zNl3/FUt3hlCNlt
RjauePLe0szrI2rexS7dyFslxrxVel2Exd9fCunvL+8bQOrGvT9kBC5Y7YkjsJFA
HSOPXKMu1bUPMThMWGkT0z9sWW7z7buQzWPaESMnsYoSmQcwF3HPHqE+jxOz7UQ3
9cumNclc5/VPa8nMXvlmRRWiVM2aKUHWbTUnBSjeeoy2ZJ/9vodvrvU8QNLTevDq
ogNXnX6Se4X/vMiavta1xvggX+xHs20BUBySrYyR19+ixGMZTGpMWwflEBo4mPvQ
mnInL0zCRGAUz4saUivWkOISpglynTgI5q9pTMko9/pjAcDtt65MIzCuLk7cPv6O
a4C45NgRvQsKklKWMtmVg7kyaixHqVM/gnuNPKMwC7TKopDWhFHK4Xz90ZDsA2dY
WjPOs0enuUgLovU7a4aPZi+cmOG+9GwJTlHeZXTtruEa7x8qKP6cjmGR3HgWU4bC
hLMOnHCPNGVTl7W/AVpnHGUlzU9v9KX+FvXqtOQ/YiDFTRkRvuBZ2jr4qU+vXHgf
eq6iDf/Bvw3V0AxbWLjFMgAyJpK9kqANcwx1/5okESpXcG7WDkoOUW3cBNl4vcIS
FzqgDbY7p+cjpoFyNmh7hkDVnsbtI9v+PqZII+/DWB9891d0rnZKgakkmoWTKf0m
bFBPZD71/gngEks36TcwwcYrxPpy5KQHBz7Ds/LK+LYdCh6sy2fDR/Y3WLiWvIUq
jhKlgAk/GM3df6djahTtcohlEdDESoBz3R+XIb14NZ5mIQt0I0J0R1nXsLuAWOel
atGhIG4i7OESxlroCYJbIVI6AMzpX7sjmYvr0VG8zJvkZXx/AFfn/HUg/AEYJskV
o9q8XEQ2ZmX1rrpYuwAw2fpJ8WL7ZH4IFc0YQ8SE4MK4EMk5la/fbYGrt3HsItKP
uKRn/BWebKs8bsCWjTdWCGCfCc9ATtymesOc/vcGsgg8a+u9YZ0CobZUkJHvpPgA
+TNJrqhX2X0eCRH6p8R+ro9jqsl5iGWo1rtFo813SwBbr4Kq+aDnwTYgelGektwk
+iJEJ2f1IucjjgVQ6YIsSjlYun23H2rCdDe8R/BsDKw9vkZVBH0Q20Il7gMrms6F
3r5/q43W+IptPtwrm88DnKm97NrJ5XJTynrOQ7XTCpRBwjE0lwGizGxpxREVc1gr
Y5RGSkLED1EftSCWGeotDJ3l9mdgTyFh2lh6v9m08THcN7p5LdrQYuZxRkUttERp
ZRNB0xzfcWwB9PrV5440FqPLCHFmv/yVB3Q41hNo+VOdyzeGUu5iv4JM/j1N8LqQ
E1qrEIaA3uNIT2ca1JGHB2PtGWwoKdUMUk3TmGkdBBpCMK3xdDsjGW7A13kNy0yl
QDR9t01u102qhjL/3rQ2mXc6Xuwh5/cwqdmBycpGF1CdDrK9yLJUw7Mbrhra42wS
iM0IVmesImUq5T8OFi5SBJSCGzhGbl7wcCfP1LKxFE9isTiJNLRV9M6lPa25T8iS
fIwNKNScwERPGavbBhfAx9VkOnJptI3c3OtfJS7Y6BgTTOX0qa4eeLIOUqvwHDEy
uKyJRzuf1CLDTs9/uhC57uQ9uZBlgszSPCenr088o0qmtyRYqoWJrywLb/FsGjmF
4AJq85TTascNa7fHIS0zISR5qZSl2U/KY1zy9igoXH/4PTPiYIbxE3v55XKcJedF
ILUeZRhE3nv8rMTVvseIAT4VGScn2hIxyiN0CRnTpwwFYnWL1Tb5Jp4ZRYMYHfiz
5y6T2qykfzIvtMvufIyYiPRw74TR7YFZM9DJZUxdOe0wVoneC2pNhVU58iC8fYFX
pgUftMmew00YA8+UNpPlclo3igVN1QZHadApRhl7cdfkiRi5ILpV8Jj6mxRkTKcZ
g8UitdDdlts2HFQizznnBFAdqr+c6LHDV/gRVwEEqEU1toPg7cMAWvx9dwKv/ER+
aRYyV3xfLFZ72wJvAniUK+y0lAqVKJ1BFkkajbGZw/s8CFHz0rHJWWtfnlUZ0BNZ
tDLQ0wZmmGns9oBoacC/lHm3aYwCaw93DBdA+9FRpxNg5OpTtOoYQ4cSZatqfH76
Wqi7AGw/grE4nOcPh7Y+rv131KR8aLG/hvuTnpNmr974yT3qtEbOdKlKYdHNJK4F
kw3UGQp2Sbsm32irwpmusEcE/qjtgaFXHlwpzXDPCXAvOhiEAO4uwZw/cDyW4D5X
q50U0sYtbOiL9i4zZqoL2SIV68cHkWyINhrs7qMaV6vtRz6H6TyIy2JGWVb3IJVq
Ov9Q2TBFGatQMFQfkMWhY3sKFzM7OYXrWJQXuA7VbzEOPHZ5ktZZzYUlX4CoNrrS
Pmjq+JjpKp4Z1vH9NPJWpmF9hWnTTG7i9sYd2NxaAOBKOoblSn7hDV/oRmWLW9r9
GMQnAkH1c8Wx3Wp32yLrr6v/AsvBTG6GTL2quIkQKM05WOQNRmNoPSn39PbISdSp
5v/089rrZx4m7Za8SEzdcNOMrN2zHMfMl8v2BTJWTBPo5IYggHckVr2xBTxdtFG9
pEgqC6lRpNT0XgFL6mgsSmyCQFqXpeU7LUKD7jmCJNKL/XH5294AWT9z9Q7W3IUK
s/VidYkX/N9Z53L3SHwjBOOL8HlDwxlmI+B3IQnevVGPMkCgHEYyva+IOib1vsQ1
wdKYFGdZAVg9x9DDQj+LCV1TDvVTkn3aQdFrVbmDBAQDv1Soj4TmPN0c6ISP3y4f
NuKzhRag2wc9pa5KkxadRibgLi/GYPCZV4/7UYMhctyqq1cTtDWH32W0yrsMi69c
qPpNZT4Vm1XoHCca6KEFSc1+4KWTGo5XlXiwEyQpg8AS3EOUrISi3Zi4uzlU8/eT
kFSBkShDfXxQhTFOeR/JbZ9dOrnpblE/YgBUUzplnHVqmVZZd73hBcK2FFrY0uVb
n9fHUTSOzt0VohsmwDB2IurP/zweIqHjcnImDG0xrHvCj8LST54a0iPDIzAL93Ew
1einfjSmNPwlZytpE517/F+nOt7H0MM7y0m7YQezyEJGaBGeq+BSw/xNxoFKwJMB
xOiUyQR55/ZsksOmXZBGI8ALtQmq/fnhomggZe+6bKrjGBaGbUw1SJ6nki3wYkI+
4kbIWGCuQeQgTCE6Z2gR1F7QLP9x2xhrbk0UTXrxPh5D/7imK8JKDO5nqFh0yv3b
LZ0Ud2OoaSPRq8BU27UM5nL+y+UESrMJ77kxJuBQ58QdA7c59cXxatU4K4ytKF0s
HzPgwOnTwbJW55e6WnKnxxH3eKA7XSi7xrIu4r3Z+FJGgaYwSZusj6+czK14RaX1
xnAOKQ7rpoHNQn/ea7RbNQBCYwDYxK10XyEulTeKJ8j9179b0422DrBbtHzYofOq
cVC+vP+ev/fddocSjG10mnSZdp20T8komhxit6YuJYPpjjfs42DPsv8LfN68zrhQ
cD6UKOZLzOKGfNxguVtonuKVzkEdf4AAgNQ1xnvaFNSp1CG7foEJC6LgTupLEwpR
lt3tEDTyLnPgA/xtAKoMjfYaUdAFIpWXoZSvfTH1TX44CSE5AbZNSLmgzKTgUlm5
x/rIKXHnLH2SYvdJrg9emR3e43tHyKxFd0ksyWduoxf7djNxHGfCznytHrtp3l1U
iAO7L83HYA231z2sNcGnjxrw+WyBVYwUrvISq1bXedMAPNYbtJLqnZ+kIcEqO4OZ
h20p4aW1gluCHOCXP66R9Tm7Nz3h7DdbT6g1QXcdAmSGpwNXkem8Adc3fECn8j/s
cZdnV1pghYBauyCMAWg4zel2BBHnk8+zyEcCRv8yc4KV82a4V96BbnmNC9UV6pqy
V+f/Z00ak4CkOsLMqt349bCMdSmaTGtCHEAkWicVzuuU/G/uOZbljrG4E/4z2YJS
I+9X8bN0F8N3oONOqL3pXYTurY/eTGAv/NPFw8EDmUvrnYSjm+EWhCi0DADUn96/
e45etejaaDGh51Y4jOVN9Wb8tDJBNIta7dmJNUfytPhCRjFFW/1PKrFX/jci2bpH
exroPf+efK3LSC54U1WEzW+RGeKyBzJhr1rHp8QdzP4wE4nCzF4NE6vRViATR/Mt
Oh2k2WexXlDN7w2I7psFQxuj4S1FLrFo6rsSDZk+SyHXwLZ+1+j+zrf5/lljv+Pc
/y93OEtvJ1VLbAZ2O9XBhKyP7CVRoaLsaFVVHaZD8rTWU11al6sTLdSBg01Dhdjd
jZnDzogH3DJGh0qz6OWarKFNJbG4cQspohMTg42EJT0rv4SUJ2ZV0KCKCZRvCD9e
2Y5WeFG2V+gYMIqklM/KZbKdypuuSO+6C9B9zOcpIiaroYYprkyGr4SS+F8lgUUy
rxm2YPJp2N2XfW5b5qrghjqDXAW3jKUTMq7TvbooSFVEt8YFM6cTxGSBl4cJAmtZ
bZq0DsqGLT3E4KEs2CseiL4AL02l9Nz2j3JYyul2uYtuXeXZsPzYOCqu6pWaXt76
dfosRvryiiiyuWD31m4ElrpRAI0MuBnA2OF7KfUdgQGdVyDrwy1K44EVm2hfKC65
tnDvi7bR0g2yICeg8FS7oed1hUAOp0uhabcFIQs0v2yH5VadD3ZiQMRzgBGQ2hiZ
PLR/wrFUMMkppk6CTRuDec8Ve8q5UVPcyC2RLwYMsFeL+3db7ttB0/NTZGmnmjPN
g7SXVvHGATW64tSHUarL2BjQ+RkoYkZBLTD12IQnhVoa1gVM3mxZoZYdM4TvCm4E
+YlXt677wiTmuaIrP04wu6cBa2WicqpirbvzvbG5AKN6gV1uoye9y8SkJuK0M1zp
0S6SF8KbOEkBUIfpPC1526vzkHDGk4Su+OavA6br/QPNFIVbPCCmRXspnxZGZLvm
6emuzBnjfdlAWAe4jSiT44Zaj6EE4F3We2FV04XVboWMHIugIG6ttcJdw9kcl/jN
nolzGt/MhC3YZN3gu7Co+nwG/kaL8uRez6ypOWpObivGEUWBh0B9DHyAQGj4uq55
HZ2t0sNqvh6qfjWjwt+XbjxE6ctxs+IHBMURmSl0sHcEvP7CtrLWahDVLGZ7es76
KT443G5c061//IlBFC00Km0TLbSINdcSXT5YHuTA25AKCD2Y8hylbirMv1S4kfbE
gcAh61i5ooqsQAil/wpN+uXxRGCqYtL9I0wI49U5io4M68W2hqUDNC2NFg7ocxzb
jVkL/vMbVgtB4nTwCOGGiQMVJV1lO/Ek6cMiEdV4UP2HLhs16Mg5fzCRwhvOHhT2
us0O+IDWP1gdWYniNat12I3WHsx8IzLohmeM6yfX23AMpR3CdZjy0CY9lLBIZvfh
nk/Uthve1ZZ5wt7smjpvhwaciEbMegn+5yz6udp5ybSYw8snhfBL2GwApt5j+zDG
/XJQmgag7TGO6I9Hb7xuBeqNBuih8ryrE4mowcyWAtyf/rXLVRnhQ9n+GacOffsR
V+F1e6H1oIH4AyXLyKw5FfzOE87oAwEw5fC4PLLqG20i494w+zyoB9XjPacQUAm0
5RJokMAMzkkTIKHZKZtFlPW4uat4E6AhI5oblE5dbseXkaIeeFJZeRGRcEszyIIt
KffOauVsPVLhzkGh5bEIXkD5aXvKyfgqD2SPxv+4qg5BvsZvgTGPh2Zrr+PSw/3C
Taxqx807wqIWXPrQ+T+UPoWGvCFaq2P82BCTJS9eB4byZSuE2DgpbchHtTDtL48B
Z7ghe/FH/85B8HHx4IocRHkUgrVKH0S4k9Wh2EhxtOMSfo5uRejNScgnWKa/PC00
sXG+Q9mbbHLFfRt/CDc5GGS1M+gMK8EfDeJk/j+yd6u29PixZk2Ld2FLEdXHsium
72TqEJzw8Z/F4kJXmUICmS6tHi/TW5px2us41njYMfL8KG0qAVz6B4VdLCqbrTig
tGtAIJsUEqMjpfE31eh6LzduSL6SC1YEw06I22ThA+fVoY12+XUnu1X/R1rvBI3I
tcU23u8sIECtSOLwacZrlvokqV5s0w2yA8d6WpHtDu3OvO8A4SKpaNLeY1bgXyKU
wYKiqm7iMNbFyKsZ37AHv7/uevd858yadRTAfdj+TZaU+wwgQ9Ah8LXjeB0eoj7F
O/dX6fhdbW1PGEdbW8TekuqoXcSxAah9JOcGoQetnWl4cYm7G79qJ5HDpDRA+/9Q
jY8YANEbpP05zDSpQZ1vczN256cE15lGYcqWTbaIpM2kcM+N2wUk1uc55qNv9dTx
gA53sbJ6wqM4aVKthGa37CuybXmZebB7HJpp/JOhblD2rABenYyNTVRNvpNQO5nF
LYsZF3hkCUE+cnHy9P4RrcDqisD/De9hY0xvzrFBX6/E+P7M2TAlt+CpzWNDuocm
APLFpB0cZXA66FlM5tLBgk6fMQ9ZmTiZvKQX7H3ccYcyic+IzpczBwH/KbUYdU5b
RPdKSb5Bt5y+FQPMJSZcca1AFj02FQ8iTVdF4ChwQD9nISY5hJYQccu9n4LtvzoS
wEWnBRmqXGbbL2laZlcYK8rLFplpNDWUoQs2RaDO0Mhwl7lkfkLvk+QVI/qvD+27
oeEACMhoAU/+BsN76z6jisxV9ON9MqozuWN9SMos6tKVuGzpHUUp7TDkFNnCE0xe
1mEMLZDxyrBDpVp5l5/2kc33eWruFnHrGZkyvTHX5eCC686osHuhv1Qvahhr8BQf
Bxx4600rsO5VxgL+wsz6xCgTOScWKmQzZO6/T3qcDdDgYvJrBzHHLM/aRagNwJEj
6DMLb++I4rvTWTzYd+9jXar+SpvSiAvIoPUQsWba40bbpb7BAFQlEnf4GAy9puxR
xhYLD3EyZ0S9iPRAINwqX1G65D2F2SYt15y6feJOdBbNmlkLFePqrjVkuUrGsN0F
ew8c77wB1bbULbV3iQF/eCCVFu2yhXrAFKtYbgOqdGcAxi3C97vidDqvpZB9f3iT
1PRdlyucUXQ3HPwF+a3UWYeOIFS8vbxTvwSnfa5ZfM00/EdQDQfQNnSwYp+iJmH1
Qn6g9GCu6XwH8fWmu1ZOmVAQtUob+FWuz3tzaPgVssMpVg/V87ApcWu2MnscGhsX
nLMBF0UG3OrR0Dd55S/QstwD9MV5KviTdnYImETn8pizZMYQuvkfxFePxdpiFrpN
y/9jyNcJ3CCUhFXyTsfKmVmJl50FURCjkZjWj2uGGh2DJPVl3Q/C1jzYxzgVJ/Q4
IX6DRg1vAsVB9V0iCZ3FjCmcjP7hAoMWKqV584Xcu1r+9Cg7L67L2EbnZcBnFuJ4
ai70Odb1xNo36N9MTHbT++NNirf5qUDqEohShRXJTQxrut7DX6WTA03NIQwIjWd1
2qL/M3CV6yBf2DJuJAeJ5brUd6iXUGjahGr4ek2Fo2BezIlqiw/nkKsNWfM4WiEy
6aoITnzyc/RxFwqEx15SANTvicDwGZelcZe/pjPWgjg9wROuEWc1uhRskrAEfrR1
ZHflWVok1y/SiOibk/oWr/yrn94dIkvcnETvH6kXUnVtFEtH4Hc9p3ontzg9BA47
ZhHt+fCi3f+qPEXantHm2m/WUsD3B4JdVj0cuoN4NTNFC+XLyyKldMRAGd0cUknF
j5/FEoYns205Nk6UEmvAiA4TzMfdwpwAPD/85/UUVFF7fatM3q91yIpafqkbxIwn
Md4hAbHNtINZKpTnOW0owJbYDOJy27ZFwfMnHnOjPGJ5A27Ofawo7Ln4Oyt5tU9j
3temoNX4Us+Cv9Xw0+D/aca86LF3O5iZbzfF+sJV4jboknO8l8eW3Ckmb/NoSBrk
j8nj63jqvxO+H/aX8Mr1XW6dDGVLrhYM8pc7Zxg73LOB8T32z9FzNh+P5/yNTcDa
zuAYhcdF3MiW6nJIobdoypW/2ZVPSi/Hx+ET4rhHkGui8zUfkex1qRiz5svq0tke
e/cACvlWfuCigk2wfDVpVuHnBs22dnEKNUxWKCTZADEgvL5fZDdETvRNE3dZT/9d
u9ag+fELPw3GCAZg2E8jLHXZs1KUw2DTwOhv+vp+lEsU9YIpW/jO6wth5xxhkRdx
G7MWqleTe6pDsH/Doof4KVJNuX38yYQA622ld55svR8tAsTf+O5eNoQs8lyfq4I0
IRamjxLQXrFEvSIi2pOxg/aPjI76KN6aF/RG3iQH9s4YT0FoeZXyn/F2lVP7BCU4
fmcZIEK80ZKrsPeq8BXVw0MX+tCZcIaLG0+rfpl2jVcVNzIlBKm5B2a1Ug7zBE+F
faxMMByKd8ARLnx0ex2XVvvMQFGG19BzbuUZHWNtIauRI3vcTkphHjSKL2IoIhTN
iPsKmRpxVwlffpN76vPy1Soxl82DEuw6S/xLbmwDf0cbWj+MOS+bmRZUdsczqcN5
49OvJNiZEzW9y3Iwe5doQALQ8IsrfetA2/SrzSRkOYAC7gSHIvbyszfRIMH+foyC
o83XmCxKJYPhLnhbvsx+rKEbilMYl20BntjZudkCvWAdNd3/wYR/iyPwbvaXAkd5
/TN6DJJSObXeyI3Vv0+nesREPwQJM6Rzy+mmj9U7268v/Z/EL2HvPg+daD+l2HLf
GASss0XyWhM/C4phJ03PMRgvlr00d+R9EzdxEmqqiDCHR3itz/I2D0Uz2JFqqXKV
94Z5xgDLOcWErvbq+4TNXwFxh13chgHcN0yobeEcYo5TMkavyxbmEIsKlTT5agJU
87wieKsdW60vAurR0fwtc7W5CUkQwBgH0DwCk80lGFkyac6VfCUrE+tWXfRUIADY
Cs1ELB3TBAUKCBvN0tovi0CvkSGGZNEqCDSy3yMSfVnIHXvD6ht1onmyq2gBSGpQ
XtOaHJ4Zimq+VE0K2NQ6xPPPUdHg4+bcUDFZ3yw/SD82gL3TXJ77ZCtsT48XvZzI
fb5GPTuVcGFZq9fHC8fyROokyxODp+Hj6290dYWoc3uC3eB6n0lcWkiRgFgIYPWP
TmjLDQA157TRCjvoj9tzt0L3iC4kLq3p2LmuDFVHvmuwkumlH1S8aAmPmEejxLD+
CmNE0HNX/amSUQiajmGAlXohGx+Pm/9QVfMK5RhPgdLzZOSC0ujsu61zlEnmZL7f
GizM0SDvplKtp+jUuaeuBnRcd5XROKtFa8YkwEZwROMCJL0cH6+V5tjSWdSBa8S8
8sWe8sTC4bxwyFRWs2oBqGv41RKthMAzufm+AE+XrEl819C+COsmLysP9EnuGmoJ
oL+dHTbmVDd+maqOfy/PWwEX+/oq06z67KhgnPUdQMiswHW7an9Nc4L11SU3Koht
P04UybUDo623OylnUjTyBLn5GG2qqWx8STI20omPQbBj/o0wSRJ0WKtGFx2EHMeJ
7VBt7FSQUs9G5BwJp7FR/YcQLHzlke9NMyy/WSaaK09NqW/lQmy0ni75OPohTRTc
UUpbn+qOO/ebJgAGdfhBY5quzFTElJm0PTBEyELA7iub6oniGqhs0WEj8MNcyjsW
/lTJrxXVT+22Gs/cKsE1Nm+MtqILYwZZ0/wm9yRDgDjizviRMMoynWaMd0Uwm/f6
XGrijx/fpXtK9nYZ7nlYTtseihZP9se14CR7fdkwYT7MixKT2kVwn68TFGQUKX+q
pL3n6uwWNLjBIEVS4I09n7Nh5P9DCCs28FNUe5z53Wcwt+16t6MFrKlPkswDCj+z
Lr+qbAmAEWj2/WDDzzhwhsTRYsTEr2daSlNDsakgUNKFxmKQqP5jGyvzbZbLdN7o
E5dBayX+W8ek3fHMWA1ZLeDWgq+vPXtFea+O3H8rM2Ej56V9uCvpRoVXVPo3ydqj
iK6XqiEZL6i3Pc4pjSmWWZJCgkC2XIFhZbO0kr+4pimDfNhU1f6o5D3UEXST2ok6
+AgWfaxxiMOymE+ioaxHNTkdfX+ou/KWqGOdVZ1L+WqYh6TgKv190wRO13qEpyl+
J6V8mAGv7wUJOxNoEGG/l2eJCTeoFgcA5YSYksYw+n4NYw7c9zcn/Xte/bY05vAN
sJl1zOT6BDeqxH/JEMOUDHR7ggspIAinwJo4bmC6h8iGYJ18odk7OIhHEFVuorYo
3H5Rg/1kr6wW3Mc0EoS+sawOTE766hNocrclwIfvZKHsKfB4dW9ogXVPuygKxL90
KwDTseJ1UxAc2/8xBrao4U6xThFKbLlX031GyWoW/xLCSyCBlAlU6ANLRzuJVBqh
YMLkssp/zsvNX19MK7SFyLExuqCdoGaqHs7nQQlNNZ5vAljDsDEec8lggWQ29in8
NliQbzO7esnwVE6NSUT3JRdgxhwArz0qxr0TeQghttrCtjTuAet66wkhSyvq2r6P
+aiW74AJQaAx6Ssv6hOGTWre7AKQRemKyLeCN+kHx08sIVmz6ASkSMqdJlKfTepr
hLUJr3ID2c/3v56d6k1iOGP+JChDTIX1EYIAvf0E00au219gBU2eOjgrWofry1Ld
e6MYsRpM2XO/Jw1byePxH/YVxf6lyLPX/khCm+ClSjw9wEbO2rmJZPd4OmYLwGOf
AkoHC31+8h5c/sMeF1uRaTdtoJsnyPvFMFnjFS0/I8gCPFet++QpIgjB4y455w03
SYRL9EDtvCBv3nPYoMK4bN75bqzFUi/StCgNLNbFHYbi7Uzfn+5ABKxsyClv6dL8
Q0OpqN8aRfd5SiGtEVMKrD/Jptwq9u3qKWO5i2iIE16AVGq6Sx0hvZGo3F7UYFMu
UFZU4dEy3sr0aO9rquARvv8lxzdcC+/cPolCP+eEA6DNQ74qk9u0OzMX1yiu4CO2
DS2X9mz4CdE/wq8xdQrv0xVyHYJO9OQPLd+cfnGyZExvduwL4BXPbunCphFFdkMb
bdnkHSD5jUb79NsWqJeSdtbLnkaPRWXRi7ws1J29xkJ9lZGEccE571cs9bsnskwC
Ay8CtB4we/AFbVVF6KarzIkOd+q/Wd6guzS0oP5g8KJt4/lmVRD7fCjWvU9QNpKH
KyLvxvyAk7ussUB2OOLM2hW3tFIy8I4EeoIun/YxNCYxU/4FEwunzkeMhdeurwdA
uttYSeWtVjZobDwbQrlshkV+GsgWte7y+ZHQPC4E61syx3GYzLbhcpMOsdcplE9X
LRDcjHFXRgoOr8Kfk2XSrsOBQKvOoXMI5C4PLNReouYx/wN3L/mQqQ5QR2oao6B0
yqJv172eJ8BwAYEEKwTkadta4zuPD+CdFvI8JqZt6wqK1QQzK4ZVi9qxHJNh+Y2O
MbHqDdWH9Yc+DuNTYF6oX7y5/6bt35PC0A28w30FdOzJilk1iiZMzMFticrEA/wb
HQrzlyVn93VzSkjRzdSS/NK78UWLo8mmVGKc/dVoF4TdxZk/xhzkdzJXRWB1g8pV
9NuZZ2S2ZNdaXVggAFxV4tgV0mbiAq2zYf5VxyP4wjUZdk4UftcgT4xnESwy+M91
3wRWYkvq2Q1ZB86TkoFBV5Cd8CmC06c3lptEU3a2YR3cR+LtgylmupmVGAZcgxwT
hGDGNhIL43v8PTzAebof0E5EFOxOIJGLgbKBdVumdkktUq53AbyFVuy9nST5G/Oh
nLK7/IVMxqPED+XoXmQKqtZfIYSF0lfRwE2wTSghQuTyAcOYckbLQWZAxCepdUwU
4sRbad5jOrqXztk1yGCA3Cj9OyF7OfwL6iII85DJKKcQk+sAn5NsKtE6UCX4aZfW
1bKHWwYtEZwrjbrK55tGc1qJH+pXVAa6iSy6oHI/I98AspyJP9CHEAPqFCWCClqU
fj2krtqn6B1MmJLFvg0TkFX7firrB6pveASRCyM2FyECOKoh3C7xxgVpJTVvvf8w
kiQqY+wtQV+uf5xzI/1zNNM9q5CwV5vMfMadK37/X3tgMO6jxyUslu7x+xur7RGK
7rpRaVnSNEPHAofRx6eVo41D+w52EhxofzLOwXVRaSEGCMp7H9MW1GbFy11vBPfi
GpRJ+tkfkiue9u4jb181RnrX9nlXHmI6+Mss57p0CLvCBb7X1imkGXQjv3AE7LMG
Eah9KCsuNLluxS9cqpt+Htt395CwAg1KyfpijigZ2HBe2me+DAc4dqEp+DAIRMqQ
ES/Yge9BLBAdM1F5gX1eGh5/fDoHkUt5zdHdunwcsmIQWuGgfUKplQQMBGFT2FHU
38Ft5IbIit4VhVYTSPT8OxtBxLF/yWGazBm/awHgiTte916Fu2tFycJgTYXROI4y
+UkGHVjLv9zWyBnuHy6H2MyLsT/1OGWhsx1MJalMjGOjUZBhcCBM1v/HuuBH5ljm
XbuLNtIb8XTkCwTMge3UV3f0qlxkGOIHIqFHTKPT1kat98dJ9vGAJm/w6cJd25YV
KvmwWG7OEcwCNuUwuh6Lbxw/Xg6XeUlsR1issVtuDJLm7Up0AIfz96ISDDQ+IwZV
W692hAU9iibAOAdVVK1R8MATXd2DOFdpmnqlWlUECDkIL6Y8KI0nroB0cgnlWYDx
VUCYtFL20fOM/PW15h9fpQaLx6ZDScKgx3JLDsBZssNbSq8715wmFq2OZR5Fw997
+Fbmz7YSLWetqeQ18GnIOdEFSmOsaf60GiBUCD1n2iorL9Y5/XNXdLMJhVkomvpQ
Xd+LvWt8TrAlsJQHXqhZCussXi+h21SiE0Dt9u8yHZmvSWg1w0ss/bMxPcO3KLLr
6HYoxJYZfP0f5a2jwtFAdOXo72NmNcCG3nNacQom4P+d1f0xmiFMnriUpO60Ou25
ljLw1HQsV1NnLDuom38H3JD2d2/8+u5TCmZcFRxjEvuIFccoHEATMSwVObCbCEV0
P3aAupJeh/Qa3d5y0oTonUt+0FsLSB/HITy6gf99dnnsVRETeOZH3erz4fb2v3Ma
dgZt6aTDxeihOQBSTZ7qsifMVc1hQ8o3u4LNYCSRMZURxcNwupplYEZW5h2zbsA6
j7F4fuCg4/VneouBBFjbfOi9bWDhQNrpiMYuwaA3JWN8/2xe9f/lYjRou3S4IZXu
GR2m34RoThFd0EY6P+HYjcJ06cQjsnAYG36bxkygDfyEkupCsgVVwcYMmf8mry2A
dlIiYqOIfdW/rFyc2TYF4R6yday8weVxD9bqJu4qImcfGsfPc8D3i6K6qk6Ypbep
UmZCiW7yts0IcWLNkUwK52+t5cfs1LC4AbGxP+/ATKP77k1zptBJrFnjMAWyTzTm
`pragma protect end_protected
