// pcie.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module pcie (
		input  wire         npor,               //               npor.npor
		input  wire         pin_perst,          //                   .pin_perst
		input  wire [31:0]  test_in,            //           hip_ctrl.test_in
		input  wire         simu_mode_pipe,     //                   .simu_mode_pipe
		input  wire         pld_clk,            //            pld_clk.clk
		output wire         coreclkout,         //     coreclkout_hip.clk
		input  wire         refclk,             //             refclk.clk
		input  wire         rx_in0,             //         hip_serial.rx_in0
		input  wire         rx_in1,             //                   .rx_in1
		input  wire         rx_in2,             //                   .rx_in2
		input  wire         rx_in3,             //                   .rx_in3
		output wire         tx_out0,            //                   .tx_out0
		output wire         tx_out1,            //                   .tx_out1
		output wire         tx_out2,            //                   .tx_out2
		output wire         tx_out3,            //                   .tx_out3
		output wire         rx_st_valid,        //              rx_st.valid
		output wire         rx_st_sop,          //                   .startofpacket
		output wire         rx_st_eop,          //                   .endofpacket
		input  wire         rx_st_ready,        //                   .ready
		output wire         rx_st_err,          //                   .error
		output wire [63:0]  rx_st_data,         //                   .data
		output wire [7:0]   rx_st_bar,          //          rx_bar_be.rx_st_bar
		input  wire         rx_st_mask,         //                   .rx_st_mask
		input  wire         tx_st_valid,        //              tx_st.valid
		input  wire         tx_st_sop,          //                   .startofpacket
		input  wire         tx_st_eop,          //                   .endofpacket
		output wire         tx_st_ready,        //                   .ready
		input  wire         tx_st_err,          //                   .error
		input  wire [63:0]  tx_st_data,         //                   .data
		output wire         tx_fifo_empty,      //            tx_fifo.fifo_empty
		output wire [11:0]  tx_cred_datafccp,   //            tx_cred.tx_cred_datafccp
		output wire [11:0]  tx_cred_datafcnp,   //                   .tx_cred_datafcnp
		output wire [11:0]  tx_cred_datafcp,    //                   .tx_cred_datafcp
		output wire [5:0]   tx_cred_fchipcons,  //                   .tx_cred_fchipcons
		output wire [5:0]   tx_cred_fcinfinite, //                   .tx_cred_fcinfinite
		output wire [7:0]   tx_cred_hdrfccp,    //                   .tx_cred_hdrfccp
		output wire [7:0]   tx_cred_hdrfcnp,    //                   .tx_cred_hdrfcnp
		output wire [7:0]   tx_cred_hdrfcp,     //                   .tx_cred_hdrfcp
		input  wire         sim_pipe_pclk_in,   //           hip_pipe.sim_pipe_pclk_in
		output wire [1:0]   sim_pipe_rate,      //                   .sim_pipe_rate
		output wire [4:0]   sim_ltssmstate,     //                   .sim_ltssmstate
		output wire [2:0]   eidleinfersel0,     //                   .eidleinfersel0
		output wire [2:0]   eidleinfersel1,     //                   .eidleinfersel1
		output wire [2:0]   eidleinfersel2,     //                   .eidleinfersel2
		output wire [2:0]   eidleinfersel3,     //                   .eidleinfersel3
		output wire [1:0]   powerdown0,         //                   .powerdown0
		output wire [1:0]   powerdown1,         //                   .powerdown1
		output wire [1:0]   powerdown2,         //                   .powerdown2
		output wire [1:0]   powerdown3,         //                   .powerdown3
		output wire         rxpolarity0,        //                   .rxpolarity0
		output wire         rxpolarity1,        //                   .rxpolarity1
		output wire         rxpolarity2,        //                   .rxpolarity2
		output wire         rxpolarity3,        //                   .rxpolarity3
		output wire         txcompl0,           //                   .txcompl0
		output wire         txcompl1,           //                   .txcompl1
		output wire         txcompl2,           //                   .txcompl2
		output wire         txcompl3,           //                   .txcompl3
		output wire [7:0]   txdata0,            //                   .txdata0
		output wire [7:0]   txdata1,            //                   .txdata1
		output wire [7:0]   txdata2,            //                   .txdata2
		output wire [7:0]   txdata3,            //                   .txdata3
		output wire         txdatak0,           //                   .txdatak0
		output wire         txdatak1,           //                   .txdatak1
		output wire         txdatak2,           //                   .txdatak2
		output wire         txdatak3,           //                   .txdatak3
		output wire         txdetectrx0,        //                   .txdetectrx0
		output wire         txdetectrx1,        //                   .txdetectrx1
		output wire         txdetectrx2,        //                   .txdetectrx2
		output wire         txdetectrx3,        //                   .txdetectrx3
		output wire         txelecidle0,        //                   .txelecidle0
		output wire         txelecidle1,        //                   .txelecidle1
		output wire         txelecidle2,        //                   .txelecidle2
		output wire         txelecidle3,        //                   .txelecidle3
		output wire         txswing0,           //                   .txswing0
		output wire         txswing1,           //                   .txswing1
		output wire         txswing2,           //                   .txswing2
		output wire         txswing3,           //                   .txswing3
		output wire [2:0]   txmargin0,          //                   .txmargin0
		output wire [2:0]   txmargin1,          //                   .txmargin1
		output wire [2:0]   txmargin2,          //                   .txmargin2
		output wire [2:0]   txmargin3,          //                   .txmargin3
		output wire         txdeemph0,          //                   .txdeemph0
		output wire         txdeemph1,          //                   .txdeemph1
		output wire         txdeemph2,          //                   .txdeemph2
		output wire         txdeemph3,          //                   .txdeemph3
		input  wire         phystatus0,         //                   .phystatus0
		input  wire         phystatus1,         //                   .phystatus1
		input  wire         phystatus2,         //                   .phystatus2
		input  wire         phystatus3,         //                   .phystatus3
		input  wire [7:0]   rxdata0,            //                   .rxdata0
		input  wire [7:0]   rxdata1,            //                   .rxdata1
		input  wire [7:0]   rxdata2,            //                   .rxdata2
		input  wire [7:0]   rxdata3,            //                   .rxdata3
		input  wire         rxdatak0,           //                   .rxdatak0
		input  wire         rxdatak1,           //                   .rxdatak1
		input  wire         rxdatak2,           //                   .rxdatak2
		input  wire         rxdatak3,           //                   .rxdatak3
		input  wire         rxelecidle0,        //                   .rxelecidle0
		input  wire         rxelecidle1,        //                   .rxelecidle1
		input  wire         rxelecidle2,        //                   .rxelecidle2
		input  wire         rxelecidle3,        //                   .rxelecidle3
		input  wire [2:0]   rxstatus0,          //                   .rxstatus0
		input  wire [2:0]   rxstatus1,          //                   .rxstatus1
		input  wire [2:0]   rxstatus2,          //                   .rxstatus2
		input  wire [2:0]   rxstatus3,          //                   .rxstatus3
		input  wire         rxvalid0,           //                   .rxvalid0
		input  wire         rxvalid1,           //                   .rxvalid1
		input  wire         rxvalid2,           //                   .rxvalid2
		input  wire         rxvalid3,           //                   .rxvalid3
		output wire         reset_status,       //            hip_rst.reset_status
		output wire         serdes_pll_locked,  //                   .serdes_pll_locked
		output wire         pld_clk_inuse,      //                   .pld_clk_inuse
		input  wire         pld_core_ready,     //                   .pld_core_ready
		output wire         testin_zero,        //                   .testin_zero
		input  wire [11:0]  lmi_addr,           //                lmi.lmi_addr
		input  wire [31:0]  lmi_din,            //                   .lmi_din
		input  wire         lmi_rden,           //                   .lmi_rden
		input  wire         lmi_wren,           //                   .lmi_wren
		output wire         lmi_ack,            //                   .lmi_ack
		output wire [31:0]  lmi_dout,           //                   .lmi_dout
		input  wire         pm_auxpwr,          //         power_mngt.pm_auxpwr
		input  wire [9:0]   pm_data,            //                   .pm_data
		input  wire         pme_to_cr,          //                   .pme_to_cr
		input  wire         pm_event,           //                   .pm_event
		output wire         pme_to_sr,          //                   .pme_to_sr
		input  wire [349:0] reconfig_to_xcvr,   //   reconfig_to_xcvr.reconfig_to_xcvr
		output wire [229:0] reconfig_from_xcvr, // reconfig_from_xcvr.reconfig_from_xcvr
		input  wire [4:0]   app_msi_num,        //            int_msi.app_msi_num
		input  wire         app_msi_req,        //                   .app_msi_req
		input  wire [2:0]   app_msi_tc,         //                   .app_msi_tc
		output wire         app_msi_ack,        //                   .app_msi_ack
		input  wire         app_int_sts_vec,    //                   .app_int_sts
		input  wire [4:0]   tl_hpg_ctrl_er,     //          config_tl.hpg_ctrler
		output wire [31:0]  tl_cfg_ctl,         //                   .tl_cfg_ctl
		input  wire [6:0]   cpl_err,            //                   .cpl_err
		output wire [3:0]   tl_cfg_add,         //                   .tl_cfg_add
		output wire         tl_cfg_ctl_wr,      //                   .tl_cfg_ctl_wr
		output wire         tl_cfg_sts_wr,      //                   .tl_cfg_sts_wr
		output wire [52:0]  tl_cfg_sts,         //                   .tl_cfg_sts
		input  wire [0:0]   cpl_pending,        //                   .cpl_pending
		output wire         derr_cor_ext_rcv0,  //         hip_status.derr_cor_ext_rcv
		output wire         derr_cor_ext_rpl,   //                   .derr_cor_ext_rpl
		output wire         derr_rpl,           //                   .derr_rpl
		output wire         dlup_exit,          //                   .dlup_exit
		output wire [4:0]   dl_ltssm,           //                   .ltssmstate
		output wire         ev128ns,            //                   .ev128ns
		output wire         ev1us,              //                   .ev1us
		output wire         hotrst_exit,        //                   .hotrst_exit
		output wire [3:0]   int_status,         //                   .int_status
		output wire         l2_exit,            //                   .l2_exit
		output wire [3:0]   lane_act,           //                   .lane_act
		output wire [7:0]   ko_cpl_spc_header,  //                   .ko_cpl_spc_header
		output wire [11:0]  ko_cpl_spc_data,    //                   .ko_cpl_spc_data
		output wire [1:0]   dl_current_speed    //   hip_currentspeed.currentspeed
	);

	altera_pcie_cv_hip_ast_0001 #(
		.ACDS_VERSION_HWTCL                        ("18.1"),
		.lane_mask_hwtcl                           ("x4"),
		.gen12_lane_rate_mode_hwtcl                ("Gen1 (2.5 Gbps)"),
		.pcie_spec_version_hwtcl                   ("2.1"),
		.ast_width_hwtcl                           ("Avalon-ST 64-bit"),
		.pll_refclk_freq_hwtcl                     ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl               (0),
		.in_cvp_mode_hwtcl                         (0),
		.hip_reconfig_hwtcl                        (0),
		.num_of_func_hwtcl                         (1),
		.use_crc_forwarding_hwtcl                  (0),
		.port_link_number_hwtcl                    (1),
		.slotclkcfg_hwtcl                          (1),
		.enable_slot_register_hwtcl                (0),
		.vsec_id_hwtcl                             (4466),
		.vsec_rev_hwtcl                            (0),
		.user_id_hwtcl                             (0),
		.porttype_func0_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_0_hwtcl                    (16),
		.bar0_io_space_0_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_0_hwtcl              ("Enabled"),
		.bar0_prefetchable_0_hwtcl                 ("Enabled"),
		.bar1_size_mask_0_hwtcl                    (0),
		.bar1_io_space_0_hwtcl                     ("Disabled"),
		.bar1_prefetchable_0_hwtcl                 ("Disabled"),
		.bar2_size_mask_0_hwtcl                    (0),
		.bar2_io_space_0_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_0_hwtcl              ("Disabled"),
		.bar2_prefetchable_0_hwtcl                 ("Disabled"),
		.bar3_size_mask_0_hwtcl                    (0),
		.bar3_io_space_0_hwtcl                     ("Disabled"),
		.bar3_prefetchable_0_hwtcl                 ("Disabled"),
		.bar4_size_mask_0_hwtcl                    (16),
		.bar4_io_space_0_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_0_hwtcl              ("Enabled"),
		.bar4_prefetchable_0_hwtcl                 ("Enabled"),
		.bar5_size_mask_0_hwtcl                    (0),
		.bar5_io_space_0_hwtcl                     ("Disabled"),
		.bar5_prefetchable_0_hwtcl                 ("Disabled"),
		.expansion_base_address_register_0_hwtcl   (0),
		.io_window_addr_width_hwtcl                (0),
		.prefetchable_mem_window_addr_width_hwtcl  (0),
		.vendor_id_0_hwtcl                         (4466),
		.device_id_0_hwtcl                         (57347),
		.revision_id_0_hwtcl                       (1),
		.class_code_0_hwtcl                        (0),
		.subsystem_vendor_id_0_hwtcl               (0),
		.subsystem_device_id_0_hwtcl               (10337),
		.max_payload_size_0_hwtcl                  (256),
		.extend_tag_field_0_hwtcl                  ("32"),
		.completion_timeout_0_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_0_hwtcl (1),
		.flr_capability_0_hwtcl                    (0),
		.use_aer_0_hwtcl                           (0),
		.ecrc_check_capable_0_hwtcl                (0),
		.ecrc_gen_capable_0_hwtcl                  (0),
		.dll_active_report_support_0_hwtcl         (0),
		.surprise_down_error_support_0_hwtcl       (0),
		.msi_multi_message_capable_0_hwtcl         ("1"),
		.msi_64bit_addressing_capable_0_hwtcl      ("true"),
		.msi_masking_capable_0_hwtcl               ("false"),
		.msi_support_0_hwtcl                       ("true"),
		.enable_function_msix_support_0_hwtcl      (0),
		.msix_table_size_0_hwtcl                   (0),
		.msix_table_offset_0_hwtcl                 ("0"),
		.msix_table_bir_0_hwtcl                    (0),
		.msix_pba_offset_0_hwtcl                   ("0"),
		.msix_pba_bir_0_hwtcl                      (0),
		.interrupt_pin_0_hwtcl                     ("inta"),
		.slot_power_scale_0_hwtcl                  (0),
		.slot_power_limit_0_hwtcl                  (0),
		.slot_number_0_hwtcl                       (0),
		.rx_ei_l0s_0_hwtcl                         (0),
		.endpoint_l0_latency_0_hwtcl               (0),
		.endpoint_l1_latency_0_hwtcl               (0),
		.reconfig_to_xcvr_width                    (350),
		.hip_hard_reset_hwtcl                      (1),
		.reconfig_from_xcvr_width                  (230),
		.single_rx_detect_hwtcl                    (4),
		.enable_l0s_aspm_hwtcl                     ("false"),
		.aspm_optionality_hwtcl                    ("true"),
		.enable_adapter_half_rate_mode_hwtcl       ("false"),
		.millisecond_cycle_count_hwtcl             (124250),
		.credit_buffer_allocation_aux_hwtcl        ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl      (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl        (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl   (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl     (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl       (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl         (0),
		.cpl_spc_header_hwtcl                      (67),
		.cpl_spc_data_hwtcl                        (269),
		.port_width_data_hwtcl                     (64),
		.bypass_clk_switch_hwtcl                   ("disable"),
		.cvp_rate_sel_hwtcl                        ("full_rate"),
		.cvp_data_compressed_hwtcl                 ("false"),
		.cvp_data_encrypted_hwtcl                  ("false"),
		.cvp_mode_reset_hwtcl                      ("false"),
		.cvp_clk_reset_hwtcl                       ("false"),
		.core_clk_sel_hwtcl                        ("pld_clk"),
		.enable_rx_buffer_checking_hwtcl           ("false"),
		.disable_link_x2_support_hwtcl             ("false"),
		.device_number_hwtcl                       (0),
		.pipex1_debug_sel_hwtcl                    ("disable"),
		.pclk_out_sel_hwtcl                        ("pclk"),
		.no_soft_reset_hwtcl                       ("false"),
		.d1_support_hwtcl                          ("false"),
		.d2_support_hwtcl                          ("false"),
		.d0_pme_hwtcl                              ("false"),
		.d1_pme_hwtcl                              ("false"),
		.d2_pme_hwtcl                              ("false"),
		.d3_hot_pme_hwtcl                          ("false"),
		.d3_cold_pme_hwtcl                         ("false"),
		.low_priority_vc_hwtcl                     ("single_vc"),
		.enable_l1_aspm_hwtcl                      ("false"),
		.l1_exit_latency_sameclock_hwtcl           (0),
		.l1_exit_latency_diffclock_hwtcl           (0),
		.hot_plug_support_hwtcl                    (0),
		.no_command_completed_hwtcl                ("false"),
		.eie_before_nfts_count_hwtcl               (4),
		.gen2_diffclock_nfts_count_hwtcl           (255),
		.gen2_sameclock_nfts_count_hwtcl           (255),
		.deemphasis_enable_hwtcl                   ("false"),
		.l0_exit_latency_sameclock_hwtcl           (6),
		.l0_exit_latency_diffclock_hwtcl           (6),
		.vc0_clk_enable_hwtcl                      ("true"),
		.register_pipe_signals_hwtcl               ("true"),
		.tx_cdc_almost_empty_hwtcl                 (5),
		.rx_l0s_count_idl_hwtcl                    (0),
		.cdc_dummy_insert_limit_hwtcl              (11),
		.ei_delay_powerdown_count_hwtcl            (10),
		.skp_os_schedule_count_hwtcl               (0),
		.fc_init_timer_hwtcl                       (1024),
		.l01_entry_latency_hwtcl                   (31),
		.flow_control_update_count_hwtcl           (30),
		.flow_control_timeout_count_hwtcl          (200),
		.retry_buffer_last_active_address_hwtcl    (255),
		.reserved_debug_hwtcl                      (0),
		.use_tl_cfg_sync_hwtcl                     (1),
		.diffclock_nfts_count_hwtcl                (255),
		.sameclock_nfts_count_hwtcl                (255),
		.l2_async_logic_hwtcl                      ("disable"),
		.rx_cdc_almost_full_hwtcl                  (12),
		.tx_cdc_almost_full_hwtcl                  (11),
		.indicator_hwtcl                           (0),
		.maximum_current_0_hwtcl                   (0),
		.disable_snoop_packet_0_hwtcl              ("false"),
		.bridge_port_vga_enable_0_hwtcl            ("false"),
		.bridge_port_ssid_support_0_hwtcl          ("false"),
		.ssvid_0_hwtcl                             (0),
		.ssid_0_hwtcl                              (0),
		.porttype_func1_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_1_hwtcl                    (28),
		.bar0_io_space_1_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_1_hwtcl              ("Enabled"),
		.bar0_prefetchable_1_hwtcl                 ("Enabled"),
		.bar1_size_mask_1_hwtcl                    (0),
		.bar1_io_space_1_hwtcl                     ("Disabled"),
		.bar1_prefetchable_1_hwtcl                 ("Disabled"),
		.bar2_size_mask_1_hwtcl                    (0),
		.bar2_io_space_1_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_1_hwtcl              ("Disabled"),
		.bar2_prefetchable_1_hwtcl                 ("Disabled"),
		.bar3_size_mask_1_hwtcl                    (0),
		.bar3_io_space_1_hwtcl                     ("Disabled"),
		.bar3_prefetchable_1_hwtcl                 ("Disabled"),
		.bar4_size_mask_1_hwtcl                    (0),
		.bar4_io_space_1_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_1_hwtcl              ("Disabled"),
		.bar4_prefetchable_1_hwtcl                 ("Disabled"),
		.bar5_size_mask_1_hwtcl                    (0),
		.bar5_io_space_1_hwtcl                     ("Disabled"),
		.bar5_prefetchable_1_hwtcl                 ("Disabled"),
		.expansion_base_address_register_1_hwtcl   (0),
		.vendor_id_1_hwtcl                         (0),
		.device_id_1_hwtcl                         (1),
		.revision_id_1_hwtcl                       (1),
		.class_code_1_hwtcl                        (0),
		.subsystem_vendor_id_1_hwtcl               (0),
		.subsystem_device_id_1_hwtcl               (0),
		.max_payload_size_1_hwtcl                  (256),
		.extend_tag_field_1_hwtcl                  ("32"),
		.completion_timeout_1_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_1_hwtcl (1),
		.flr_capability_1_hwtcl                    (0),
		.use_aer_1_hwtcl                           (0),
		.ecrc_check_capable_1_hwtcl                (0),
		.ecrc_gen_capable_1_hwtcl                  (0),
		.dll_active_report_support_1_hwtcl         (0),
		.surprise_down_error_support_1_hwtcl       (0),
		.msi_multi_message_capable_1_hwtcl         ("4"),
		.msi_64bit_addressing_capable_1_hwtcl      ("true"),
		.msi_masking_capable_1_hwtcl               ("false"),
		.msi_support_1_hwtcl                       ("true"),
		.enable_function_msix_support_1_hwtcl      (0),
		.msix_table_size_1_hwtcl                   (0),
		.msix_table_offset_1_hwtcl                 ("0"),
		.msix_table_bir_1_hwtcl                    (0),
		.msix_pba_offset_1_hwtcl                   ("0"),
		.msix_pba_bir_1_hwtcl                      (0),
		.interrupt_pin_1_hwtcl                     ("inta"),
		.slot_power_scale_1_hwtcl                  (0),
		.slot_power_limit_1_hwtcl                  (0),
		.slot_number_1_hwtcl                       (0),
		.rx_ei_l0s_1_hwtcl                         (0),
		.endpoint_l0_latency_1_hwtcl               (0),
		.endpoint_l1_latency_1_hwtcl               (0),
		.maximum_current_1_hwtcl                   (0),
		.disable_snoop_packet_1_hwtcl              ("false"),
		.bridge_port_vga_enable_1_hwtcl            ("false"),
		.bridge_port_ssid_support_1_hwtcl          ("false"),
		.ssvid_1_hwtcl                             (0),
		.ssid_1_hwtcl                              (0),
		.porttype_func2_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_2_hwtcl                    (28),
		.bar0_io_space_2_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_2_hwtcl              ("Enabled"),
		.bar0_prefetchable_2_hwtcl                 ("Enabled"),
		.bar1_size_mask_2_hwtcl                    (0),
		.bar1_io_space_2_hwtcl                     ("Disabled"),
		.bar1_prefetchable_2_hwtcl                 ("Disabled"),
		.bar2_size_mask_2_hwtcl                    (0),
		.bar2_io_space_2_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_2_hwtcl              ("Disabled"),
		.bar2_prefetchable_2_hwtcl                 ("Disabled"),
		.bar3_size_mask_2_hwtcl                    (0),
		.bar3_io_space_2_hwtcl                     ("Disabled"),
		.bar3_prefetchable_2_hwtcl                 ("Disabled"),
		.bar4_size_mask_2_hwtcl                    (0),
		.bar4_io_space_2_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_2_hwtcl              ("Disabled"),
		.bar4_prefetchable_2_hwtcl                 ("Disabled"),
		.bar5_size_mask_2_hwtcl                    (0),
		.bar5_io_space_2_hwtcl                     ("Disabled"),
		.bar5_prefetchable_2_hwtcl                 ("Disabled"),
		.expansion_base_address_register_2_hwtcl   (0),
		.vendor_id_2_hwtcl                         (0),
		.device_id_2_hwtcl                         (1),
		.revision_id_2_hwtcl                       (1),
		.class_code_2_hwtcl                        (0),
		.subsystem_vendor_id_2_hwtcl               (0),
		.subsystem_device_id_2_hwtcl               (0),
		.max_payload_size_2_hwtcl                  (256),
		.extend_tag_field_2_hwtcl                  ("32"),
		.completion_timeout_2_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_2_hwtcl (1),
		.flr_capability_2_hwtcl                    (0),
		.use_aer_2_hwtcl                           (0),
		.ecrc_check_capable_2_hwtcl                (0),
		.ecrc_gen_capable_2_hwtcl                  (0),
		.dll_active_report_support_2_hwtcl         (0),
		.surprise_down_error_support_2_hwtcl       (0),
		.msi_multi_message_capable_2_hwtcl         ("4"),
		.msi_64bit_addressing_capable_2_hwtcl      ("true"),
		.msi_masking_capable_2_hwtcl               ("false"),
		.msi_support_2_hwtcl                       ("true"),
		.enable_function_msix_support_2_hwtcl      (0),
		.msix_table_size_2_hwtcl                   (0),
		.msix_table_offset_2_hwtcl                 ("0"),
		.msix_table_bir_2_hwtcl                    (0),
		.msix_pba_offset_2_hwtcl                   ("0"),
		.msix_pba_bir_2_hwtcl                      (0),
		.interrupt_pin_2_hwtcl                     ("inta"),
		.slot_power_scale_2_hwtcl                  (0),
		.slot_power_limit_2_hwtcl                  (0),
		.slot_number_2_hwtcl                       (0),
		.rx_ei_l0s_2_hwtcl                         (0),
		.endpoint_l0_latency_2_hwtcl               (0),
		.endpoint_l1_latency_2_hwtcl               (0),
		.maximum_current_2_hwtcl                   (0),
		.disable_snoop_packet_2_hwtcl              ("false"),
		.bridge_port_vga_enable_2_hwtcl            ("false"),
		.bridge_port_ssid_support_2_hwtcl          ("false"),
		.ssvid_2_hwtcl                             (0),
		.ssid_2_hwtcl                              (0),
		.porttype_func3_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_3_hwtcl                    (28),
		.bar0_io_space_3_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_3_hwtcl              ("Enabled"),
		.bar0_prefetchable_3_hwtcl                 ("Enabled"),
		.bar1_size_mask_3_hwtcl                    (0),
		.bar1_io_space_3_hwtcl                     ("Disabled"),
		.bar1_prefetchable_3_hwtcl                 ("Disabled"),
		.bar2_size_mask_3_hwtcl                    (0),
		.bar2_io_space_3_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_3_hwtcl              ("Disabled"),
		.bar2_prefetchable_3_hwtcl                 ("Disabled"),
		.bar3_size_mask_3_hwtcl                    (0),
		.bar3_io_space_3_hwtcl                     ("Disabled"),
		.bar3_prefetchable_3_hwtcl                 ("Disabled"),
		.bar4_size_mask_3_hwtcl                    (0),
		.bar4_io_space_3_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_3_hwtcl              ("Disabled"),
		.bar4_prefetchable_3_hwtcl                 ("Disabled"),
		.bar5_size_mask_3_hwtcl                    (0),
		.bar5_io_space_3_hwtcl                     ("Disabled"),
		.bar5_prefetchable_3_hwtcl                 ("Disabled"),
		.expansion_base_address_register_3_hwtcl   (0),
		.vendor_id_3_hwtcl                         (0),
		.device_id_3_hwtcl                         (1),
		.revision_id_3_hwtcl                       (1),
		.class_code_3_hwtcl                        (0),
		.subsystem_vendor_id_3_hwtcl               (0),
		.subsystem_device_id_3_hwtcl               (0),
		.max_payload_size_3_hwtcl                  (256),
		.extend_tag_field_3_hwtcl                  ("32"),
		.completion_timeout_3_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_3_hwtcl (1),
		.flr_capability_3_hwtcl                    (0),
		.use_aer_3_hwtcl                           (0),
		.ecrc_check_capable_3_hwtcl                (0),
		.ecrc_gen_capable_3_hwtcl                  (0),
		.dll_active_report_support_3_hwtcl         (0),
		.surprise_down_error_support_3_hwtcl       (0),
		.msi_multi_message_capable_3_hwtcl         ("4"),
		.msi_64bit_addressing_capable_3_hwtcl      ("true"),
		.msi_masking_capable_3_hwtcl               ("false"),
		.msi_support_3_hwtcl                       ("true"),
		.enable_function_msix_support_3_hwtcl      (0),
		.msix_table_size_3_hwtcl                   (0),
		.msix_table_offset_3_hwtcl                 ("0"),
		.msix_table_bir_3_hwtcl                    (0),
		.msix_pba_offset_3_hwtcl                   ("0"),
		.msix_pba_bir_3_hwtcl                      (0),
		.interrupt_pin_3_hwtcl                     ("inta"),
		.slot_power_scale_3_hwtcl                  (0),
		.slot_power_limit_3_hwtcl                  (0),
		.slot_number_3_hwtcl                       (0),
		.rx_ei_l0s_3_hwtcl                         (0),
		.endpoint_l0_latency_3_hwtcl               (0),
		.endpoint_l1_latency_3_hwtcl               (0),
		.maximum_current_3_hwtcl                   (0),
		.disable_snoop_packet_3_hwtcl              ("false"),
		.bridge_port_vga_enable_3_hwtcl            ("false"),
		.bridge_port_ssid_support_3_hwtcl          ("false"),
		.ssvid_3_hwtcl                             (0),
		.ssid_3_hwtcl                              (0),
		.porttype_func4_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_4_hwtcl                    (28),
		.bar0_io_space_4_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_4_hwtcl              ("Enabled"),
		.bar0_prefetchable_4_hwtcl                 ("Enabled"),
		.bar1_size_mask_4_hwtcl                    (0),
		.bar1_io_space_4_hwtcl                     ("Disabled"),
		.bar1_prefetchable_4_hwtcl                 ("Disabled"),
		.bar2_size_mask_4_hwtcl                    (0),
		.bar2_io_space_4_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_4_hwtcl              ("Disabled"),
		.bar2_prefetchable_4_hwtcl                 ("Disabled"),
		.bar3_size_mask_4_hwtcl                    (0),
		.bar3_io_space_4_hwtcl                     ("Disabled"),
		.bar3_prefetchable_4_hwtcl                 ("Disabled"),
		.bar4_size_mask_4_hwtcl                    (0),
		.bar4_io_space_4_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_4_hwtcl              ("Disabled"),
		.bar4_prefetchable_4_hwtcl                 ("Disabled"),
		.bar5_size_mask_4_hwtcl                    (0),
		.bar5_io_space_4_hwtcl                     ("Disabled"),
		.bar5_prefetchable_4_hwtcl                 ("Disabled"),
		.expansion_base_address_register_4_hwtcl   (0),
		.vendor_id_4_hwtcl                         (0),
		.device_id_4_hwtcl                         (1),
		.revision_id_4_hwtcl                       (1),
		.class_code_4_hwtcl                        (0),
		.subsystem_vendor_id_4_hwtcl               (0),
		.subsystem_device_id_4_hwtcl               (0),
		.max_payload_size_4_hwtcl                  (256),
		.extend_tag_field_4_hwtcl                  ("32"),
		.completion_timeout_4_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_4_hwtcl (1),
		.flr_capability_4_hwtcl                    (0),
		.use_aer_4_hwtcl                           (0),
		.ecrc_check_capable_4_hwtcl                (0),
		.ecrc_gen_capable_4_hwtcl                  (0),
		.dll_active_report_support_4_hwtcl         (0),
		.surprise_down_error_support_4_hwtcl       (0),
		.msi_multi_message_capable_4_hwtcl         ("4"),
		.msi_64bit_addressing_capable_4_hwtcl      ("true"),
		.msi_masking_capable_4_hwtcl               ("false"),
		.msi_support_4_hwtcl                       ("true"),
		.enable_function_msix_support_4_hwtcl      (0),
		.msix_table_size_4_hwtcl                   (0),
		.msix_table_offset_4_hwtcl                 ("0"),
		.msix_table_bir_4_hwtcl                    (0),
		.msix_pba_offset_4_hwtcl                   ("0"),
		.msix_pba_bir_4_hwtcl                      (0),
		.interrupt_pin_4_hwtcl                     ("inta"),
		.slot_power_scale_4_hwtcl                  (0),
		.slot_power_limit_4_hwtcl                  (0),
		.slot_number_4_hwtcl                       (0),
		.rx_ei_l0s_4_hwtcl                         (0),
		.endpoint_l0_latency_4_hwtcl               (0),
		.endpoint_l1_latency_4_hwtcl               (0),
		.maximum_current_4_hwtcl                   (0),
		.disable_snoop_packet_4_hwtcl              ("false"),
		.bridge_port_vga_enable_4_hwtcl            ("false"),
		.bridge_port_ssid_support_4_hwtcl          ("false"),
		.ssvid_4_hwtcl                             (0),
		.ssid_4_hwtcl                              (0),
		.porttype_func5_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_5_hwtcl                    (28),
		.bar0_io_space_5_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_5_hwtcl              ("Enabled"),
		.bar0_prefetchable_5_hwtcl                 ("Enabled"),
		.bar1_size_mask_5_hwtcl                    (0),
		.bar1_io_space_5_hwtcl                     ("Disabled"),
		.bar1_prefetchable_5_hwtcl                 ("Disabled"),
		.bar2_size_mask_5_hwtcl                    (0),
		.bar2_io_space_5_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_5_hwtcl              ("Disabled"),
		.bar2_prefetchable_5_hwtcl                 ("Disabled"),
		.bar3_size_mask_5_hwtcl                    (0),
		.bar3_io_space_5_hwtcl                     ("Disabled"),
		.bar3_prefetchable_5_hwtcl                 ("Disabled"),
		.bar4_size_mask_5_hwtcl                    (0),
		.bar4_io_space_5_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_5_hwtcl              ("Disabled"),
		.bar4_prefetchable_5_hwtcl                 ("Disabled"),
		.bar5_size_mask_5_hwtcl                    (0),
		.bar5_io_space_5_hwtcl                     ("Disabled"),
		.bar5_prefetchable_5_hwtcl                 ("Disabled"),
		.expansion_base_address_register_5_hwtcl   (0),
		.vendor_id_5_hwtcl                         (0),
		.device_id_5_hwtcl                         (1),
		.revision_id_5_hwtcl                       (1),
		.class_code_5_hwtcl                        (0),
		.subsystem_vendor_id_5_hwtcl               (0),
		.subsystem_device_id_5_hwtcl               (0),
		.max_payload_size_5_hwtcl                  (256),
		.extend_tag_field_5_hwtcl                  ("32"),
		.completion_timeout_5_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_5_hwtcl (1),
		.flr_capability_5_hwtcl                    (0),
		.use_aer_5_hwtcl                           (0),
		.ecrc_check_capable_5_hwtcl                (0),
		.ecrc_gen_capable_5_hwtcl                  (0),
		.dll_active_report_support_5_hwtcl         (0),
		.surprise_down_error_support_5_hwtcl       (0),
		.msi_multi_message_capable_5_hwtcl         ("4"),
		.msi_64bit_addressing_capable_5_hwtcl      ("true"),
		.msi_masking_capable_5_hwtcl               ("false"),
		.msi_support_5_hwtcl                       ("true"),
		.enable_function_msix_support_5_hwtcl      (0),
		.msix_table_size_5_hwtcl                   (0),
		.msix_table_offset_5_hwtcl                 ("0"),
		.msix_table_bir_5_hwtcl                    (0),
		.msix_pba_offset_5_hwtcl                   ("0"),
		.msix_pba_bir_5_hwtcl                      (0),
		.interrupt_pin_5_hwtcl                     ("inta"),
		.slot_power_scale_5_hwtcl                  (0),
		.slot_power_limit_5_hwtcl                  (0),
		.slot_number_5_hwtcl                       (0),
		.rx_ei_l0s_5_hwtcl                         (0),
		.endpoint_l0_latency_5_hwtcl               (0),
		.endpoint_l1_latency_5_hwtcl               (0),
		.maximum_current_5_hwtcl                   (0),
		.disable_snoop_packet_5_hwtcl              ("false"),
		.bridge_port_vga_enable_5_hwtcl            ("false"),
		.bridge_port_ssid_support_5_hwtcl          ("false"),
		.ssvid_5_hwtcl                             (0),
		.ssid_5_hwtcl                              (0),
		.porttype_func6_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_6_hwtcl                    (28),
		.bar0_io_space_6_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_6_hwtcl              ("Enabled"),
		.bar0_prefetchable_6_hwtcl                 ("Enabled"),
		.bar1_size_mask_6_hwtcl                    (0),
		.bar1_io_space_6_hwtcl                     ("Disabled"),
		.bar1_prefetchable_6_hwtcl                 ("Disabled"),
		.bar2_size_mask_6_hwtcl                    (0),
		.bar2_io_space_6_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_6_hwtcl              ("Disabled"),
		.bar2_prefetchable_6_hwtcl                 ("Disabled"),
		.bar3_size_mask_6_hwtcl                    (0),
		.bar3_io_space_6_hwtcl                     ("Disabled"),
		.bar3_prefetchable_6_hwtcl                 ("Disabled"),
		.bar4_size_mask_6_hwtcl                    (0),
		.bar4_io_space_6_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_6_hwtcl              ("Disabled"),
		.bar4_prefetchable_6_hwtcl                 ("Disabled"),
		.bar5_size_mask_6_hwtcl                    (0),
		.bar5_io_space_6_hwtcl                     ("Disabled"),
		.bar5_prefetchable_6_hwtcl                 ("Disabled"),
		.expansion_base_address_register_6_hwtcl   (0),
		.vendor_id_6_hwtcl                         (0),
		.device_id_6_hwtcl                         (1),
		.revision_id_6_hwtcl                       (1),
		.class_code_6_hwtcl                        (0),
		.subsystem_vendor_id_6_hwtcl               (0),
		.subsystem_device_id_6_hwtcl               (0),
		.max_payload_size_6_hwtcl                  (256),
		.extend_tag_field_6_hwtcl                  ("32"),
		.completion_timeout_6_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_6_hwtcl (1),
		.flr_capability_6_hwtcl                    (0),
		.use_aer_6_hwtcl                           (0),
		.ecrc_check_capable_6_hwtcl                (0),
		.ecrc_gen_capable_6_hwtcl                  (0),
		.dll_active_report_support_6_hwtcl         (0),
		.surprise_down_error_support_6_hwtcl       (0),
		.msi_multi_message_capable_6_hwtcl         ("4"),
		.msi_64bit_addressing_capable_6_hwtcl      ("true"),
		.msi_masking_capable_6_hwtcl               ("false"),
		.msi_support_6_hwtcl                       ("true"),
		.enable_function_msix_support_6_hwtcl      (0),
		.msix_table_size_6_hwtcl                   (0),
		.msix_table_offset_6_hwtcl                 ("0"),
		.msix_table_bir_6_hwtcl                    (0),
		.msix_pba_offset_6_hwtcl                   ("0"),
		.msix_pba_bir_6_hwtcl                      (0),
		.interrupt_pin_6_hwtcl                     ("inta"),
		.slot_power_scale_6_hwtcl                  (0),
		.slot_power_limit_6_hwtcl                  (0),
		.slot_number_6_hwtcl                       (0),
		.rx_ei_l0s_6_hwtcl                         (0),
		.endpoint_l0_latency_6_hwtcl               (0),
		.endpoint_l1_latency_6_hwtcl               (0),
		.maximum_current_6_hwtcl                   (0),
		.disable_snoop_packet_6_hwtcl              ("false"),
		.bridge_port_vga_enable_6_hwtcl            ("false"),
		.bridge_port_ssid_support_6_hwtcl          ("false"),
		.ssvid_6_hwtcl                             (0),
		.ssid_6_hwtcl                              (0),
		.porttype_func7_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_7_hwtcl                    (28),
		.bar0_io_space_7_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_7_hwtcl              ("Enabled"),
		.bar0_prefetchable_7_hwtcl                 ("Enabled"),
		.bar1_size_mask_7_hwtcl                    (0),
		.bar1_io_space_7_hwtcl                     ("Disabled"),
		.bar1_prefetchable_7_hwtcl                 ("Disabled"),
		.bar2_size_mask_7_hwtcl                    (0),
		.bar2_io_space_7_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_7_hwtcl              ("Disabled"),
		.bar2_prefetchable_7_hwtcl                 ("Disabled"),
		.bar3_size_mask_7_hwtcl                    (0),
		.bar3_io_space_7_hwtcl                     ("Disabled"),
		.bar3_prefetchable_7_hwtcl                 ("Disabled"),
		.bar4_size_mask_7_hwtcl                    (0),
		.bar4_io_space_7_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_7_hwtcl              ("Disabled"),
		.bar4_prefetchable_7_hwtcl                 ("Disabled"),
		.bar5_size_mask_7_hwtcl                    (0),
		.bar5_io_space_7_hwtcl                     ("Disabled"),
		.bar5_prefetchable_7_hwtcl                 ("Disabled"),
		.expansion_base_address_register_7_hwtcl   (0),
		.vendor_id_7_hwtcl                         (0),
		.device_id_7_hwtcl                         (1),
		.revision_id_7_hwtcl                       (1),
		.class_code_7_hwtcl                        (0),
		.subsystem_vendor_id_7_hwtcl               (0),
		.subsystem_device_id_7_hwtcl               (0),
		.max_payload_size_7_hwtcl                  (256),
		.extend_tag_field_7_hwtcl                  ("32"),
		.completion_timeout_7_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_7_hwtcl (1),
		.flr_capability_7_hwtcl                    (0),
		.use_aer_7_hwtcl                           (0),
		.ecrc_check_capable_7_hwtcl                (0),
		.ecrc_gen_capable_7_hwtcl                  (0),
		.dll_active_report_support_7_hwtcl         (0),
		.surprise_down_error_support_7_hwtcl       (0),
		.msi_multi_message_capable_7_hwtcl         ("4"),
		.msi_64bit_addressing_capable_7_hwtcl      ("true"),
		.msi_masking_capable_7_hwtcl               ("false"),
		.msi_support_7_hwtcl                       ("true"),
		.enable_function_msix_support_7_hwtcl      (0),
		.msix_table_size_7_hwtcl                   (0),
		.msix_table_offset_7_hwtcl                 ("0"),
		.msix_table_bir_7_hwtcl                    (0),
		.msix_pba_offset_7_hwtcl                   ("0"),
		.msix_pba_bir_7_hwtcl                      (0),
		.interrupt_pin_7_hwtcl                     ("inta"),
		.slot_power_scale_7_hwtcl                  (0),
		.slot_power_limit_7_hwtcl                  (0),
		.slot_number_7_hwtcl                       (0),
		.rx_ei_l0s_7_hwtcl                         (0),
		.endpoint_l0_latency_7_hwtcl               (0),
		.endpoint_l1_latency_7_hwtcl               (0),
		.maximum_current_7_hwtcl                   (0),
		.disable_snoop_packet_7_hwtcl              ("false"),
		.bridge_port_vga_enable_7_hwtcl            ("false"),
		.bridge_port_ssid_support_7_hwtcl          ("false"),
		.ssvid_7_hwtcl                             (0),
		.ssid_7_hwtcl                              (0),
		.rpre_emph_a_val_hwtcl                     (11),
		.rpre_emph_b_val_hwtcl                     (0),
		.rpre_emph_c_val_hwtcl                     (22),
		.rpre_emph_d_val_hwtcl                     (12),
		.rpre_emph_e_val_hwtcl                     (21),
		.rvod_sel_a_val_hwtcl                      (50),
		.rvod_sel_b_val_hwtcl                      (34),
		.rvod_sel_c_val_hwtcl                      (50),
		.rvod_sel_d_val_hwtcl                      (50),
		.rvod_sel_e_val_hwtcl                      (9)
	) pcie_inst (
		.npor                   (npor),                 //               npor.npor
		.pin_perst              (pin_perst),            //                   .pin_perst
		.test_in                (test_in),              //           hip_ctrl.test_in
		.simu_mode_pipe         (simu_mode_pipe),       //                   .simu_mode_pipe
		.pld_clk                (pld_clk),              //            pld_clk.clk
		.coreclkout             (coreclkout),           //     coreclkout_hip.clk
		.refclk                 (refclk),               //             refclk.clk
		.rx_in0                 (rx_in0),               //         hip_serial.rx_in0
		.rx_in1                 (rx_in1),               //                   .rx_in1
		.rx_in2                 (rx_in2),               //                   .rx_in2
		.rx_in3                 (rx_in3),               //                   .rx_in3
		.tx_out0                (tx_out0),              //                   .tx_out0
		.tx_out1                (tx_out1),              //                   .tx_out1
		.tx_out2                (tx_out2),              //                   .tx_out2
		.tx_out3                (tx_out3),              //                   .tx_out3
		.rx_st_valid            (rx_st_valid),          //              rx_st.valid
		.rx_st_sop              (rx_st_sop),            //                   .startofpacket
		.rx_st_eop              (rx_st_eop),            //                   .endofpacket
		.rx_st_ready            (rx_st_ready),          //                   .ready
		.rx_st_err              (rx_st_err),            //                   .error
		.rx_st_data             (rx_st_data),           //                   .data
		.rx_st_bar              (rx_st_bar),            //          rx_bar_be.rx_st_bar
		.rx_st_mask             (rx_st_mask),           //                   .rx_st_mask
		.tx_st_valid            (tx_st_valid),          //              tx_st.valid
		.tx_st_sop              (tx_st_sop),            //                   .startofpacket
		.tx_st_eop              (tx_st_eop),            //                   .endofpacket
		.tx_st_ready            (tx_st_ready),          //                   .ready
		.tx_st_err              (tx_st_err),            //                   .error
		.tx_st_data             (tx_st_data),           //                   .data
		.tx_fifo_empty          (tx_fifo_empty),        //            tx_fifo.fifo_empty
		.tx_cred_datafccp       (tx_cred_datafccp),     //            tx_cred.tx_cred_datafccp
		.tx_cred_datafcnp       (tx_cred_datafcnp),     //                   .tx_cred_datafcnp
		.tx_cred_datafcp        (tx_cred_datafcp),      //                   .tx_cred_datafcp
		.tx_cred_fchipcons      (tx_cred_fchipcons),    //                   .tx_cred_fchipcons
		.tx_cred_fcinfinite     (tx_cred_fcinfinite),   //                   .tx_cred_fcinfinite
		.tx_cred_hdrfccp        (tx_cred_hdrfccp),      //                   .tx_cred_hdrfccp
		.tx_cred_hdrfcnp        (tx_cred_hdrfcnp),      //                   .tx_cred_hdrfcnp
		.tx_cred_hdrfcp         (tx_cred_hdrfcp),       //                   .tx_cred_hdrfcp
		.sim_pipe_pclk_in       (sim_pipe_pclk_in),     //           hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate          (sim_pipe_rate),        //                   .sim_pipe_rate
		.sim_ltssmstate         (sim_ltssmstate),       //                   .sim_ltssmstate
		.eidleinfersel0         (eidleinfersel0),       //                   .eidleinfersel0
		.eidleinfersel1         (eidleinfersel1),       //                   .eidleinfersel1
		.eidleinfersel2         (eidleinfersel2),       //                   .eidleinfersel2
		.eidleinfersel3         (eidleinfersel3),       //                   .eidleinfersel3
		.powerdown0             (powerdown0),           //                   .powerdown0
		.powerdown1             (powerdown1),           //                   .powerdown1
		.powerdown2             (powerdown2),           //                   .powerdown2
		.powerdown3             (powerdown3),           //                   .powerdown3
		.rxpolarity0            (rxpolarity0),          //                   .rxpolarity0
		.rxpolarity1            (rxpolarity1),          //                   .rxpolarity1
		.rxpolarity2            (rxpolarity2),          //                   .rxpolarity2
		.rxpolarity3            (rxpolarity3),          //                   .rxpolarity3
		.txcompl0               (txcompl0),             //                   .txcompl0
		.txcompl1               (txcompl1),             //                   .txcompl1
		.txcompl2               (txcompl2),             //                   .txcompl2
		.txcompl3               (txcompl3),             //                   .txcompl3
		.txdata0                (txdata0),              //                   .txdata0
		.txdata1                (txdata1),              //                   .txdata1
		.txdata2                (txdata2),              //                   .txdata2
		.txdata3                (txdata3),              //                   .txdata3
		.txdatak0               (txdatak0),             //                   .txdatak0
		.txdatak1               (txdatak1),             //                   .txdatak1
		.txdatak2               (txdatak2),             //                   .txdatak2
		.txdatak3               (txdatak3),             //                   .txdatak3
		.txdetectrx0            (txdetectrx0),          //                   .txdetectrx0
		.txdetectrx1            (txdetectrx1),          //                   .txdetectrx1
		.txdetectrx2            (txdetectrx2),          //                   .txdetectrx2
		.txdetectrx3            (txdetectrx3),          //                   .txdetectrx3
		.txelecidle0            (txelecidle0),          //                   .txelecidle0
		.txelecidle1            (txelecidle1),          //                   .txelecidle1
		.txelecidle2            (txelecidle2),          //                   .txelecidle2
		.txelecidle3            (txelecidle3),          //                   .txelecidle3
		.txswing0               (txswing0),             //                   .txswing0
		.txswing1               (txswing1),             //                   .txswing1
		.txswing2               (txswing2),             //                   .txswing2
		.txswing3               (txswing3),             //                   .txswing3
		.txmargin0              (txmargin0),            //                   .txmargin0
		.txmargin1              (txmargin1),            //                   .txmargin1
		.txmargin2              (txmargin2),            //                   .txmargin2
		.txmargin3              (txmargin3),            //                   .txmargin3
		.txdeemph0              (txdeemph0),            //                   .txdeemph0
		.txdeemph1              (txdeemph1),            //                   .txdeemph1
		.txdeemph2              (txdeemph2),            //                   .txdeemph2
		.txdeemph3              (txdeemph3),            //                   .txdeemph3
		.phystatus0             (phystatus0),           //                   .phystatus0
		.phystatus1             (phystatus1),           //                   .phystatus1
		.phystatus2             (phystatus2),           //                   .phystatus2
		.phystatus3             (phystatus3),           //                   .phystatus3
		.rxdata0                (rxdata0),              //                   .rxdata0
		.rxdata1                (rxdata1),              //                   .rxdata1
		.rxdata2                (rxdata2),              //                   .rxdata2
		.rxdata3                (rxdata3),              //                   .rxdata3
		.rxdatak0               (rxdatak0),             //                   .rxdatak0
		.rxdatak1               (rxdatak1),             //                   .rxdatak1
		.rxdatak2               (rxdatak2),             //                   .rxdatak2
		.rxdatak3               (rxdatak3),             //                   .rxdatak3
		.rxelecidle0            (rxelecidle0),          //                   .rxelecidle0
		.rxelecidle1            (rxelecidle1),          //                   .rxelecidle1
		.rxelecidle2            (rxelecidle2),          //                   .rxelecidle2
		.rxelecidle3            (rxelecidle3),          //                   .rxelecidle3
		.rxstatus0              (rxstatus0),            //                   .rxstatus0
		.rxstatus1              (rxstatus1),            //                   .rxstatus1
		.rxstatus2              (rxstatus2),            //                   .rxstatus2
		.rxstatus3              (rxstatus3),            //                   .rxstatus3
		.rxvalid0               (rxvalid0),             //                   .rxvalid0
		.rxvalid1               (rxvalid1),             //                   .rxvalid1
		.rxvalid2               (rxvalid2),             //                   .rxvalid2
		.rxvalid3               (rxvalid3),             //                   .rxvalid3
		.reset_status           (reset_status),         //            hip_rst.reset_status
		.serdes_pll_locked      (serdes_pll_locked),    //                   .serdes_pll_locked
		.pld_clk_inuse          (pld_clk_inuse),        //                   .pld_clk_inuse
		.pld_core_ready         (pld_core_ready),       //                   .pld_core_ready
		.testin_zero            (testin_zero),          //                   .testin_zero
		.lmi_addr               (lmi_addr),             //                lmi.lmi_addr
		.lmi_din                (lmi_din),              //                   .lmi_din
		.lmi_rden               (lmi_rden),             //                   .lmi_rden
		.lmi_wren               (lmi_wren),             //                   .lmi_wren
		.lmi_ack                (lmi_ack),              //                   .lmi_ack
		.lmi_dout               (lmi_dout),             //                   .lmi_dout
		.pm_auxpwr              (pm_auxpwr),            //         power_mngt.pm_auxpwr
		.pm_data                (pm_data),              //                   .pm_data
		.pme_to_cr              (pme_to_cr),            //                   .pme_to_cr
		.pm_event               (pm_event),             //                   .pm_event
		.pme_to_sr              (pme_to_sr),            //                   .pme_to_sr
		.reconfig_to_xcvr       (reconfig_to_xcvr),     //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr     (reconfig_from_xcvr),   // reconfig_from_xcvr.reconfig_from_xcvr
		.app_msi_num            (app_msi_num),          //            int_msi.app_msi_num
		.app_msi_req            (app_msi_req),          //                   .app_msi_req
		.app_msi_tc             (app_msi_tc),           //                   .app_msi_tc
		.app_msi_ack            (app_msi_ack),          //                   .app_msi_ack
		.app_int_sts_vec        (app_int_sts_vec),      //                   .app_int_sts
		.tl_hpg_ctrl_er         (tl_hpg_ctrl_er),       //          config_tl.hpg_ctrler
		.tl_cfg_ctl             (tl_cfg_ctl),           //                   .tl_cfg_ctl
		.cpl_err                (cpl_err),              //                   .cpl_err
		.tl_cfg_add             (tl_cfg_add),           //                   .tl_cfg_add
		.tl_cfg_ctl_wr          (tl_cfg_ctl_wr),        //                   .tl_cfg_ctl_wr
		.tl_cfg_sts_wr          (tl_cfg_sts_wr),        //                   .tl_cfg_sts_wr
		.tl_cfg_sts             (tl_cfg_sts),           //                   .tl_cfg_sts
		.cpl_pending            (cpl_pending),          //                   .cpl_pending
		.derr_cor_ext_rcv0      (derr_cor_ext_rcv0),    //         hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl       (derr_cor_ext_rpl),     //                   .derr_cor_ext_rpl
		.derr_rpl               (derr_rpl),             //                   .derr_rpl
		.dlup_exit              (dlup_exit),            //                   .dlup_exit
		.dl_ltssm               (dl_ltssm),             //                   .ltssmstate
		.ev128ns                (ev128ns),              //                   .ev128ns
		.ev1us                  (ev1us),                //                   .ev1us
		.hotrst_exit            (hotrst_exit),          //                   .hotrst_exit
		.int_status             (int_status),           //                   .int_status
		.l2_exit                (l2_exit),              //                   .l2_exit
		.lane_act               (lane_act),             //                   .lane_act
		.ko_cpl_spc_header      (ko_cpl_spc_header),    //                   .ko_cpl_spc_header
		.ko_cpl_spc_data        (ko_cpl_spc_data),      //                   .ko_cpl_spc_data
		.dl_current_speed       (dl_current_speed),     //   hip_currentspeed.currentspeed
		.rx_in4                 (1'b0),                 //        (terminated)
		.rx_in5                 (1'b0),                 //        (terminated)
		.rx_in6                 (1'b0),                 //        (terminated)
		.rx_in7                 (1'b0),                 //        (terminated)
		.tx_out4                (),                     //        (terminated)
		.tx_out5                (),                     //        (terminated)
		.tx_out6                (),                     //        (terminated)
		.tx_out7                (),                     //        (terminated)
		.rx_st_empty            (),                     //        (terminated)
		.rx_fifo_empty          (),                     //        (terminated)
		.rx_fifo_full           (),                     //        (terminated)
		.rx_bar_dec_func_num    (),                     //        (terminated)
		.rx_st_be               (),                     //        (terminated)
		.tx_st_empty            (1'b0),                 //        (terminated)
		.tx_fifo_full           (),                     //        (terminated)
		.tx_fifo_rdp            (),                     //        (terminated)
		.tx_fifo_wrp            (),                     //        (terminated)
		.eidleinfersel4         (),                     //        (terminated)
		.eidleinfersel5         (),                     //        (terminated)
		.eidleinfersel6         (),                     //        (terminated)
		.eidleinfersel7         (),                     //        (terminated)
		.powerdown4             (),                     //        (terminated)
		.powerdown5             (),                     //        (terminated)
		.powerdown6             (),                     //        (terminated)
		.powerdown7             (),                     //        (terminated)
		.rxpolarity4            (),                     //        (terminated)
		.rxpolarity5            (),                     //        (terminated)
		.rxpolarity6            (),                     //        (terminated)
		.rxpolarity7            (),                     //        (terminated)
		.txcompl4               (),                     //        (terminated)
		.txcompl5               (),                     //        (terminated)
		.txcompl6               (),                     //        (terminated)
		.txcompl7               (),                     //        (terminated)
		.txdata4                (),                     //        (terminated)
		.txdata5                (),                     //        (terminated)
		.txdata6                (),                     //        (terminated)
		.txdata7                (),                     //        (terminated)
		.txdatak4               (),                     //        (terminated)
		.txdatak5               (),                     //        (terminated)
		.txdatak6               (),                     //        (terminated)
		.txdatak7               (),                     //        (terminated)
		.txdetectrx4            (),                     //        (terminated)
		.txdetectrx5            (),                     //        (terminated)
		.txdetectrx6            (),                     //        (terminated)
		.txdetectrx7            (),                     //        (terminated)
		.txelecidle4            (),                     //        (terminated)
		.txelecidle5            (),                     //        (terminated)
		.txelecidle6            (),                     //        (terminated)
		.txelecidle7            (),                     //        (terminated)
		.txswing4               (),                     //        (terminated)
		.txswing5               (),                     //        (terminated)
		.txswing6               (),                     //        (terminated)
		.txswing7               (),                     //        (terminated)
		.txmargin4              (),                     //        (terminated)
		.txmargin5              (),                     //        (terminated)
		.txmargin6              (),                     //        (terminated)
		.txmargin7              (),                     //        (terminated)
		.txdeemph4              (),                     //        (terminated)
		.txdeemph5              (),                     //        (terminated)
		.txdeemph6              (),                     //        (terminated)
		.txdeemph7              (),                     //        (terminated)
		.phystatus4             (1'b0),                 //        (terminated)
		.phystatus5             (1'b0),                 //        (terminated)
		.phystatus6             (1'b0),                 //        (terminated)
		.phystatus7             (1'b0),                 //        (terminated)
		.rxdata4                (8'b00000000),          //        (terminated)
		.rxdata5                (8'b00000000),          //        (terminated)
		.rxdata6                (8'b00000000),          //        (terminated)
		.rxdata7                (8'b00000000),          //        (terminated)
		.rxdatak4               (1'b0),                 //        (terminated)
		.rxdatak5               (1'b0),                 //        (terminated)
		.rxdatak6               (1'b0),                 //        (terminated)
		.rxdatak7               (1'b0),                 //        (terminated)
		.rxelecidle4            (1'b0),                 //        (terminated)
		.rxelecidle5            (1'b0),                 //        (terminated)
		.rxelecidle6            (1'b0),                 //        (terminated)
		.rxelecidle7            (1'b0),                 //        (terminated)
		.rxstatus4              (3'b000),               //        (terminated)
		.rxstatus5              (3'b000),               //        (terminated)
		.rxstatus6              (3'b000),               //        (terminated)
		.rxstatus7              (3'b000),               //        (terminated)
		.rxvalid4               (1'b0),                 //        (terminated)
		.rxvalid5               (1'b0),                 //        (terminated)
		.rxvalid6               (1'b0),                 //        (terminated)
		.rxvalid7               (1'b0),                 //        (terminated)
		.sim_pipe_pclk_out      (),                     //        (terminated)
		.pm_event_func          (3'b000),               //        (terminated)
		.hip_reconfig_clk       (1'b0),                 //        (terminated)
		.hip_reconfig_rst_n     (1'b0),                 //        (terminated)
		.hip_reconfig_address   (10'b0000000000),       //        (terminated)
		.hip_reconfig_byte_en   (2'b00),                //        (terminated)
		.hip_reconfig_read      (1'b0),                 //        (terminated)
		.hip_reconfig_readdata  (),                     //        (terminated)
		.hip_reconfig_write     (1'b0),                 //        (terminated)
		.hip_reconfig_writedata (16'b0000000000000000), //        (terminated)
		.ser_shift_load         (1'b0),                 //        (terminated)
		.interface_sel          (1'b0),                 //        (terminated)
		.app_msi_func           (3'b000),               //        (terminated)
		.serr_out               (),                     //        (terminated)
		.aer_msi_num            (5'b00000),             //        (terminated)
		.pex_msi_num            (5'b00000),             //        (terminated)
		.cpl_err_func           (3'b000)                //        (terminated)
	);

endmodule
