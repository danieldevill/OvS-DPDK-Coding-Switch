// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OGmMVnWTKxsTXx6Nudo4JY6g2WSogIxRYK598Cn7HFNpH+uJ3hgQdWhzktIYS0sQ
7/ORwThEPbHiWJTHMdAylJeuwgu8FSvc9VCQBxPUDnPbF8C9jztXuY7jmBGzxzyk
Hl75PzPos0z2wm+rreIlsq1fGkaflNdCNRihFFwkoCs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 123904)
BX8tdi5bsYSBY0s8IVE8Z7NIyakkKkZySK13Q+iOqKrK08nZ/ttrw9NXEg9nP9JT
aw44EhUSo3eLEjtwU2loT1S4uvfDTCoUNQg4b79FTk0sBKvuOs63wItGml6d+gl5
uUE2MqTFExWPBrWqtRaVWMZ/FURPZnc30iM07MGlX5OX9ZAE2m1ga3ppeqx5hYQu
J9EX2OxT2SgZJLFd83989MjQTjPHfcdkidBtnd4tBPd35Qk86/xHKDm/eQ/KQOGz
mWlz/VVZu34l4g470GOdVZOfnqMUR2KrptcDXOdZLqKdXu1MQm7VLiBrDtYu7ZtV
rugcMAHCOF5HGOsYiBBpIMqe8FyJWgjSC9KGxDNng3EAGhIdOzO7yPXW8u+jjhUw
mHJoEDUXQgLJCEfNNeDonK0TtNPsEO37cABTTbj0ULlibRgUiD7h6nuiYQjhX7oi
tbGlmk/+KCNm9B5w6wmIn/Qk9UuDxHJvFYjjIC0/mp7uknYUJ8eFyB7aDEtD3geo
Dd5VjpMSEd8vfkay2MUW0KY7v0+qlY9t8ZbU+tv4+BQncjiMW9pQi9fnRC5/reK5
ElnZTj0ZJsfxR4Dtwk22vnZx0u42HHjYdLJycSKJ0yb6E4nr7oqCJ6GW/zJ2B/Ze
Kxeopw1KyYC14MrbEQPszGn9qCXHFNLSgDBZ/oXtU46wthDWp2f5guoRMCuMMlbH
FbPCnSj3/vhBKmvPYrUIByoZhM70FY5ztfmsl5jTMXuyg7hHcT+N6Ra2lcr2k0Lu
34KCfY897S3b1saSiBWLGWzcrQMSSmJXxsu2m781bg/5+pBECN6goB84gn3iXSyp
s+Jm1v8LXK3qSET2dUHkIgsVOVBaeNh6BHhb3wKhIAopG/Na/spQwgmnury8hMLJ
wEQg/wtzzuQ2vmZFjYLQZs3IO4SkN/QByoc51mlZmXpe1S22CyESQpbntVSTJw6a
zqKOz1IInHg6ijslthQXVp/KHE4X4WXXM3jZ8M1yX10R1jz1eUhACKwMLM2wkB97
VQBLAWL54G99AKRJM5lf59F+HvVVTHfZeHLUEgkt8dNE8QSPVH60TARoo63wjREi
9BpgVW7Or+jb+aV0CYUYT1PMTznqYos9qw0sQpWAXqDoATiL9hOkdg3XBMgMoLYR
6Z1QZenr0U6M5JAJ3QbdmKWoFC6GksSVQVFZbveVE+lbVPgpdNsg/8sGEGt3gy7Y
CyKCkQ20DBajPljSOEc+pWB0SnxTWCaHqOpNmB+LYQ0Rjde6YfWkLtmEOHqXNoXX
M3cqnljzOpsJVG9C1vo71rGOQ48uGoGal0miwohsfYbS1K2SfO1eo89lr1cj2laT
WnbTUpfOwclqVeUdEUgqudRnHW/pFLwfnfWenGhlbkjq8zzMyNaFoBJJIRqszPNl
1X389rD0Rnmta4BNDlKcqM/OpLspEB8XvdT+PQLg2QmIixpsMZPJaL11b6gm8UkK
THPkP9irWYZT0SlXbm+vqWuNajNM+en2edD3zl5cfxVdGVhcFviKjHyQ7WBfh94n
OlAY/jab7HORgkcvTp41qnCfv9l7VVJ85va6vKhi87E3hmD2hyDD5vFk9qsJIIsX
494HwC85GjqWrRRvgENMSHkQqzPy+KSPc5MulDkh8GXIalkg9S9RaV4N7K/qPSU1
Ds3cCGWuwQ1fmMD3/pWx8Gu6xWwXRLNGzPH3OXjqxt+M99K7MciTiHKhYsb90Bf1
rHPM16rEtLC9y2nZFMBe3s9UUyUS3su+nFzgn2so8bEJlF9jpQuYRTe7nK4dEPM6
fKw1d9rTSIRlDMjCkywkmZBPNCHd1+daOeLqUmFQXjttNNRAVymGrKmFYYTJevRp
GaXGZ95RY6wwZ6U7Z4bQHHGGNPRhdYirZqI4BYpTGHODiJo3ScmG6vxbulfXjDD4
VSiq2QMZKy7IiTf9H9lQLDwnODOCsNNYbnCTwJcrCTM2QTRRLD40dAaaPdOvOxyM
W487mYGtDGhy0xkZCu1VrlDMKUJ9vmJGCdOYgbaxu5kqinV02G9PuEWI91AgYEDl
uGd5pidwFUi5iAH8csQwOitWuXC9wL9zcysiN2isgb7lMjjqMnQBF6Z7KOo+V3/r
69mLWvJWbXaHPSYIIa7yai7RGO20IOadBfvONDJXjiI8Oyyy0kYF4rRzEOefbA2X
8jiumcq7qjc74SnCSiOGlFk9lAphr974eucu9LPGwzQCIPTpESY+wqaqxK2oFXU2
ihmcsE9vaayDiCvuCmlcagk7vCg3ShbK8ccLhgGM4JJ6sPalMcgpTu4YMoMrd1N9
OdFGxfEv2B1nmrmpGP6Jhcj6ivDuPC5rF/P/37oqkkxajV/q9kLLCygHlFYFWHJq
Dd2+dHnxBhVcUEGGJjJPaUsk5PhN2Jvw7akUIiY5l6WbOVTb4ZhQxjtayxyHAefe
Jb6zsm7GcyEcjYC8WpSPfpDdBLhX6ZFbLWUBt5bDLX9VxYb0l6jURZ1+Zo0LXypl
GUVH10iFGRbaIwil2lwetyRGvfyKhsdMtBAE09lXrPp9PhEiAyueWchK1ksgMHyZ
qt3AQlATugqterGWdLDVpMLfSQNARRlVkfZBgw9vomnmKmmiCqg0EROlt3cFlYyD
hszfwyN0lv/sYeldMFOENX/+ermeOuKWRIVx6v2Bws+scm45ixVKgjkyziIZM/fs
kij75829pNwKlrN6TwEMwY/cRj1jwgz3oX8b1mVx5c1aLyKPHtynduSrM6f+pTw9
l7jLrN9k3y9H+qCKYpfMw+50no6TPWgPXjys7nwPytPM9n/mE6XIZjbYpusnCmFS
bdMQDdBwL+deyI/i8eB4QH7W1BcE1zyK9JeVriXe1KjtwgvVcPsXuuuHwbmr1TqP
cK6yWp0EBZbO2CaV83BQCVhD8htIT0kVuhAaHhJp8zNR93eJRnlPhOvm2UzgHuyc
st/5TKbu6zpmdmOg6PsdDfWzUcgfFJ1F0A1XoOYZHI6WjL9q3tr5ktR0TySogOg/
Bq164h8KEjfeTcFMivQaOWcCB8SPNwT5YcRb7DV8fW3tdKOQF8Lx3vhFRJzXKw/m
lj5hJmsuefVJfRFZHv5FXG+t3CBEYnp2huX1mwjitf+hzTSQJtVHuqA0xEhaenKh
54by4jsmyRul0BqIVpV07je1fiteivs6u2PTfbz7LDGiDKVYDM4vbh4vH5LPupqU
ZfdM5lej8gX1cDhgYZaQsZRVPWy5FxfjZkdKftA8f0jnpvH3FytTmsUmgyzy3akr
GPqG6HYNYnFJtHDA6Ru1jGDOexQkRYzgUcdpaPCy8havrSM8t2jYQXR9rcNBKtcu
ZhsleaEo/rmVF7AELDQN0+4sZWr6vQK+cgpmK/CwOr/uQ/2uO1FdqlH0VWN0GAjh
mpOzfnj1kKWoAefUqAdULia2mJm4ZhVD1PAJiivQFOfMl1Q2tc+flUDXsoD9xeMg
2XIaq4nvc5NtptAbpIc8MUUlrOvMw5aV1KDqDB22GPb+HJspR4z5tn5GV/G/rp1F
cHnFw+EtrSUIEfXy0PxSDStSpSFjqdSZfQ5v52duiZbvWYFhwQy758mM/EHyUTxQ
QvY0WTgrMVMtfl1CQ8ljWMADyDNvyLOYvg3PdlqzBmGNAH5RqDd1fT2+lK12VndP
RZFYuA+w8xPjmB6c+tng0EQ6oWDxGdg1IS4EMg+GEHAqu4N+IbO1z1W4UuSn/uiq
PLbIiFxyO2lM4BByae+7IIkDS0Swx/9MaQPQEGxElZ/6T8jQaQFkCx1DV7Io5CUo
WshkWk51f7+940K197yKm3OhFbonHlnc8q9yZ8YKniXO9I+B4sbQAAlChz5cMtij
ipEI2zt7fWpetRhP3++mEtJmzk3pPlGzjuwcsfqxVa6PkBkfpSLab23LF7RxlChB
vbbsS91JW7UAQu/WqQ2Y9aF7zW2un6ZwWhh4nqC7nCmmmZcTwt6kx9kdOl72QjAv
GNzQ9wQiWUjRmaJqVFHzIUyPPkel2AH5tqy7NhSBJWmLxHEYF8QsgvXf1WW85LkB
Df/Bv6LKbpodt4mhUgKwZkYCL9sgA5dgioxVU0BWz3XXkQw3VlVT3IoZYChD65ZE
X6AhzBPn+aOLHU4WNep8iHm2Cp0T5VroT+e6jHWebFnnU4U6pqPMJt61LWOu/dkv
cCMkirtxrN8znig3wtUp/YlBu4Q/XukqXl6c+CZko0oAfA/9FWHcYnFK+W6Hnqjg
dJzkfaElodYGtq96qHzDyGF+UMQqo+bBMVtaLvZ+ifGVhyUeAPb8KL1VBzpkP+Vq
s6of2qiicMFokP0p0OExh45qKecEGS1YRWJu8gg2YUgLSFq+F2xOy1nFqLXIX47a
iIZQFnhtZqswEgxyTzVVri02h9NBKI+iDxh2pCe93h/ol0fYpCpVK+DxnQVnVb1K
Oln06tV+QV/sJS/DgSIbRG1nz/3DH8C1xvtCItprrvCIvOLUACsK+4iNLX1nMXcm
f3OuqJd87L0rjyAdxYych6Rh0Xa7NaCz5sfEvX7wuMGDXiEshrAPQGk7wXv/nbJn
3H9vP1VESJro0xVyeMrsiLW9B0gZzFIhNiQfG2YLUZ8oPH/Nm0XyqJ0iTZuHMJNn
q+UxP4yOwWw9DE039UuAvzkXZpVoRObcAoEh20Bhm9n0tGA92/fGs+aoC3AzTAzG
5GjiO2ObyrnDko55TDFVTuubdLrOB0GbSFrPvf1ba3CIdIFDjuMKuCcYcSBXDKso
ev7N2mC7uRF4efKbWtQ7HAohq++CCICmF0OTa4RBS48xQsS5sONjNg5Oq1vHBQ3J
1OKrg2fsta63X4fm0ugIfNSeOzDMus5rtnrBAJrMnGyog9RRq6FhLiVSRhNHv0E7
BnLQ/kAzwUrEH7w5ukihLwVj2BkI/E2+By9PzJDi8ckgfOpBkpLlj/DmIdiJSPnz
z2m/pSvtgGOOQakolqX1MqO/11MLNgm7xo+5rAjcinqBmLIscwREYy3nk5GNVIJ4
uQjWKuy5olRlfQzK1dtdTqoQEwsvPVPXxxGEjA51kL8/0Uj0QeNuRqkxMjXeKdbq
Dg9hzFo1JJfSpQrEk4K+GT+f9HcW5y9u9hraIAEbifTsFpz5ZFG3VslyT0Yf+UqD
Wu4nbm8NZ5Qwe+L5JX98Bzlg97GOgrnYyGNDGycrTOlk1Dmqg7MYtLrRPmVmRpiE
ELN28b06oJFavK/Fu7VpG/FM34/05tdfk9bihWzxj7oR3RTNS8dxouQC79BqKTQK
wmSp++eAFPv8+bqDdXtM97TfEhvvjb6B2WCGDrCRISYndN/FaepK9FcW5USrFDgq
H7I2npCNVpuSoE8fjjnXAaTO+B/iSW/WshZPnSiYz2OnIz41sqEVzx8kP4hA789o
lZ0L9C6+PDIZ/qcGNsVUN4wOYLNjUA64LqRcYZvdYPIuMNJVL3DjsyeAK/KoZca+
dWlxQSVwPC0WO+WRBsVvmB/7ksW3RqIEwbhCJnUM88pot9KLDP2ZxVYOM2QrWiR9
D8o/tzK27BMFV4psp00vZRByzRbSWDhRortWprFh66yNsm8nlcbHyeWvp5y/id01
dNltp+3LAd+WV2G5LKdl3yJvsGLT3/Gcp7Rt01JR8u/qpry/KtI93jSnBPUjdlmS
t/ScfxJzJM+V4UJi8QSpPPzdKb7s1O5ocKvIbigX0Hsi5a1riJNF1YUEfW6FkEVx
Y5pMJpod1MbItOFXpPt/yzgAxPersby2jCC6eguCguGfr/VauPWFnAeJnAi6K9nU
BmKp+DkTL2Bi44GGHBMvNiBr4NWhA/u8aYkDuF984nnsamORhu4W18IvtdAVdF1I
/v7kAUbJa742GhdQN1SYGwIIEgmIODYixPq979Xv78roLuVw3S/ITURBPe2FGeOd
AZtLCMW3OGNBzX+VyHLdsxjYKPEVS6Ym6PQDgKvMugkDPBnD3ORcL45m4R2yOfk/
Xus8iK0MqkPa0IbAHtd+zJzcxg4xEEC5Vm0V/9EtvF+pMDft9Yproa8hIVCpcHUR
yxHGtBH+nhGEix5n9X+SWA5YWYVhP9o2gKNiRUWGZD74zC41BaKNWGDZGiYO2hp6
WrVeK8GEo9ZmtMk6HsVZUB8bOK60NLTbhVvdhVHEtvf5XKxNE7NNjbnUfLH7kekI
Qa/tC0Eyev3FbXMbHOY40Rd85PS/ndt/BZBDjs5zvE6Y6KaLlI1vGNf7ntGH6j1z
vRzDjzr4+WtuSEjfse5JED1M5CF/D2M4KTppJgHPhDVuRI4M/zerSEHhhZ3LulxZ
WKj1zMq1nD5MlmkDwB4ilh67CrN0WLUd2xxzHNmyJMfrAyNwDS39a0nD897G8BaG
bbC9+40xHY3pV5aWSLPBHnbiHUvH0N06YA1P/PkdPW1kmmZ8BrIcNQeHJz1UnAyw
kMV20hszn5BTbA1THt8J6whxVFs3r/xvEBGFiYlQsCT0Fhu3pzrL0eNXPvdwakFL
Z0ab1x00if924I+QQ6dNwRg1aw1af4dFTnirb437g08S7/OoQxwtngIVXVtxhysU
YdZXrwzG0ggzdI6L1iczzbK1ZjKwn7iMlLwSdoPn9hHoYEGSuB5e/JRLEYkjteLZ
7fMtsGIDpXPqbkmHKHGJh+fShm1JnLP9KFXjp4/7UDC/Ll8aLqPIgBeqUZcPRgZL
B9yZ3SIWxdlQFrwGPqLsdfIaryRJcqiRlL4I9scKCYrQQ50apFfsXF1fXpFQIaKm
0H4U10ZswjXq5RoplR9rV94J+DnN7UHVnPtCbGDNKTdu535+5FcJNZz+fSkUAPmK
xEdUFqZfT3caZH/wT2FPg984/p5/gBRSpDqOXRLyYkjlE4Crgkzr/V8L5A5kF8Dj
lAJTkOW9iH80YFzo9GuOkRjwJZzX+GpIu/YbtcKnZCypujzQfa8Rcc9+lxW/Hfu+
3DNZ12vAO6OQV59OBLh9Wq+1j6EOMPTPg2CTrHHZp6MPqSPvgQDhb7EcIZUBjLUL
Db4KfBj5mRBDoriCnmNNZeF20wpo+w9AYLn5LcuQFUlaQBHwbci8b2BLdpdu5t26
OoO3yWzK4yEVrkf0qptzxwU0EnZ+wF1h8ZXJglHNQkQzeKVLvrRh82Yd+IeNBR8C
6SsH+T3DqRIvHGoyq0IdZTK7RhL6wvRRraV4uNYedjryveEsfT8n0nZ0/iiZ+DsJ
hlIgeb2CfbfpV5twCfctTEBOqn8lLKAyYibMsaOUgHpY5vtkst54RYO4A//i8Ox/
M1OPD4kof55/Z4CeFHWOEVZ03lsmWHdbsEMZZ8kjSG47SVkhNx5mht0KenMnKEcd
8YskraXEA7hukcvLfQ6cQBz4QUxoWt80+mnrPg93g0r4404ZtNHBtdybwiu/Dxmp
UAf1M4TJT1ni8SMzw8KdK4izsn+EVE534L2PWsYNFdMxNBZNMevljSuRVd2CuGts
Royse8rCBgRdqV9/tttT+a3Lb1p5zTF1VCtuEq2FqjWeRwhfdjQg+Q8c7gfo4+Da
iHQpgb6VbQZgn+ejZVqzrIc8TscvCXRxWT3t6FzHNuuUWvZCPTYAqB8e4TE0GiyB
6zT7lqjxiF0PvkLq5ddIgxH49jRPKdXP5YOlTVBAqJrZD939820EJ/FVxNYhPdo6
QW5kLQgmhiSmDT7YqeZTFcnovTd1B2KTKF1zbcmeI6/vCJzJhXJc7Jhl67XEl7Mg
c6EeQ8ZelNXyZfsdLRta4nwYxsVVw68HnbxBUkaAI594+mqn69VT51Im4WJZsPlM
sAbWW8J5WoVqRDlEMhLXP0S5XZR4ZaNUcK//FbKB02TLyVb2U9xG2USwWEjoOGcR
MBNMOj6KfNmDAAKZSiBPaeDAZ/xpCr1dGmt4l8IQi4pFmcuHBcpSaVPpkdgQNy3R
zfVXBy8QZ3RzWjBqkmVXNYv1OR/Jtii4nAsN93SB/w5RvKDdXaKEAffNo0gUZP/1
iJLSZlqTljbUBOPk+NFGN3gBC3l/O4Dq/TueSG7YMgvSZc0y6FkP/zVD57eWub6M
h76J4hDXQrqZcQWDYbIY7v7XlU590dHYSkoel6meB7q29uTCQd/WNKa1Ws0vf2JF
NuIsR+l10apMAfHJgKVVeK4qNsMclxIQRodp+EG5XRLllnGP7vlPg02E54DRZTCq
xs7ewmXjoHE9fR68MQAPDCk726UD7CTdZQM6hMoO8DinQEQAJ4w4aR2tlzQvoWnn
jtpWbp/27UQyBbo/XpZo9LcvIk7ZV5erH3K3azcaiD7jiVq8PJ+DcQWM9GMAyTKV
EWjbYfpCoEwYNsu3O+I+B+jUodchYmqxbjwb1IOGhi8hftbKGErElePseuZAvuEg
8MC0NIDpmdt1aKWyNTotBd7owbRhIJ24JW701DfCaJxy50Z6aWmjsalX4Ugwc/Df
2JbuNUZbPlWd+a5PMMb8L8GjrDv9ho4/aIFaAF8SpAE5q7VUvJ4SSCLMrsdmOJRt
stImoE48H9zvvctVKSwA3O9fO/C36UugEpv6vG8ZyaN/xGhX49VJWWRgoku0zZpH
MNRSzgPrVhkttz4s0nMY+oOHiuXNKy/wgVX7abRc9rzeipZQry6/vDZ838KKfv+M
+zPkYL2vkPbuHMyggEbydl4nismjowmt8DkCqQyRWBqtVxh7ZpFIjW5UvSoBlb8j
JYXiE9ciVjKdVz7M9BRlpJ/VNvXtUyLUYq9TrmThLNyzxk806o9OH8BFRLHl+bRA
E97DYzdCn4T5FBKTMQwDoMlj1sqrnvaVpjGH0rStKn64W9ZvgzUuKfG9EzMOSabl
l1hk4e6OMRana5YJljsluCNUhk59YBaeTZBYUC6bPFPKZ8If3rdBgcDxqOdDr9/c
PZbcXYY5//9FUwweBvIG91D6rXVIz/oFQCWzv3EUV3D4wlWWHkD0Pc71fRKU1gTl
DZvU/dNHF5z4aIDMRCDiDWvBnxSBX5HMTxC+d+nrSamZRjOu1TYlid5tZzGnudDL
K6+4Iryv9cydMM/molLbD45j9g7Ith8gQ1GdVTU472tYIBwOA0nVreJ9Y2rzFtOZ
KlypAus+0EYc16tk49X91PfpDgh7s9+YUeAonTpAefzaWR5h/HHN1xPX8xojVNUo
0GeThRaP+s2FqVSMdj8v/de+WPrGAP0EVKWlyrVCa48lvOsI1b5XIbkb8yVasKLH
lxyqp/Ummt49JwqD9PDcH5bmOfDs0P0tO5hAAvIhmc/XaH5PngOEAGmMtlBytgV9
w19QX64kYQokr4LkqauUP1RE9tR6usxlTDHcjrPhMScBkiserq++HCs2kluz/hB8
iF8JviwVIqlh8Wke/7yCvrCF3tig+kXVP2RG5K6OGFTaXwsBDd5YNEuOL/1urNqp
qeAJcxgiDuFt3QojygfhHsIn02Io8P/nLmxTG8s2j0ZAofzGbF2J4uvC4IpllsRy
W93ygIgmagg6LW2kFvoAASvdJeCvGdMyYDoOsVIqGo8K0Z0C3ixbI5mG00qeAcnv
w+m4JJyyV7MBFz4RAoSkB7ih86jmvxumG/mrPTQgmkKTamI8dchdroeqSrtPSgHC
fMjpkYs0Sv8wnQt1dYql1lhNuNOJLdyXsBQM2PH5aCmdj6R2rs03p1gPXS0AbhCb
Q4gVBq22kvTwn8oY7q8rkkz7WuNurtNw2zJiymK/VH3hSD8nQUzVFdI3nopH16Nb
AhnD+9XYC70CfKjcmw7fNleS4e4yK/2/d4Hz1/1QJqHLX7tOqCdLUbJ0ZXrVpTh1
es2grYql5Vjdue4fBNa4hiRQ4oxj6fMLcrgocasXAbJ0kkviYD9kUFftI8DlF8dh
vgDBNDsE8kUlArE/U4bIcAt3tYnKO8BeAi5PHcWfA0iOMBOFBbTQy5tY168s9jwq
CSwpyTtuA5vRsqwIR/mXjYzou8qshCpFJ+P7NIlMCizxs+QRCNDG2q3FauxtcSze
TQYILJcWai4PYoJvo+pah6UkEcUgov4sVZ6tDHsFEf+dzSsZ9qu0HvVQr5WWWVgM
uTlTExEEaU8Hp3tF0XR8a6CuJ+WCDlwyThMzxoXIjtxa91A6kKUpl+OXFwVqo2F0
7Z4z8XxHY9+VLpSbVOyIZq3a4mvmww4dK5TZEHutJlxKhzDmhPPtOcrcx7pZNrkb
aBxCHv/8uCEmoziMfPPOPzEEqoj6mV7LOx1MWelu1iqh5pIELgUNhuc+yk5aiKpr
GSJkSrIrhhy1iWl7Eaqn1LWHkvIuqkpWDTjrEKmtDxLrz/X4BQYhubqe+5RAH9H/
TpzWjv+4WzlbQfX3mMydSdAzGbJ0G8Cd/BsmNsuB0L/XwPdBRElFUrAvkRzIP/rD
utZDJokOg1fpktswOi1AR3mDdeGiIkrvqUsygCoo0cyZIAvrSKgAonzVH+3k2CNh
t4FQ+ZpFs5qR31PTYC7Z7oU9f1JI/0iuuxvD4dLRBe3lleoCUJ91TvixREYt1xcN
t2dp7rM+OYcwtF+zsHoYlhzbvd2fAc1CDgzfZzgB+Dgnt87SrJI4eaNWA7EMXNqG
CvXJa3ZYV5pLsBJWRfSC9D4xBt0PQrAmjCey+s/yTpJxCL8IEJzJS8O2tVWFXT0F
61CLOvTw90+fd23YXAiKCSyfNES+VXAdNXZ5kTtyd48qf2u1EYTc5ClMsDC+W6fU
sIo6DK6811ukgV2Wco0DBVoL7pBelxGo7QYPdcBerwyGRfaXK20ZPua9lZAtHjJr
/MvTdipP0z6kx+kJNpveh96JlKcqTPAr8fumz1uxjvA+4cJYhdy/yP6YUiwRasig
8X1jW7ZCYXJ+iE8uyZkvZO3hISqOAafswpA65QwVkPAJfl82CR8HN4ULl0zSMEv9
oO+vaVozCzb7rRm9GBidLrG9XualCwHngdIk7WIvRy0zqbf9Z6bzl/5FQImPbHzc
NoVj21Ggw+6FLLCcmCoipt7mLtYCVnCWVhpigvdHo7OtL43BI2LklnXKOv/zH7RW
79DPBL8cPeJWu7cKDhteuo4v2Gb8MF7zxK9x3wgm9BTED4HSZ1DZZny3eIVDkJca
rffxxx0+cJK760wzJOLYzNE8B0Fbqf6q1V/p3LUbJODhQLPXxp8pPe5BZQxO2IhT
D61PwA4a2SYBC0ol3ffBZ06BNh9SbRa/KdPqMQrQcoFVRpgzuEZon99hncBFM6Tk
bVkYyj53PbxX5ihdGjCXGQQxawZojWeJ3sWNjEQ4cRu7Lg+vplnC8qSF9Tp736Ch
Sft8Y4Ka2wErbawsQz44SFD3kAJ0G3VSQ+0cJAJgTez3tzNH98+LiWpw5QXXRtZ7
k+GESFWazm+haHGAH8gK9CzaM/fsUKU+HQi9H87aVJDBRZ7h6W13GhRLU6+MKqk1
oDxAmc0E+c9Cqp7Scu2KaBY2sSLbHEfnyAKgAYpVCZfhOE3kR3lVgJn8kzAwWJaE
tra8/G/T6q0HyTFROjmxkwLlU8hfwdCJ7y7qZNk3PcCimU0EsBTwHcqCaQB1E7bG
Dg813W8dQBt0jbVlnIMYp852ZOHc4tZdmYCL0UEUIvSRhrDfYBIYRb2DjVPhy+xH
O7oc0kHKp1k9zSN1L8SBxLg2yoCaVcm017sRoVPwW1G1Ou6QwcV/fL8TyrAAl+Er
2FPiutWatxy9s2cigl+J9DM9q9U3iejDKLYYE5UETJkm27pjZKyNQbjauw/Jg6pT
OzRpDXty8p22PlFAzKIqHxE1hoLAGOtZtorijtkPjGagaVmhotaIMBi5U/79w2j/
m2EShRaBm37iLkMk3pXFkZ74yXBt9PDXumyHs2H0hNcJcpJ7kVJZZp1f0Y4mbsyQ
kV69HvW5bha7TXSZWjxbfMmNcoRWRY7UU6od/UwYoh1pPcK8ZnAz4DKnHsHdX4Em
m0lkVCi8ORjZitTvtx6WXijnMP7ohhzaZQbGKlHYBNgJdJPo4s/pRb8SqNZnUFqp
+jxsro92IV0yd8Ya329Y1ECiU4o3NaFRWjpRKPX88+WO+BiXR2ifKvVsWn/O8vCb
fiY0aGpzSccaWD+UhWoefX9P5tpRQI4jq9nFaYv/U8l5JX0PRrs/XUa5rNmniJiR
tt840D2O6wljcmUxurpjLrZVCVfuAlhZnlSsvRw9CKwONFTJoiyNa/YVj5/x10i4
Fx/28AqAaZh/FVDmFyiMe4I7relVM0uFI3PCrrN7dk5nroD3mtLC4BDQMw9390CV
RZBvjJ/0DjHEAjqg4lQfubcZI0q+4kqNmJFU3ZEwgWxVSC812PXjAsI9U70/DEvd
oQAyoApnMbBH35WBNRhe98wSAXrF/yMdX+n1m1LUy2GJ0quxkobnGkLlvtHJ69AR
GUC0uzAj6hjbjJdA6tiFC8Zs557MeKGUfj88H/UiqHyvCFcDF5Hi2Kw09i+LvDYF
ak+DM0GGkNZz3XzUligY/3ydaHtjOPuL+ExAnT55YPzu+dky0MSgnCvybY9MucyE
lRHuzJb5wqaS33Bb/UG65T7Lsp7Xy3OUvIOGKlVPNf7f83dPTTrFXmNzFp+nYx3x
ESzkc50SyyrIQ8/uNEu2hXSGKVTX1dmWjkOHPdhw9COPFWDx1TQ4otx3HUPWZtY1
6sQ0TlqHtZaDbt0gMHlanpJGk8X5NmuRMAe17/HKurICHFQ8L7QiyoujsRBvmCfB
UQNpenh9V/xKWNWataXICZCNPLAtq3uofKJZHlhgq4gCLTppT1UDTca7d1p3ax0K
cTVrwe4r/hbq8LO1LZ8gYWD0eSyI2ya+PZAjMJrRLbF9No8ASfGHDcxsPJ9liYdr
+o1NbvBR5Jwontg1gNxjT16LhYdMJqAIpZsViqASgwvrk3E1Lain/sicPIGkYmk3
THu/Vy2jRMA5KfNODHi5fq5gz+vUBw6hs3Sh5MNrc3n0iikni6oVfB85QZQXdq8B
9Y/D8QFrlUF2XNw3SvstbkUHbNh7UdF9MeQPSJjoZFJH8MIN29oKnkdWOOyk5yZz
nYyT4sK2VIAX7d3mWjAiuTik3BMjQDcfQzwJIFMKMSjwW7Zb6N+k3z+/ghwnLTg6
ybLWgm+gY1bH+kbCXugC5Mu/JbBJdRuJLg4souTiecbhKwjWWDtuHPmdS7mfHM0/
bcA0AmflR6XBZY2RA39S5mg62nELbupWrr4A73s8UzJPPCK3VtJcscXoCjX2DJed
FvReoWBzyPd+UNak70SQgw+c5F3ZfIohuGF6knx6zakyQF1BVnHpyvStVIZCdFIA
oANqTiQNHnVeZSTGVWnr4vUdUyHZxT2le3kwti8JBl7jyK9rV+dO0gexJeu2eiDG
f6P6+6XgZOFmWN/KANkfZAM1K90Fd04YpXHPexz+XN/ak5YUzRXzUOZOsh2naoHD
ELXK6emPyKhyim2WAUu+MgUqB/ZZzrhK3y4fgDy/V9eGdz6Gb+WaW8KD3sLXFNYA
EXfRiLrOe7+3bfGy773ucaWQtOVQAVvHXL+Ndj82SKwZKzheuL+cRwHZoWixJ3kq
I7hR84rMQQOgQRCaoJjn8cCrfIwmIDdC++CK85YGhJO/uL+M1otURRuLhHwIXdY5
jSkQfimtUpluvMjjYk4BsvrKPKNtQ9ryY99Kj0G9b4saDh7sHnzl/83jG3s0vk6o
S9L1jEAP6sU4mnrKAf2B8CAnXylPqQ+9V8y9OgfUAREjhy1INjgTxxyWu+Gil+O/
8nryDQ80GdTj1xZk05QvgJkcMvPwssiKiVlsLdXXs6ltuuXIeadbbhAUM2KVISL0
RzD+w3po+OKFysfpg7//PzPVc4tyxg0CeBYAHdqGDHMTOot3QIQDsAZ75mQEd3PI
XAVsHvVN8y4IcFtdedH38++TmkYlwqZdGgWqRhUd9yPfaoedK8LWT6Q95P9Gi50W
47xUXzyli2gq9qg98g0YGE74TRncxwGamPr+CqrLhBUusRIA9WV+64gltb93Med/
TsjpNxhnwzS0zBJHObQxzp4MuJADKHCWGFUKG95iNuTWlrxDCE1EGjYxOuEHtvGH
+dxf4cc9cZ0Cvi3d+swo0oVpasxKwcZI3WngIqvefdYMYI92HOL6J/yjYOJm2RQc
ZZAWW7hwnGAlTjqRmqTTrAPb1kTCk+kgotiiGU9Ktp+zgAwwR9z5e4eOL0ruEzGJ
vpLGQROa5B2ZXFAzrPlB94Trqft2JgtMUBIVupYuTQWYTwOsFFg9gBkOGxi/dbfN
m888S9SbdUoj0vp+Hy7hyC2Ww2UnwPjtv4EAMzatrPEiq5Ej9p5vqWJEMS8lcBAB
HZGLPY62iSiz3+/t8aHl+HlBmmjbYgsn+lJydyi9lbJmcVW1p6YhcYG1U0JDV/KS
F0m+9VViK1OSusDed13SSTjVa7FWGK1J5oNyYX2Et+51dJYyq997GpkldcbCpLda
khZobC3CbqVEYgZyMwGwsfzyVSu8yJkY4QX0GvDuwkRIOYeiPU2kZpMTx0Oow8+U
D3JEiwHWnivK9Jpw+I4GXnU9yojee5sYr6jXZZnncbUmgfo/DWAU/LR2IIXtG5nW
XSctvMDqeFzdMibnCiLlkBP42spkrdxcNOQHTJRKa9TWpW2RiV8x9I3I8x0fA4MV
FXRbd42u+1N6Ic+BkZf5y+VKJPYYTBCcxAPZ4GYeaE8/XL+8Ai0xSt2ORym10isj
hhrraBHCr2cGjfKNW0MIhtGLjw1FoRPa0F5JjJ/PfQVwKgh2KLsEFl334hP7QzrA
vwWY+ZHcrObcuo8LcNAVU9U+DQcT0nVak/zoYcbHq2tZhqz1I7QcWP6llX01/e1D
dURgZcvUPfKW7/VBGuW8Sn5VR6OtkvIF0J8n/045zDlbjheCw4PHVClZklTKQvza
syeeYIJMsddRECZcISvlI5Ybpyp1QzIL64AIk2VOLnx/+txcoIYyqzqC8CiS9w9o
6uUgjCrZQWHmAselkhB2ymyQkwcTndG35zGFv2y6i0LJuoNQIP1vTBRSpRaxoco6
VooWahAh1l3h3N77J/qawByTzwL1Ez2OlXtI4SEvkgYVBNI11XNhe5+IRL7Q92w6
/GSuseV0mdqASfl4sZO40TBRVG5nfU72u2rEWStut6+fqvxU6PgxsBA5/Ug6EELK
Ws0wxuTY9Ib0yi4k7aGnj6Q9vLhlIsU+tNtYvFnGj3LtIm/HdvThnOBgeyk0bky7
NDNbdCa26Nrb5jTwaNgWgeWUmq5a2FEP9Y7tGxSIcRpZJiqneEV2k6iC1vxdiY3c
rfDuZqJlAl/0DDRRRt02IHBmq/Fq8C4wJoCul6cli4rdJoEXkrRp1cQD0thbtqFf
y3i1aVMn8rCdXfDZbQx60MW2u1Mw1hXczZcRVBvxYOmDs80QjKq+bny63Fmt7N5I
wXzl8pd7yff0S2FvRPSi45Gb9kqtHKbuApUpI0lzSv3EFVuaR2t109YKMx03ukOl
ET9DgyazOJLgdaw2HPxArY6EraRJIfYlPIyZKDzRPnB1zee4nYUSg3zRbfqOEG28
tnopuB0EH2SgcENzvmavssBOIaGrsq2t+sX9Y1frfY/fJkaVDieEBytaZNI7psBw
dwpbkrUk7w5+CQ/fOL+Z0oBkDyviXhZhdbGvgaoRuARkvhbyMgF7sycP6KiT3pkg
MMBfsMGyfdp6DJzQRoM8GmknwUM+l+lpPbBvcyazJ3zFEK1Nb8PDUWhb1pIfK+DA
gcWJEarWBBBRr9od5eA/sL6irNRg062on95ggySX4+MVbnZmN22MF9jlP4ItiEYN
2GUM41PG2gAfKlcbeHW52Orbtq0/aftACtoXARzswTY4Un5JdNS6gZuqZT86T+ZT
gCGYC4NsRj1x0C7Ai/fkgXOw89FQl/RXCiTj7FYJz1OoVfM1VU4INnAM5Szt4BdA
YmiWwyvxcVZpMH0OCvjiiUDV4uSK38DQnHBujiyZZ0lLyP/aIZ1g1l1SGcvg9PgO
XCfrTgv/ehKJOvyPlSO2UpwiIu+p7KMuTlmWddbaa4/NiAKf5QGM5BBf4O5bOrrY
Q9Bt6scp/Y+nJZSf06KjTp9UXEvIcnLu3UlUhVKmcflsJtEhtpf0VbmvOZ8/b/in
xNpwlVvHO0hfBDS9S6Y3muml8WswDpahbO/i27+qOC7+5qLEoOO2DUlHKQxEX9x+
Fc+x1mcGzBbzhGIg+k6HeRcK22hTF/6O69l2JaFmjCVKPwBj/t5HtBeg1jboWpf4
E1LfSAsT8TIAHTOGJqxeBEfufbuNoKcDnJNt0D+et3njub85H+V9lKHgKWHtXR6q
9yQMklSEpjocWTI1TCRfR2K11NbcjJ/TvD4Npkj6J37SADN0kPcggL1I0UAIZk7e
x5RPzzjfOk8p4Uv5swTS7LvCWNdP0jhR7P3KsrL1j4QbapliMyhYaMb1jQo6mH9U
JyVsJU+D6GtDyEB1DAgsZYjKv2Khcs389N/9JqwJquJzGVvilMweUtgAU/yp6n/K
ljEqVnktYQ9yFbMSZvqdxcmEZsFmSf4F/prFzToXQlcLkK/z7Gc2XacO4DTTQLTn
Dp97rSoEDSSswBRlCxDWQGrmQ4Myu3NGJS4FKJJItZ0WdDNXc/SFK+LbqYK/0lod
lxdymGdL4D7E7gxBEL+JkpIDF9ejMcmi+0PWW+A2zAOHre7azaTHRnTf2sHFLQv6
p9BpsmFtVWhCQEc2eFU9u0MREOnOm1iVf6klOTBlDQs7L6R/q426bV93UDPjODt5
AUmk83xtZdNt4LmsgjNeRtECShUV/Fbo6h6BCxRbGmEc078FVPkZ78tE+zXybRNz
CjT9010rizIlpwU3cFW6r+A6dCxwU3OcvI3PVyyh12Uqvf4yEq/Sp52rJH672GHs
m7yJzrk7JoeOchVx6rUxFBDJjYj/ecwPUTDKOQJVDhz1eHYEb95Z+ZELqwRBAe0D
4gsJkzIQI0v3Ble+5a/Zw26VD+cxNJr9mYSCgbWiFF/oC6djavjEWkH+laI8FuBu
sn/TnsFgqMuFk/mf+emcGyuIaUn1GCVvtMBHHtsLjbS+Rn7sRoY0KzuKlHqWJDc9
7nSyDU/sAifwUHT16qlNlDQveQof4spJ4AFRWglpG1youW5dTc8nctpwTCkNPqfT
OUZ3gqru5KsWI2oppbxvuZMVIEPxnDmz2rCacz3LSxqSMx+tzgyYOpnHLjbEh3bS
aRwjkJMSQXWNsP4UBtmVqE98zPmsfncPdDuQtUUQ5CV6ivkNtGwf/enOtL0CkKX+
EXETnJhaxWYDoURqCaA8vF86Wpm4kM/S6QTwhJV8qX6fnktnPvPOXEE+cprO2oDY
4j8H1K4HvFi2rTsL0t1Mnjo0yLEUffvyTjI4JSI3pzl7WNJDOhZBfpk3DJSlfOjJ
e532et08np5qBpNyAEEvLknVdwDcHwC8ax1P9xnD8o+71ARrgHwV0VoVwy6rG93+
+BGtMWZpB+Oq9QfZC/a2nlTSWyigtKQryYu+si1HlZLB0+AmIF/zESzUPJqoNUt7
12UmUYXBVwSL1GR1rV99cgnK3a2gyvxqBJ3Uytw5IYRzNz0TF+4y6PaKB6/sP5El
9kqjHiUMOd2hrpV5xe7T0sPK5mKEUV36K9S/T4fxJAqiZN1AXOtCbymC6hBOtxbG
fhRFyd4m7KuB/7VqipSh8vPFFC4DBTmblkNN/yWNRLRNqjWBsBJrA5KtWly7Pcq+
x3/7OeB7oJzsAYMUvj2ylqI21xdwjDycNWKtNh4+4Byx05teQ0sXn15Et8W7mrFE
DeQsMUs8+MhprKaT9rL+hDt9IykkSSTvRWyFfGp3vJfbmZpinZjTTX6KXGbOSe9J
ENfpvLt0PF9kkJh4imvheB7fS97zmvumML1YRiK0GjTekimZlA8mpCRPxN6oJegQ
cCdNa03auEQY9WM0tqQuJQubc6c8BKuQOgMXD6AKtDaqpzsbaUh7qA/5dw7n8bwW
j/EtfnuuovjbWTWG1Vfy+FfGtT97p1xM5DSh1FzuRJjSa9GtHo4omWchje10tGFu
xPyWzTKlU8ov3pU7/ZfvKCz8wNgBZz+9rNNlxJQwfbOGaCAxyEIVfAl+JkTjHE4W
6DguuNLhxbz4K8SvairRYVI1XD+OC3dH1ZzR72Sh1dVyOUWXDnk+z/UXDio3eNHh
cArIV21SWyJTavf7oAn5kKrnKK4HCF11J9UjLBxmoz72pmJiJLJpMQNjywOe2Ams
+eBWoRTWTyIM0cgj5wdnI1vwBJ8nKEvwqZpx7oOtXdQcglNCDDMZKqtRpiI/e51t
IEYjlSeEg4lwMISc80UpsLUcyaQI97NPG79G/+3l1GSnZjgf5QFPdn1KTBXZRuzA
c1/VZhifMxpy9h5dO2OC240il/lumGTZoTWl60d522T6IzmxX33OkEg/7ZiDr90Q
nwArZ5k1CzWcUGXBHmKDKo9z+5eQqfU/bNMUFrwNpRqAxGrUG6VN5x0fGOoOUnhT
ifpvNFOoBpaubq0T2xtquCBsKRQ3nf7EAPKvcihrjKPAbDnXhPK7cgVJ/aWulQOL
1TEUf5iiN4zguO0QDGPladef1BX5yp6h2++10O/jmpK1ouPlL6qWR4VaWTZYKpgT
EOgWaBqp1+cu2i/aroW4M5Cz2YIAP29h6BrKfYISc9U7LnhLrf+LwFLyfUCJh4sY
rRloh93ZZGn4hYVwE+spstmjxEhVK5gTSZQkvhXO1GAgZQsZ/pu7FkR3lx4scla8
YTpl2C2PnpIKynxu186ljkLCoYgdi9V0aCcUWSld+tkF8wY6HhFHs/Pc0F1zVecn
u41fwy5S/bGZiyUE7L83tCLV5QQoDymO6xncE2dUtSY6YJEmbRKLQjKi8vpxx5ar
g3mr44q6ha+Lo6WaC2bC+xN+7T5uUZ+i3m4drt430qu+oVwiW1qMT1E4hCmBX9NL
KBJQHFWWQlEbR7pexfJ0HHpJ42meyLcj0xN9D8hQTlr7OxrdmVUc8205r1fBqnq4
eL2BT6MbklOwLijPGbYCRik/6NnSLo0huQOqco6yk7prN1dqqqhVT/mRppDdmj7d
CpWAnR5l5bKjAieqihk8kPKPydFef1i8LcnqdiSoNhNXcGQLxWktvaBsMHMJt1gC
atSDLpar1/sonB0elaDxe0snQC42EOdYO0ZbjCy1mifk2YKPTqDDFjIwOgRJEXsf
wnfRm/Zya6drAQNDggRziadLRKe0lCXBX29CyLxSiMyqu15Nfhi/kSLA/iPQ0HOF
3qq6Xgq074wsdEuO3Hr7FU2RKmkY8l1QBdDuJaRF1ZSklVvQF8B+0+PaYAoSUwMw
J3t0fkM7M477lasewsV/EMK1kOMh63uk0omoJWtyRDMjmtoE/jKQ6cgDujTkSwmf
NNRrkzVv7/6XvGTTckWOF1miPIUXT8lAgIhKVgeaXDlrEVQrVHUGdgK5kgYeGPbv
C1bMDiYjhylMdF6lX8aHMAUkSxa7AkPfQoa0yes4NFyPisuv0m1veUZZAWbsq2Dg
GWUYVQomgpR15CghdUUPxESoKgfcGKZU2UWD5zYcCCwKXOsHrU/w1cTWAOPCT4mC
7d+EIwE9QGxYdCUfKTya+vJYxpIckUty2g5vJN33My2oNf+i9bu364p6t5wazsSZ
vPd1BNhua7gmvMpCVDUANKBv0soOT8J1NRJ1C5OYahNfsuSrcV3n5oI1Yf/34SqP
2t/NjwEvv8W8flaWp41VW+c3y3Wt6UpehBhUREUEXqgHodzsmkhjl6Tdu6WrV2Vo
HFMh4QsW42i1Uan7gXKuvvLPEvhrpRh8npwOfxcLOAM9S0zrcZ+onu1mnXtfNp3R
Q2J3J2SvOh87on5q99H+AJZyndczZXR0BDBDEBcVB8C3wLAevYXABZWZVl63gKG1
RuhcvsPfumiryevxxu8A7+TV6ddB9Nwib6gB4O+JxRw54RxFvBku4JtPJLwZtJPx
P4OTnzfZTgoF1bUjvxhrySCxeZ1V7MDiUmaFpuG9yvsPA8Pg6VlXpEVx7ICumT9S
0rc1CV2zCZmFX6zueW8lug+gh5Bkun8M70ARZEC+mnxZq+iHBq1DYu2CouXfGxPK
8nuVNpyBfYvmbPKQ1K7v2rT/zB4QnZRVMbXyRv3Sr70Ujepx60lBoAT84SwiwWd6
wy+XqVq4lVe4nofAZ7g01Wj2q1p07f5SWOu0N8uvVbzuJe2kWjtsWdqUB2bzIWI3
cARGARLpeYCimYwKaO0W0YfuBHmJZm4h/ZFtXY+xCd0S9qo6Z5v3a5HLi4ovn/Z7
29zPSj+2Mrkb+Gxlrnjp5Iwf/83kbOtuo3gNq3PCsdYr117uE86oncBU3OhhOgvx
IpTavRtyZoJl+fZWSmDzye9sYtdgLLnlhGitoqz8m/ixqVgZJeciZvKdviGPodGd
UmQGuclc+nKPkjGAs3NWMcfAVI8OJHZfQiQP+ZQx6gLEovFbC3+tTIcfjKYrUuTK
DflFnPp3I4i03k7T9x/Z9vmgANogonrVRcsQg4KaKc7Jl37l1978pBHw+dA4axYe
QGos0g7/QZACfA87tvjGSJjlGRS3tjs750p70n43/gvMDpAJMxAAKabloIZjcVsv
EAjMb5H62wmFVnIVaPljQfFu88vLs21h+JzuQUPK3/+raklUt+JpgvgbvCngPnAu
IWPtGPyTN8XmIow1erQ7eiMz9iCp2Ccs+hYGmqBRkfxL8SMbFnhRu9fWpTCAXQIh
ovz7If6oU9+8McSZ7NP1lBQuM2CYgKk6UWBlAoed/Z2AbIf26X4gSFtyUXGCs89/
KDXORWvnEdBaAqLTsOYoOR4H37ie6Yc4XOZB0FVVfX3BJRNYdH+L3nqaViDHaiOj
UjEKQftDwiZp2GePyrbhu61xLKO1Nja4dz3DUIEUiHBKUqhbWE46cW+c25GhG+vN
q5GSaF+/J8Npi7K18Rwp+4cjqj4hh9aceKvBXdGX3JtCdMQP/lkHxY90pyadHDkk
TuReawizcMgPjADhdCHQKakHHfgZB/iVgEIRBNxG5UNtMYBaTRAiJy0t6zfRPuV+
kSYQVo2hL4vUh6D8SQl60G/RQGDI7JeuPBlZQ1M1QcObQlSUUqhQzLv8O1Z1bOZz
t1znoFTYd4qxTn89GoalHWVhkzB6cQsFexdlWauLbykxLeUfFga2drAYv+3EGnnv
fR1Y7AsMdq44WvEBZ9AbWgN2nG46tpQxNVsrc3MthFZXE1x3lkB30Z6XuUz2XQu0
1repvpanUSqG9qih7HiEcxcoD88ly7U3YVX6HTHk3A6qphusSe/Goxbem3Aaox+c
7QK44VcnBNTaBOyiaXRah4EvQKWnDG1BIGn5n39KSFvl3h902TTakN7PlI1bIkgq
DIFbzlXYlBuFNpQijWKhBp0MVVr+PCELa0q31ahdXXGTNT4aqz/Ge+Yyqqh6Rahf
UkaOA5bdBxuql3kipj6hwmY/IrY30nJ6mnu7uQWP5//coc/N3enxIrooY4tf9jww
7yvNCpm0qSmHyNh/5u69SXP+Zdy/gtjyR6wox8QsJ99Fjy5lsaw5RVf4izdqRUlz
iOmRUzH+ZcaScjp4HYVLZSsxVJ44JvFvTBaZODHD3Lvv3X9NJLUvEQcKvtQxWg8Z
PowtUrRnrXlNSehjkCH3E7msPRNWiA5JHXvGR7bYGtIBIH2bc3oNu5Xkq2t/BBou
NPUtA1m6oXS6wiLiIEiBLSEK0usLbwikTfftjLzTvsXtC+foxNEDLz+G9yVfpanA
MPN9rmnGkl0Cgnt3vnTv3ZDpLGrceL6JYMo9LyKEuHBVQxDaDwMwyRhM0TFRZ0xF
gg45dKKgUHAVAhUcTviAGZ8RJ542LMwAwfLaB7BxGccjbGZ3PSjUJLNSiWFi/tk5
LrA7G62DnSIP8D80o8w5SGvt78GNmwHx1zXnuRw6MJi7kpQsqs5uO69ytAXil8ld
mmm80vyZWxZ7arOx8GQWQsCH4SQnMUmN5WcU8kR3GNsgExLz9mKbkh4G39XxAcht
LPn7mIzgmLG5pYZhu8be6B7hYTU9D0UUNDT3xzYLV2xuPjyEJgW+PZyEyppyrzXk
lt751iCLg77ex0PcrAQXi/e18gG8R1Eu1FvObj8a8i+LUGT1LwWw+u6Y5yaGoY/6
JPkbtE2b9V/rR+YF8Wd/Nsr+gW17a6XoehcYZptb0rgV53nHvvhY9eidkvFdJItA
y9AGqJiOCpKBbKdEzRzNodNYWOlx9faygnY/17BjR5jtYBFDpz15YVzimCDO/uOf
goDoGwwqBKpULgRKmf7hxza7DOCqwRrhzAEqF405Wg4wlSWjnqejUbWFvOp2NVoR
Q/Sz0BOo5E/PhyjYDq6nVlXqeUli+/WU7SBQOre0ZBtl0WnyHAu5dDxf5hMiH31g
Sf5+6DqawOdRC3eO9/S4LhLJmcR1ZmJHgXT0koiKHFOSg5GT4kkM2jA9Bt/Ib4vN
L8e+5uKW/lvLMOvzG3IMekDt+omLMI3C5JqYOzcCGQxcg6WD6oKpaDPyr9HckVzx
dXqEnJvyNPEV8uw72+gQMArXkSCOx6AkA1fptJUwgWnNe4D+S+BsZ4Y8b4BrBWCW
BvDxLL6tAGEMBArNnL1uBJfnAeexm+TjYw+B5aCtu+X8HX/QSaY4c/yQbgO35Pfg
xIHwCoclhPEKJV2ZvBfONwFJq6pJftEPZri2ut2M/IynvWdacZbVd4DOSp+Dh9bo
QpjSRSKxWqFBZP9irltQimIO1k38YDfmiukvaYs6h2dkdHneHNZFlSiuh4OhteMu
qTsnHN0Mi8fYNurbDBpcZWUeS/WSNf0D3VGvQCk6fF0QWb3x+L16hsvws3I1hCf8
GrvLD8AKyus0R0AddZhFn9/pmFGtGKx+6E8UaqpZ+XAJ/0o2y/vQzuRxOSNSkRpe
zHUuiMqW4Cf2hBkaxhu3lCk52D3vFziE+bcYigMvkTiIsVIFJLyBVISXxImp0b55
698u6uKgnasf+90ufOMqGCd2uFkeilFe2p70OFXqgsV2O5afKR3Wqn9dcGu6PyaW
+shTlMKRmsj3x5z4x8Ds4Lh9Ho+3HCu0Eqcmu0YbOTaIELu/Mm+88abpZnzlDq2W
yFKrwSRXqfESNigPTZ5vGBLHxf7rkH5+yLfhIC0NM+ln66cXN7QfJWF04njCvGqN
gBAbUF7C/5woMzwSQyNiRFkxX+f8xnhgfOTf1SrYbQba/x1xoyAsuoswo51zag9M
yfrAJp6lJrkrfWz3ZLZpyXNEu8/rqkesnvuZqrraQ+b14Xs3u7iEThE/p6lKir5q
hSzQFGk5NARsVAUzLwIDW2bNQTWXMh1gCt2WvvJOKeYwL6yAX8mRxmDGH1W+yPl5
cHu6M2wZyr4N/jSdbEdiE+ybsh6F9Zc48wnjgymvTVF9HbQqmfRgSrWdgRQgEbwJ
B8YJQ78zNnAJnrr9cviwohnGrgUla91ojPgsJRjBTVIeESRJ1gn02czksWB6wqA0
lNy3vJQetUTp70bDnoCRfCtblbeqk7UtM3n8tZWWpwvu7mN5wtrV4ba6oI8J+375
WddyjLSPHn5uJZR/DygDR0iuRXralJL2HLPMwvXoL7//nZKtd0c0D2taEgXXv6so
oIjFnb5rR5i3O4zouImB23PLG3fmdBjrwZ6ZIMqWN9lfuypvYNsvin3q+HwKOa+f
0OVdF5apBh1qfbMA0CFZiVe2nwFrApaUWtxuf9mxbB5sKE/ZMD0Q2uLyfKxpX5/6
xiutahNixlQJlbJPZbaGHGjEdHi8m1UD26Loj1jlnM1nDQqIle4av3qTcsd9zir2
a6Zv/9b3eUmiU2nEYzmZK0bfJqxD9y/pWe7GjkqKYapbuRVxpBavemhMam/LNO/e
o1mTTwedNYoKxFsnBU/NfYRxqzpE7bjZPsNltZc57rSb3QFcyG4He6T28UmD8e7a
7ISt6r5EoxzWPgFZB3Cye96jyLYt+GrmxTYiUb8wOmVp5jp02my/OmG4e35LcKXX
GyZ0taSX4L5tQzASkv3eziOLOpT17EAOzpwudyNXARviusYgObG3NJQgXQTSjh37
+ZgmPhoVFR/UCcFPqJsuFSQpctpn8wCEFdFLEFtXJhPvDCaMZfmnQB8WUnOq7xdl
8Q8e4jpj00s6sOLrABB7rbDZ4phC1Kerrb2O8UCe7xLJx2TNj654QIgWULw1Ngn/
2WNWp2ooPeyDCTrmH3DuhDL5wu5/EWWSNq4Gm7jYnVjMAlf7MaZ8UsZ0GrQlHVnP
iCPSmq18GKqT6ap+sY9lgna0e/TfxeIKnPUiJO/Wz8ARkjwPxGgvfrUj4qIzdVIm
TB3o50B+o6u4527VQTjjy24s/xldc1nrq8D3Nj8U3nuazBQMjg8ZH6MiFD28DEq+
pwBGG4cuHkRCbfzJCy5bHD1tNgKMiHBbhjVTJu9n6Ny/FIuoS3cgKSPCQbtOeCni
kWIYK+7g/cUs+js6dcta2ezq2+4J1HqdiYablqBVuC8yBO8FGOHghkCU6q6MN8t2
PgdwV9LiZTwxqzry1obhYZ+JwWQtBG8V2ZTOF5f/RS/UnH52f4I21QIFJ6QKvTh9
w2qt1zcB8C1PZxYWo0V71z9s9hG0QMNFeEgfnbjXX+FMQpyhgNpADVThPbBCRCN6
fzBqTj+JF6tLd1rf5m1CUygBEYjqN//p0naBTI+6qUROg8P3QYS76gX2sBct0JBU
erKnIqTXrVTuA4TMWpwlxyYGbfivCA8RL92/BOJeo+Ck4kmt28Q9OPeoFy6xTm7K
uniW1b5MDvL+hW0owK3nesZ5xnaJuTf0MTnrhR5oYxEa9zwMhuHW0MJTUhe1ExeR
q1/JcyhkaPI8nc+3rda5qYO0FUXIg3TxVw1BEfMy7aLFKwI/ymqh2EPNNTREUvDe
pSs2EIBdpmC9cnB9JyxPTix3zJ90tpF1Uxo1iysrIwQ3j170IQkM8gXLE+yfLrI6
8oRgJ7P+3145nhop6r8NjhYisq8q9LueXaE+/8LJoYQDl0WkVblBXWoBCmxsTnyq
cJKGuNF1uHvqhw2GhZRTBXlcM65joionHq13Jdhme6HcD1DOKtrrRC4gHiteZ1pK
OUbQAxiGoao+MOkXgLo082KJSbSGTa6/4ceb1URJ2QCYxavcpfl5l0Zqz8svPk5B
6qPwVatvCGOZlbQujZNjgrnIsLglwcpL51rw8XvQ4dhQGIWuwBDhHQsewk6peu9m
rFaH8VVdKCEGMea9MxZK+dRCO3IrzUiridfeJJeuaMtLVmmNezM59KrIquayxptW
1UGBe52NGrvmLPC+FAnFM1G+vDWdrl668NjC9eBI8p7NGdeGPfyrfKnirzVp2nP+
iDAMwRAf8mJHrGwoNJT620XmmwNMJFJuIaKwgeYANOefsZbuFKwHy21wYY5FKUdt
STbo9PYTAd7a2Grmu387ahOSd3vIi61/v4x+DhTh0C80YM3wua537e912w+FwqjR
9qCuKfcRc9gGVadhzPXEs+pNZGAo6OJYNRuvVYRBbx42h0x7hFJc2YYrHtrC7ruV
M6viRufWH1mWhbbfB4i31ER/nHs/h8Cs4/31bgNYbtd9qqpJ+MfrzuS5grsu8w6A
o5+E+8zlaUdxDX8oO2TMchg5cTrhcoprr8G/l3FB2NYzWFjQhGR0/NlwAbBD1jas
kMuRvQuAefREgpNn+2RdC+cQ/IsSsM8d70zhW5QNbNHzO6kUIyrLZF13bt12E7Ez
ByTshnVH0vPNjjrHlZHV+DcfPyL67FGGjKsSr4DwE1d3D7vp30hYZNSMaN4o61aJ
QIXycnWlfddoU4WRLFx48KXSQFGQOTlg7olfed2E48SnOJd6/9jN+6Yo186qgWWE
O5xdtm0Xg46yE3y8owlygwP/Yp7JH9l2PP1zGiRRGqS7AjxTunsVVDI7FC8ET61/
Fnf2CJQicBD7deYZdgtkMpgk3VYxAUGBHiUUbd1wWlxbpyj2y0LPFXU0UVCb7YhO
XViUIG+yFGwXlEGOWbwKXkxOIKDOGhJimpQpYDPkB71ixFkZBjyNHZrSNqKqCcJX
J1+Yqn1V6b/mkaRIhefpX8FGm3y1v+8d3E1jtzbLYMxi0lV1A7dehVtxkSjZ2znq
WpQ9pmi+zR8WTHvrL0psLohtgVVpbYvSzXGC3LAUiXZQZjskv8NzXqHTkShKHfSd
HNOQw5Y6E1ejM0JVUKBI/RvPgnSmfJK2v4EcPIDgdFIzPUGW+k2Xwv0OXVXq+7pZ
M1mKPWXWxUee7Q/0SeYh7H5nPz1XaEtWvS1n/Z5blv6vdAaGApbhZxI+ZLDkRJLS
1gRUX8wjTI0GavxsROfUaUC01SxlMPGE2eqiqOHrlvtKDLoyt8ehAGGRSJd+nL1n
10ygTE9eoGgPejra3Fh+aj+vSGUmOiTG/l9G+qQ3YWI0+qRz5GAxe9JXFLmqtpVE
N4RZDqURbLlP/2ytIi38V19N+UWXEicXx4MZhit89v89T8ebVpwQmmEKPio0BW2P
397oPoSqttIUqQihkXrpNEqVGs5wVZz3OjWGfQ+aXRNjYJRvFWGi4SZmGC7lymjc
3zwKMoWX4hk3JrLbI4EA6k0YYGTxJ0h/hVBi0NkJAiUOEoA1mF/69KoKKso+/QH2
SMwf2o+Y7clkEzDRoL8ayrnfCit64COeW1jntMUQbPEle70mwhUGmA6EQFHL+kmH
8IIE0U9xV3jFgdU/qqK66uCYmigFHvJ7+dXG9crm3Q/EzByq6KBmWAMWi/upmpoO
9oLHmBSfw1/yNN3Q7UAFUZGF0Uzz9eIcNhTjUQO4cq80lpi2LUPd0oKWrFi+gTLI
gGMZqj3jY3Lnpmw7ylKvd1WcWSNkRcLiyNXeKpW5PhJhoCv8zorpUkK8/ZqJCwbV
uwmLhH41eK9KROKnhwwDvo7TDrkqgmTZltO4absC2Hp5BnzdxUXaWOaZamB3zkJC
MJ6zeZi5QvcviyqDANIB0GJ8ehCRg1RYdL6rXrXp/dZfkrgLKkSV3igmkliV05il
aUTLXlIr/HIY2SG+r9ndujKyzVR8nkzvcw+nmdhvF/+IZKmBo/pMc4nrDF4ArOf5
bthneqzFo7hPz6Wdm6uxRnoVDpPJzsdGSjhv5YBMHlJSbJU3HEwRjubhn8BNe1nS
hDASxcBAlG7cZBiqVYX4kxJLe1QnN3CU4OB757kfDbrF3B8ZsXOcI6dgvtNScUYP
Au/0stnmPTymT7TRIJp4BbfB3nCbWrnY1Qx2bxZcNYVDv21gt5Hql35u+K8Ag1Ke
ymYAOfgmPUL2GD4qLOZrirzHLI6Eb2jH3U1ZOv8fTUBHEHV6wLLssvLAdWUDVWc6
smCYPysdVDjMf80zxVOzROkqt4m257f80lPHArgtakWxB2UqrX/owe0yDWhv3Um1
3L2rDNyBqe048VaP+ibm925ANtNZcKa/WMcD0xoIxI9hf2oHwe8hL3rSaWt0F31f
3ol2hHp6ag57W2YtMFEZf/Ox2vR89BUYLOxykGBmldrFpoGDHKb6Jiuuuj4XIqqR
mtfy+dZh+T20yDe+fnzGh2a2cmGoooEWZAJm5o3VpK4KZ9EsNflSyDC1Slo018hn
Vq6GDEFNewmTpfapXAOxUTUewu8Uo3f9Zm84aq4KezzNsIXEQkUKo6MxO3Ds2aaQ
rISLCjLQQczCqjagZJAF+c3GXaWyffZMI8BS/fUmGkE/OweNw53A7wKLpe4Qnu27
Bvr2F4MCND9R+Rm0E5BTRmnFNomxnnPloFK/E4YCf8pu1RaOiZ8LScUZMidO9ZaO
SnCJMa4VlRYv9UD3QNoHH2VEMnc/mDnGRoEoB6w3GcE6mHFd5VYJlEhtqYSbUy2/
xQnzJ4jikQL0J1lkR6b7owd690fwDfKFqkcEGYYEp7VkEquge07KTqix36BE3ti2
LrNrXlhHCPBr8zY+izJBJ6uFI7LaU0hdxoAJHesHqod1DwRT2AstnQmpRfv1WB7O
6z55XcrVKXQSqBzFSqAy8aPQyOZDA91fuoUwv2cTZf6D3PUiBDThvEEGP4P9wUrN
iMiMn1ykPi3ojA6skOyMscRNJG+hYNS5j//+bW6nTiZJoxkPsLyxsyQndMLgfMi5
8VIBXDMGO/qqOMsQNV2cbJgna1AT5M5oUsGsuObWJGu0bT0i5i+o54iRpucwrsJB
ij/ZvUE+KKOLyWlK+jupzcMLjQt94p3Nj4hNysabUuVIQlf+AA/aLooYgXBE9pdt
3mTsr2LHG575th5nGGyKRjj5mippoOcWLc3fxGOyYKX3Uj3vt7wYFh3eWbCkzWbi
uiQMGCSxrX2qh0rHkIobrivASQU5PU/2GTkWAhyjZZmUFAl6prKmkgryqt7bWF9+
jo+t+G20EhByBWK3hRAK+dpvqskepHacCWC1dNDI10jIXZsL63dT8UTfEwTmcz8J
GWAe4Rn8Kmm5CtZyD7WmE04i0DCLJPCU2ilg+s4QHa++JD6T4nxCOvfuEwCR9FwE
bYydC9SzolfNaHAu4zPEF6b0LYN4R3d00b5C6OtSvWlOZS9dV1JtsPFEa+2hdnjO
nik7YXzBJRK/v+T9N07q49UGRm8q2nB8G/rVkH7Jh6tFG02OwdJyoUvKZIT0meR7
ORQz6NtiyMCPsnb4u36mDalqfZnaTnHQxH++IGjHL2G+zDzJhTkGyyUwrftoLVtE
ZDhkuAZnJvmjVUli1XXnaCE1BzSW6t5s96PONFEeVkd9z+pKTIkUKHk2NJCiyVG/
eOJPzYqgb8mB8plWzCY/JpRWLgfVTMAXZa0WCFtSbH1cPxhg6cHHpgNxXPJga4gk
RmDNWbmCXI6W+jhHRpHrf66PSNZehxxn04CsmAyx9LmndtmHNJzuPrAgtbO1xj3x
ljBB+k+NWhp43pAgC8ums9E9fcvK5Rqrz13JcwheIUixq0VTYRLj7rOjbTRD1UjX
129d9PEGcW5X2ZZsKH3z9c01T7EoniCnTGvMc3DH6Sc5Skn6VWkJnpa/KGw8XyPx
kViVzq58mNYsiFrRi3CLFl/3TV5m3q61nNYLpzsEIZ9G99kGDbZP0eSRzE8KCGJj
khq7DCefj2xatGggIXylOohf/xNdLOYzlCSslz+OsqpJwTfsFUwtYHAW3Urc4u40
tpTsg3Ie3hdRNbpzP54hdQZVPuN1nH3AK7xwBtGUli92WRGHtwXGcGmar7kruBqF
iG7S+8UE+FgaYgz07hTcig4oKM0d3tOv7cgOeAMSV2Qnz3/24hAk7eHcTNHmrdzB
oS3NMcGVlSTE7d70LJ8+uETblE7q3zl0MpJ00C83Qxg29obpVOAFQY01vAnOQwym
WBC3kuM0h/TPWKyDApgVLCOj1CtNbFtEfTNoHRodLRl+3eVJdPUNiyNX+A4YuIPT
vCa5/6o/j47AB4mU+2CuN/34t8epEUp3CAoB/cHoNQ4pwqqSszz4y1sJ5Mi095pW
bY2vD1iSsaPipaLDp+K82XOzDtqKw4jda5W9sil6eBqR+RqY6haQY0U7fPWnNolR
PIzkmFHjgdBElaTu8RFZwyNVZS2PKd8n9AvKqXdzwyaMxq/hkl5EBmWsKCo07Tf7
YjsNcYffHxW/1ZxlxlPuxQWm+8G/i2M0BjbKxuQNQEqiqxf/qsYonKREE7WIpNFA
huZz04lXDdfiy81x3W0mqFW0pX//3Zh45fu/bv6/avUwECX/UABmhu7OjZgMc3bS
LGActKFSU7SUTyUJyOuCoz8qlimxuqspIjyohLaeIVYQ3PWJVGr1BtIqkhzCkMv2
ginPGXfSNs6hX0VOexTF5cgUTNmMPcZi6QdIWb4WKbEFyykQ7cAEu5Jt+25ylXpp
ilI+ICwQCpkdZXnRqZs8dJ2pwpsjP1m+8yr5VJ7yI4ohG8ebHi9WySPQsxncWiT5
GpfNy6Y/m4kCvX/kTDGj0z5gWOWC2F/0dCIMvjvgWW0OpatMXByRFJg6+/zCtbG4
GyGtRkyonQ2FlHK0o0EQL4G0qPxBBwDtyJDmOR4vTR4vk70/ExHvXEZnmrVxlYHD
fzIyRtVsD6ErsRTmfoeiYrHXIft80kvH2H+KiOgReK2IhkXvQXL37tWF1K2UwimR
FBFNWiU14KTaeh0kvu5iEzrx7A867bdaNWDScf57a5XesZPjiyk8d/DarD4UT0a6
eKEZkAxF7yYlXxVm4mGwddNszFQrHkty9TSYkL8+WuwkmJcTmFC1+EuY1WrPuwrY
9DX7qtv+e1aL/+NUjx4eHLUOn5ExsVgGnKW5dqegPEy1V/broOLxM+LKNV//sxLX
E6fTp+qtagmnN87Hi0QD9Zwvd4oHkvtf1wHn+kpTO9/JCuwSXGAwjk19s7Jjxr75
c5Ch1hRidTvuWoQzCZfkaTNCwFTXlb+M0zD0Z3K6eKBEDiI5bZHn8jAgPCtSRTD/
QPPGdDQvAFaZdsPo4CYOZZ95Zo37sUd/IP3jPKlJt5vaRYkzdnMK2+HjvRxCjeBJ
326JDOddLrg9bNJX0giB63VnKHRI/8dWuUit7JswrivAMCjXSQJkRKdZxQqfjR0x
DTlW+Bl7FNfSjF8WqpGy/WFuxCQwLkDmnlp9I9JY9eNfbEGvDS75c5+0ns/t5bDc
IXScy6Vx+n59YUK6qh6aBYPK9bN70dD5vsVFyScJGmq+KESP8iaJvfmrFZTdZEkx
yY5E6qGPkhOkq//UCJg4fLqJASC2EeRgNXNpzgcZrcgKHcMZtrzOuCzHcDkdzDrg
peWrzugIMh8EhDx/m4GR4tyO+dbWYFteGfe5i7XnW5uR6jrWBu2klkzit7b8gLoU
pjuqxdIwkdMXUmbZZFDxPMraIEG8vXAGeHjTGA4ML9S/8W1PdR7lzXgwq49qTYuT
y1YQ+TNSNS6GuBQMkV1840ODxKTBGXibMYFyj1U8K586GqmxQdxjzlIzNvA4y2d6
sjMuvgk7e6NBpDNWUhllT//E47ppGCQm59RgmZf8xfteV8WhwtsIdezVVekto9Hw
J4iQQISfhbP9rYJI7Tn7cCL1nDOw9RcVfrUrckvg3x04SEgViXsA25+rEqm1Q953
sldNJoj8Ech/7qoC14SiFCvnelmeQe85Ert4vw9s+CM8CsqIhd/yucNROgqf+0UG
uXowiWSBEZdwNvHhidcfJH0xSQw0qCzrEvCZ0UuWMLPo0GTUBEhckWmo+ljR0qwp
/mJ442K2L05U4Qg6nOOT+Irp7POAA49iEEcjyeF0zqPuvyl1Tal9xNiYlMj2AEyV
HvoqiXt/sNsa3+drNXMrA+JXDXAHVuEK/7Q7g/Xn6Q7WaV9NAmhbJ7zNdnyu4CrJ
KbOiprQfkVcayxHlWypc8S1D7q3UdVaiJHPojk7kfnBPUKIjV50iOC8AtcZ+s3F5
sA8cywS5YhNS23j5W6WLMtlcBYq0+0rV7AirOkOy1YboavrbxiWOxzN0e85Fmyp1
iKofSqWte4XROF5uk1+YSfolXJcra0wyDUeujVmuYoQWmVC+LUbJ5oaOSZIYwYnG
p2IFOcczgEqJ7Q6T+WJ5Nilg7TgVMMhX8QmehTYsCEW2lzd8ixW6zMizbws2ydQg
3HRmFEu4rGJ2qN5ePPS8Dlm44RxQK4/r+CAuQBsS2PRorcTlKUf+VbEX4INngyh6
ia8X7Qk/TsS6+mNLzP0AeymAGXGQzKThs671qorFMNDAWPplc5iTd3HK9v1kwgMh
dMtKNwBY2YgXqPoksLWkAn8diRlGymOGtMIYkmI2ltYbTW+hNFBZ8OiVSqfoUAVS
z8keUliHlLZdDgoJCBXg999WyQOIRe5ef7rL6P4o0Em0sr6wP8lZoto2Km1K68Nm
HXyyOnoK5YtViTA28q4/WsysMBE26OEXBDcGsZw/n52SfJMkYuPEvDjaFZXTA/po
BNN4NFsJW1pHYNtL3mKX2E5um17PzocvOTJC2MzJq4qr1YlH9lc/Jjh8pGz5nxyp
B9uOrUH92iLRIeghZz6hqHfO1g3ArwKhXaHMS7Y2mg/5ixSzOtyOlHqd0i0vgFU1
CrfYZn2qrMKCQElaw2uQmpOr132zSJTJUu4V3sKSc/Ze6/ujZ+n6gm6etTW4HYRs
+/3qoBA6l6IsKe1S9QW+gYEXKjOdj4QXsQQvzjCBgt0MKzeEzTL8LGksMvzcNoQA
aoaMXjcjWMOo78K57NxhOwEXGU7EIlNnc1Y8tvhEoa/XzRkuBHZKgizA58+ITZJG
04BAd5omf62tl140IJ68MpAD9PQYd+r1jRaBX7DmHrgVNMKK5DamNUuXMbKOi7ZO
3ogzmNziWEyhZmd9dG+qyeMuGumItk8UhdRsgpZSfSx0QQ5wt9WCy6/BiAyIgMZb
3dDs24FlcX3J35lsbCeNRiehO9Z1bYiwrWt1R6bVfZLcrYOk84cPqxxpGq7A9Pay
c+wnIUE2P14hTkuprjIeyPMifFgc4W0edZb42dUJYiOc2wN8lidJEBwqLT37TaeR
NVS5pNZeEAg+MDvm3NhydW+snKFTBFwOdQZ8b62UKxeNygkfLXdvf5qlDTEOtsbM
0/2Tlb1hwHU4bzlYkRkGWIwzBprZHQZY1LogPL/1RSHbXSRzw8d0vK0zM8TgUJqL
BBw7w13P2EQXxIEXZuyHQnQ1/XmehfXYmQACDjvpnlM56BI6LODEqPhimKTrxkut
7INolEqDdZO75cf4wtOw1/M7fTM8bk0BMemtSMzGMVU4v5UGkjak4zlSqOxD3ZjZ
MYqrdMp5BTFdcVfPT2WU223z5ze4SQygv7dUIsYUWUdrUA4iofv1du6sKcpEnhrf
zEa3cUtmrQzvMqSwi2GhZgymgwjfEuQpu8i5XGA8I6TsbkZxb4dmamVtAfBTc0sh
da/Eog0XMFwoubEimyz7NFq2RPMfc5VOCre/xREgSbPqdlddJLt126n4zrCqst5j
137Y5LwiYVl+4rBNsbY5Kv+SmHJte7B+TxeX5ozpNQhb5xwsI67E4XYLcs+9hjaq
47cB7RjL7NVXTLKHoI9jn2tbI4ncghPnBqjqxdFNUMOje5fg/UvlyWeSy2cW+tZt
/5zt52Hkew8R5GdhM1J2bHY7Usp0y+C0fnGy3OrGu6n4Jeorsca11U9P+UK5sCQc
ufYz4Wc/XY/I6g7TPkyWbU6K+Q8ulNuXokPpPjZyJQIJ7/AvpepiLmQ8zxIIDBSi
iBxag3NYIteZdwG284W8C7OEoRxQt3Spk9u2fxwRWMfACb8shDbxeX6whJ7fZpOo
niCEH9pXuMeBW6MQqB/6Ic97VAevAfw8ltYNvxLHdqxLqMXnGMp337VCXCh2TxWV
lOXFzX2JoBXRuzdMX5YEefp+jaZ5xmLPqZl3MCWzbZ4Y5r402Figu5npoQ7uxEFB
Dgfp5cUiI+BkYEc5fzM+UDluhSXtmEUD3UMWY3yVkuL5vHK1dj8owMFxjC/Gwv/7
sIklA0gDVhnsHqTb+qZLcArbLV0J3Z4tzrUaPQ2TtPFXLcFuZbDNCtYlwDYES1JL
VGTBptnrZ6hDj3dtJuXvW/rd5BzIPYsf6AdUB33shopTlBocE1QOeZrf2ozpPikx
/shpAViaa3CnwlBhAMim2hABedGoNmz//m/g8Ui0Rn5oHdd11U57Y5Q4AYFEdccD
ycZaEgE9//sRH4BIaj1qyEuf5jX72J76rWHPz9WT7IBv5FM5gE4IxJ8mkqQf5XIe
puYno0h9uEm13HeZ7QPLZ7tJKX9Iso2yt3Nn/tlRwMnzhtr2YneOxUrsEUOUWaxX
Qya0E6wFwLBuOUqD48YfZ0YcUi8baYCQaL44Jo0a7pbowWEIX6ySWVSTQVZ7MN3M
q+jsU0maVD2Gi0wPTDMAep7KBJObXab45nmjQcA1Qlb5KW4FqWrbbs+vv+KPK9+n
1lC8DJYmQAjnkm/C+bfZRPWNzL9+rD/ZifS8VPZrV3EaTu0hw462+lEEfjSvOYZR
mZym4f/UsO5H21y7gdJejkG+TOISf6hfsoDj274Bnk7FZNWKkQq6qhBmwjiFYiU5
L9aE1vtGjPmSzzrZFRDlFjdhUGciErTOEkgfZj7r2pY+WLHgXXUvw4mB5AxhN/Bq
qcMDhgqV1oCNKOIjeRjSbSl5DJqXzSEVxwCQphdSTzkBwX1akiWCOzP6dW30R18I
PGsCouk3qPem+e09kAIwDW1YI1wTJzkyUGtNsqcLGEE6p+LSUkqzs/N6srZXwreS
a4iQRPHGHbsi0NTzRfYKifHUtrKDg10+P//kVqsiU8QDZ3Op6NEG6drQjrJdgITX
Vivz8W/wflRJu7nBoiqmqX1svInbzemsVtrxcDB4JgA/bnJZeZGuYPYLSXUn9hmh
E6kZu5QE4M4ne41+jwFMG9KKy7ppeVkONEZZ1YzceMw5i3KuptGhqNdzoDAibFbk
bOI3N73gkZYNkE0bW8hcH0LMu7BfcE7yCpoyHuew8P5igCcEcJNN5Mck3DF1Nl0V
Qo9yhdwdAEb16vt43cWcBc9AEu19KUa7qctTUN0xbxKzLaPGZwCv3CmjFv7yarpM
HrHugdWxiTcgT4u6EModWqhtYWdErIkVdDKInBvo+BntTnVirZD6myqP9xhITcGU
YeuQ5VPJX+u1ynM1ywTTkwiGxDlanN1IP8QJXBsJUFOYN79gSfIMZMpXnl/MocTc
RfwZFnr8wJaAdRGiLQd/USYt9K3oAsBBXPCU9AxnFubieB0a436HAowUeeTdCKT4
bN6ndjKv1BFcv7nfdRRdnOo4PWLxFMdonQOp/pwGkJFx3qNM4OpzkzqV+hxzS3tc
KDuGtSQB7qPdBP3m0efFyCvXDg0LyS6Fugf/b6w1IrpXOeVlXxIUzS5mMXSFrb57
qDJLFXPTco9zM+G+t+PfNCOvsQcT8cPBuidRmlhul3Q5UIRWAnUHm/IRPP6xSbPz
dHRH5pHzcjMxglVFvPmbbUxhxQtLS1NGhR3NBKzQ25ROSccyxNn3v0W1z/y2Mx/N
KT9YKM0D+dEDn9KM5HJ+/31f6SHYcASrMLbwtuVTr1pE9yxOd5xJrSoKrfi2KtLD
5DLH2hpfiRpHNOi/nCRjCas9EgtTOMojTj1WEme9WuM07b+l6yM+g0qdNb0OWkEm
cYbDUOitl7TI0fr6eR7YC0hnZ84I2DV+3NX1yLop4yCd2kKNfmqQdL3AQwznIouy
UegUnNHouZGd6b5rVV3CjMfUCbJWL8Ks0YO1anuA5qwN80Z6Bn4Gozo6+uTimKZG
M7mqDnoh7WjcNuLwL8HbUi/6X04I4bQx+SXQwNRM036v83LXOsmvaLrcTZnX0M8L
2+CWbEbbYCFropnQUwRBdawPPa1qHgDRVSBLk5IpxcuJzuI3/VcLkK19cnr03bF2
CpZeZSjZGZ4d26J9m8v1AVMykUgXV67kz8C4dFwngqX5sxW0WTImisijZG6wBb1K
3ryIx3DfsZZN2tboDTbSaTytvzzU1yF9s5ihazDuavDJRD3vU3uYBxpuTqwGeqze
sriF99Oiy/Hgfy7B0/XKn2fLwVSZjhQkAl4WOl//r9KejxvsOGpuYYXzwum5v7WZ
ImT2xJgaipdpgKQuCwW/s7VZ3ehChh/VkCj9t2xn3eRI9X714U9KOI5VmwBWK73I
Cx64+owJZs4ER5/WDTRhEmW0R8o3ZXvHkz1ku+2t7Fs3t4YgM8LLdV/Fzed1Jonl
8Zm3MgMEp6bBi/AOc5/ZBddn2b6F823KaO8vV7nLFSz6IgvUI7LpHt1M4nishTHT
a4Ex6vkP76KZcqj898GZl7FJYLLLrwSwLZ6530xvATWpll4nKLB7kWgcPHd3ic0r
E/jZ8PzitMS0XRPHchKSurAD1vwruY6Nq7GoiaruTuoMsJpbLCXzk4lw6Kt9bjrA
zyf0D739zqYZQE34L/n0quQVfwcobjEsHR7hiba4b4iCunZT7EN6ku3EIbdGXo2E
75jN6cgsRZmmaG+hsekmrnjkZ/j6RaTlrZLOWZCLd3MZbxRYuYcOLwfs61LK9O0a
mkDmErWRY8HBXatfDcIBiHplR+XDYv3QBh9JFfLhh32hgXr7d72lmhPY6ddbdLgW
+ERL7Rp0fbu5mbeixP078EpdNRWILeshVUY8sEV1OzBzAxPiHba5rNpzPDMmE5UK
mUtBJFl+olOeFsP2jrLACPE/RuQ2php4dCvZIJoKwmejlw7DPGOmJpxc2aUUhF0y
F7R76Ul/+M7S5axIgcAZwk9cw7V8IkhOh8WJWwdQHM0/UteENTp+4O9RufLAUps7
asm4Zb8dewcbKm+x3zHR3waVWOq+51MmB0+Pe+EPHu9VKpOWcD9Wk2nLzcW7Ov+L
AOQ7DwzTNEzLkRcn/gWODicrWyqFusSSqyma5sYvZGRcocSmcALydHav27O34RxR
CtpJIO9qJgsByB2WoVW2iMSdlRPO58ep2zIGYfPxUDZR/mqxBrNTOZNn8BVXuv4G
DfVM0olZubmBh1RVAYdMmNAu4izaikK8BcQuiisjy7uUx8swfUeSYtJXse1jpvnO
t1T/M3fc7rfvjsi/IJGcvwU6QU7hwX8tnxBLt3TYo4XaZaTpgi/6c0Yx/0VJT15e
xtetXBQayT6j4yQnY6jmTJ5F2HmC5b0qmwdVNNH6D5h1FizUn5MBOnGO4givitkd
vTuQse3Ae2pNQpCHs6+0PD9eRWIFWKXG70rG6VupXSip/wXoNq/Y2ne/kFKQo53n
FCpbWuPiVBkkfwmqqzFobb6LwjDJtgvZJbPPxpNMjHj2t7hGbERjtn2ULWZrZ0nC
mxRgghv2xn247MPXfEni4cs6VZwRF8fHn6fTviFW+Tl8wwYPdhzaiRn6BxIye7Qt
ApEpiZvQZ1sb9IhnPfDw3fc+ZeKFokD3CS8718Zd2a402DPsw6Dlsx+hVzyLNiCf
0UHpyCJFlgxhKBXXtThwFBB4UWafoo/yfzTotZ34pOIqGrotPlbEOOWN4GngBhVb
pBVFvVZ/Q9J6WiBpwbWkOkfyO8ctXRkBwJDammRxuPOJbnrlab7KOoDIb2mfXNDi
GuE2WQoC8ibuPOTkGPS2qJl8TeDzUJjlhxQCfw/QPMaDQZv7D8YeEc3zCNlIP3G2
ERu1xR1ojGLiQGXlLjFd4P9fRbzjHIfKWLudw2lfUhsK570PbAkZiyRlBY5mGTFH
Qpq724UCdYOOPAWhuy68Xnl+xYxdPwbdBFEc+xBD2j9Ea4F446hbv5bZNqsc+7ML
OpGFNvYBG7C1BF4vNSfjLR3jBsIrM5unNwb1wMngZwa7JJEpnkkoZjIEELkxCHgK
ySfN0dg1yoccbMRLA21zbp+clWTO1SZnvXBHrShrcFEBZBDhDGePNeI9E5q+Gc41
X6gjwtsuEddeNMi++z0vcW/zFqy3om/pBbqJ+UteHCAgq/XYeckinDnE8Ua5V8yX
9ezvctm9Gzs6Bo0UW7jNM5GBXx5QnR17dFNc3XGj5WoztG96qhHwDwcxsq8Rc9Hu
jIgXjAT7bR36r3Xbh78IVaqDH/34Bhe+34+I7UY6mKskLF8AtW7nKpc/m42EY3e7
NF7bXWMUgKmIKlf4IZ2yK+nTYmDJfRsTORhyfwbkiZQW6n6IntudUfZtZayz+PKz
WHd2i5JmH+QyjvKNTCyH4yysJoAZ9xGRf+cj75go5N9BUIx8XJYQCE3IcnOML3Ev
j90XpcZqKz6ZHxKeuPh/T/sIleuImaiGNMyj/b65QaFhVnR0t/G3qz0Ie302OrRp
JtFRoKo/5M9ax/TZypQD9H9UZFxKzKZFFKBF7Fva8BXNOniB9tcrIJJ3kn52TLAn
+yxxYO5ZTs00wv5jsOi7m2wKUc7a0yPUlC3hbKdINz2645RckugZplf+jgsbJ2yU
ElNkUE9+3j31DAU5LV1SHqcO2nl7IB8CFLgUoAlH9pYwCs0Zr2sPE0UvWfVWerOn
hU4m7H67OlgAygQ6llzFXRzqHBJ96J+keBUyJ6n2kq5F6G817YQcOwkdn/P9iq/K
SQ9XuKV/hxrdz1ZYLKR4eLSM9+SkT/yfUJB+AZ5FK6pDvkGrsjQNtYuSzQemGFQ/
0Gr8YEORQgKx+2dIwzRZvlPNmqj+A0A2QZgY2PsUFwBQJCY9RhZRq8uy9sNhPDg/
UYDEEOygYXSivTt7+TY4R05RREmo4SCtTXtF45ls4PSzcGckvJfo3O4cGBfoKoSM
Jc5Dyq6gW0zDRWru7A5fQA25RxQ9veNoU6tXjsmGB4Dn2gB9zGyws4VjkzwGXlGG
k+jdtbUXekvp3ticoeSVmj5SXukAfLto4IDmZ20Tnjl92gMKFG85WhPhGGriPzaF
1StB6rirutWKpXMb48wqPUOOVNvjqsPkFSScXl50S6OizeDgD3iK+p9iq31ZkGlw
vLTTG6UpIQapCaYfkrknyD6jxtJ+jIkSyXIn/qMrf/E7UgA+VZWHeUBjk4dEUFmZ
1tkuqBzWlVxB/MEbfTn1yGHIzwjF148Z5QbwFBgcy4zjsCaIA9bou5/lo4pPMV0V
pCANc9Z+PzX6BTBrFbNTnsrLHfIXp5ycoio+ayKCQPNBVZSZRLUl/mHL2QIuB5v6
4cKK34oRtJYpVG/LGQI//UDlYZSk7TKqV7ECi9K/Xpo9/k/p9L2r4LsLj1EJsxN1
KFAAdW4tEBZJUjTgwdsRWHQWiL1A6tNJRqgz6M4UVBBvDJ/gZKNo/gsUZQGx3Pis
LgKQDX5t//effRcS0JTr5zqc6oai/TnQ7x0XTthACibbNyMcOWgRbSRoPx7KB2e0
vtfDaHAF+isEOeTFR+eG5+bs9AeVSTO9iLJg7SelMcLlJzDaUf2BzBs8p5Yk43mA
TfompQEiPK+pTCruq+dz8gQm1Zn8XrFG1f6Eio29n75SFU5qFljysK9HvVP8GSE7
w8KQ3VBvELoKr+irvFgZOZH3FXVuqLjIUt0wBNZ5eWpfyNWnHdv+qUF3SRw526et
40Z8dCmdL4qPkk3B7alK0ZlmjG38dz/ye7vtj6hjslWfrkpsrMCRGHTTb+QkkHU6
8Qd4o+wb0SJ8FM9W1nOX63wtlXByq64kolKvQNAujoFfq+cJKN15T9CJhjkFKzxM
KccOkV4/9Yrtpmc5aWCkQSOucX4fjKVmUREi0ZvZDV+AeYwuh6wFoje5wN5eJPcm
c0QMkCcAjK6Up8ym1qNoufwEU5L9aODRDfZaZwSKR+g9R4FrKH1/Rjrq8plW8oZ+
CClldJzCjjmGjcWyt7Zy3MZTi1wWrofk98N0ivYfxysNUzTK+06nX+B8opYoAUcs
V8xNrsG/7QQJ0JuBJ7xU5ETDXB9v8/nl7Wtv+tdZH4fzjuKfBKukveFXalh/Jd0d
RjiXj7VfBsrC5uAKVjH0lzlnRhkKLFKYW5jRBbwYVprgQD8JiUx2YeNP41tFGB9s
NXsU2BAwTvdP2CGC04wYs1Y6QSR42ZV3dAN1FWdk8FKTXXXT84SXXAamOqqTCd89
NFmX3RhYqR/B35rmIujUmnjwWvVYg8LLi0gdiy3STv7gFT6mBG3/exnd4bFyhVqL
/ZBzBPVHOj643efu8/GeL7+sQISbGNkWocZCdTb5ZDzBYK08jtfbGh7QI1R9hqZ+
q0NNcHn+UPp7GDa1vWnhjMMn5lbIwUcDMOC04OcjHnijCQtgPtkqIAK1JySjHcpp
xFHp2oRhPo7ggEFYkYEXvh7LmYrcZb7zzn+J6scp1DQWrPrtnpq4Pa8yEWwwsjyz
evlpf84S7OzGCPhZP2xoIa8/hcUAm/QmSAmbH800NLz6Yaz/+6XDHof5fAoMJBto
v2Uxio5Ux4HWe9G7MxVGAoWL5c3LxBRx/+FCI8+XGLM8r5Ilt55wW00uJt15M6G/
yJoKybYTSW7tGIpFWZOb3nENZcICmh+9GABmt2esiosLIDUvBzttytA4uKpvRCaV
qQaP0xep422Ejt2LYUGLG0U+zrmcVusMJwt1AbLcdVaveQdzsqDIKCNcDcok8kbA
03N+jBEb7maYLJTRKj1CcNg4fvoGAIAAczp96bIJ8bJu+59fH3SFoAY/89xgibeV
qUR6v/bXtLKougxPyHlpAFGYsNhPJIDMl7AYaT+myP/C5aFsE80f8N54AhYmV6SR
cR5SP5yCusm8Mk3nS/Qgdg5KrjGocd4JWBUaRhfFRl8pxaJ47VeMaYram8Ifgdpf
FfPVg3asoEPhi5Vn0JCuTCe/X8Um0Pz66rE9+MXFujLaxaOCDXbyMj+ozAW+jxB2
I38Da5QCiOxB3+ZgFJ+13hnirqA7RkLm4BzCICD8mlghKqvhKLoz5sOTPnoYibYc
ZwCLCSrOpjIsZg37Gpc/7x5TMGWtxH8pUFdHe+TwyLLdPtJWdSxZqVmaDGWedEBc
6TSSvI16mFJnEglE/nBEdK60iDEkyVecbp5wb/K7jq0uB79rE0lgfIxPFGQe9C/x
JN6CLhvK67VT729HQWPp7g/N1tf1q6h6v7n9Iz9MB1GWUHrLQLZeALN/UXScKDv9
8FMBtOMsBVj9JHntv8gS2MZ1yoQheZxp1e/yPHCqvu200ExmKL5mCWGSLUHBrRc3
kd7h12+75KTJunBCEVOCEFxCNeQnWNWNd+LTdFpb00Zj4TvIVBofMTMj1sHAoCou
Pw7xwHhIDUVRhrJ7nUnZ79QPKofYsRzRfzsknqMDnnWCgn9I891pV8s0K6RbirDb
p7VcICdfC7UuN/6os4fbFqsjb7x/QxX2KIbZj/+pq2QQtqYUNl2N0ZpZUCAhe7wr
uQYrcjys8FpSfb8IQq/gkxkPXk3mDJNJwwDKuFpgzaknMLixIoqpNosqBwREMjF9
4hR5sf/tyJdwL4HY/0yHbwsu1xjeRFuISXCOTuYF0EM+JzorClfQH6JLzgPBMuuR
KWUmP3MEgc7+xNk1Ln+YJzWC158lhI13HRx7C1L8QhjQGZPWuzH57VCtdDBzpwBh
3LLVkWW3Qg9gh2/zE0mhkopaYbZlgU2zm1JDDE8uiZbmXPlb7dikLh/2RNbToIVx
XxdOcqri7tQDJOeyJVb5c+ikTsZOmVCJ06I+mbkxtiP3ZKCAH+8UJmMeMJRzh5JN
0l6hB+LFpRzCIxpTTOO0WVDeZ+l54xLUZjHzF76/bjAheCgext5Z/id7UkSKED8+
oqYJGzq7ftcOvgE/P3MyrcNeAVRtMM1F+gJM390M8L37idAtD3icvOsQ5bCM3OEK
2qnt3dYWnlHY7XUwmjuL/acreLaEAjxV4R2Nj2NqRWaaMuMduV65s7jNprcjPU7T
2epl4bfchcNQtpUUWbKkYWngluOI4liCkDG2y9hrECx766chTVnokEri2ZmlFNeu
is5v6LiRGeCuwJu+FghD3tSfhzaVLEvQkH5PViPT6wScaQeNpEu08Auk51LTHi4+
eW1xX2u8kUtNdlGjBYWk46sqlBK/RkoOV+v8OiPEm4nvx/KacxQbQohJU2IM+G6X
CTSbAVA2EInPBjIkHxN7T49ZnOEQ/Nl8ETiR/JLY8GS82yR3SCn9DL9++mHXQrmp
QWK2BNF4MgPvmjqI1BmmrN2zSiJ1GeYAjrbryOkngTZIX/jzOfR5+CjrmbPwFNQw
Ym5nwO45oboKmZRMG9EcqqYTrjTdosrvPB8Nc3cp+4FFoagoYlU15HPuxTnAA4/y
rDVV98MT9jmt3cepUsmJR7U27CcreCkigvybokhOrCQo9e2UtTzgp7om3HdXHCj7
dCyQVwelPAdlAjAF4wUgCvP4Y9TiX8lT4Vql+fwmdncHDQIWZWqqWsHYbkaG/Tlz
ytLttswiMr6b/HICXpe2+qLcXai6Ap/BsVXwAsxXi27BhQRMO0Q/W5QmowgIdjBa
f9PdIIB10p1VKDPHcrksBgqqTfMsdAwLVftYR4BLokgiBp9ebT1+URpWrrsBpYmG
kk4bnfplddne6cz/gf8m1gi6mercdGlsokLv//HmnETU5rSoMSLk7PFyfLw8OQcU
D46SO4uf86UoNl48y196rsldDlx0AxRX4KWrFytF7TdW9RdSdNYKTuxJ71UVzl8E
yl1nKTkPLEWFo2xo+EdC9FF1xAivFJue1R7ufp/EP2dUvnyKejbJj8pXOKMQshAn
v0EWEBGbtJDSlFJPyZy2Z5+scWUj5j1J3UqzDmTZUp7nfnxHEJnvh2dGM7HBxLuY
J+pyYntjmeEzxIYMJZna6yfrLu2wJnMYJD1LSnUWB1gq9tDaNgXIG+umNBZAQAkt
x1S2g/VyyBVPbHbNY6G4usdNe83Yl4xj6Q5nEuiNpOZn1Y+bTjLsUUYK8YLWIO+G
7yLh+mS53r6GTeKA+Sj+/C74i/Z5juyh97iyXwjNXdGKbq7cgmWIYTifOytEYThg
WnmcFfGgOsgI7AE39Dx5yqJ9zs9MF5NkaHlCA9nMp0zLKWZ1CTHucw7ewdRhJYXF
Ld29fO/zokZpDlQqL3dF+WFjiUCAvXjijz89XhZv22UGYPQxgULmjFhHbxqF0wqU
pc2quLXA0Mdp/56YlnpS1wbniixivGOKtA2LLGcUmqF19KBFIuhveZFx1O5oq1P7
PT85lUHjc+Hucy9mCXQMJEV/3hejN6LxF4BGlkEvVaRIOG4OZMZX2gtfpcc/qYSm
QNr078Uxuo5xh5J5VuLXjJfVFunzUPxW5x1hKUkl6g+fPmuQ/ddkKdu64ABf4/k8
XV6nnHNVrRqvAubG/En229WDKIfE0cDHAJZRVanvzoi+z4WN5EpB59nsAg39k1BL
ApMY6mcE/Xm3ILO/QAGZ3ZZ8l9jVKDu+xvGoH7FO34yuWC6hmwiizSm0jXeNu8gx
9+srFDBb5Z+gUcPFQagjSNVM3YycH66PLsfR3KQbZvtPV77gGB7TPeBi0O+oufPD
UPM0xDGFM0Rr9rJrhbJBziHhtHfV2DlLzmKm6wk3FY8mZY+m9b2py47raP5VZljR
Wp7wyhZpmKFB0RK/dBwAe7d7JL2r8c5lfdTFl7a29Jmm5N/7d+XkQjVV7Qrbnjw2
IIMZaLP64F/l/tO2wwbrT1nQgGnfGX5hCv0OJm/VFGhPiodoqBpq6G1V1aXcOeHV
2DIsoty4aoXBZtZEn3nswiZWxY5Bj/NJ4DtQx9WnwXsnC668NslSBQu9t3ntdKmD
CrvkImnNy2U9leG3fxhlKiCbN6YlfxRPjDNW3I9MH7xTxCemELz1j1wAy/7N+wFk
EodS0vOghNHu17LtjKkNCem6aXkrKuB3JL6xVdG9joOADfWrSK++/g1lSAAk0wj+
FZyqfIKiU0dkIdqHhqGUXmPafHAYxngsLdIm1XTZtfmXU3555GISJkUWvUrVnmbQ
DHyN9Oc4uvxKAxLpC19v2G+Gw36XmCSXZFcNS7bwK3wTuHdMvDGCk9hKI0G2h+bk
lDwaleAIJ+GNlZjQw00q5LRh++QUlF4XtaF7YaivzUTH0UdTicRfDu5n/TQ6QY8G
3hRjKiCGshXsJVFGozGw0NrPsKrtt8fxrv/CJYoNBOi2oD1niNoeqFlnVlyjTmlC
eskIa7xkg6AB8Wc6AfIotBlTqveh+79HcAK2dgs9QRN8cEf46BXpYIRKWB9sDk0W
sGs+pBKUT27Kf8msZ7AkzYi7GpwS6kUtKZ6bE33o5+EDn3tdKOLuSpZl+sVzy7y/
4+rAV6FFKWAKELOsGt8G09whWw9XDasF5StGhUHGXoGm0XjAHe92vuxTEl4H60ph
Be0vUD7bFstGsgHZ3/f1eAKO6rGfKakeeMQeGtnXjNI3p6oiT4AmscHN9GYRE6Sy
yh4QDpEYJnfDyRwnjymodadOw/M5h15wOoUDMAICvmneK+FKAjmjM5EhPwytg+PQ
zc+QFTTzM3N1vK5kC/LuGjNbgHVFge9fe7a9mV2XvxHynph+5J5t8RX03PcDxqUr
tZl/PQRZaXGpkJiLuNfWTrtvk5C5npJ8qxBCg3/RsPP0B2XZxzhOBg4WiDc2tLxR
h111u6sbth1LN2BEk1Tnd7VRzg1y9MoHlYm4ZJJJRLEVHofjCcazRh5KcOLeR61L
UHnMMamMOz39wj0Bjk1ZJhFsF6gnwuuAjyiJi9xZKAwq+1XRLr9ekte3DJcwW+UK
RvNjvJQevslgvSWvk0ATrIa+Lx5AHLUT9vYCu6qHweWSzy1WnSviQ4DdjNi6ZZj5
WDB41Ou/kph8/bHkqiN3iuAjwWmu1FwvFVUL4gL4EbRWbVhc62ys+M7oWR9nNL/y
qObVa5giGnv85U8fuST5te9wLmfQQ8qxAPhKO02nJj6jJ8iiYf20Q/JgYpk0Bz42
CJIAOXbn98cSPoERIsTV75LQ99X6xbNdwSpTu++vmDwvvu3DsbFyCtxQ3mQE+391
JvdkJ+uatSEXAkRHKj7zFFoM+5457/zxlOdJo9pjgzZerEzuMYO8P2Qvg9/RTH1L
fFYYkKjYiKxrTzqZ33SyE7YayQD+OtARdRWAeKnbJUMpXNKSWXFnX6Mox0hJt+Gm
+LvrKHWUEzn1giDYed75reOzW8weOKcaKYu30R98tQxeWPDNV0oqGtMKk6D9xUjR
ErTBrSM+gOcjSbSc0UU4E/3UxUXKthKQImsPR5gRGzhJUc37wvCJGdYF2QR/UEqa
Nby+X3055IUj9Wdw8iOd3fJY2T25W65SFq7Gge+qywggKULi7FnRa9Lay/6X5KUm
NgRGZeVkL4jOa6PrBWqzfYtTeRFbECLFANnthnmIckX9FpOoZF808UY3phQh4ZPM
xPkYoFF8rdUizo/zHoKRREBubDi5IzY/To1a4mU78qUqcvw/L4EDUedP+ClU5I/I
+gbSrFZHx9VDuayMSJJzh/oRW6a17EwJ8J1IsHZM5d5t/fY83aU1vHtoGzBU0DQR
ExetKH1EO76vUfXqAV+DX0m+hOAWk7Odxmq1uYFIfsD7Fl5KCo+c/146cv+R5fo7
xRBhcuyrWDKrPgp2W44M1HY2grxPkEPGakpjCfqmINk0iM8nkuPN96D82k7TiSYT
KAUNB0iZIUyevU/5UFmUeAA7J9YhY1S2pch+ionpW+K7OsyRJ0c+XPBMp7+LUu2i
4fEk0KzHN8aOJNiw+2m5ZTyqHlB21tWgaxDwq+Hh3tIQupCmmesTiWvQY7PZhiBy
+UX10Yk+fCKBEeAttH1BemUy9C57osoklQw3rKXlcG2vVecY8xYedwil54cUZkDM
Ete173TWZgWn7xtar/TWXKFeVeArHsTFVCI/wz+hbv6u6DC2LBXFZrw/a9Yagu4B
ch1+OpuBRSYTVCfXh+wJpJx1IwTjmSphOejLVvIY/v7P5HxNjqV+B6XnC5Yj3VjW
400oOOoFupGZkaZOMMzSFKqtCAIhW8OS46b75FB99HMg9UBoyTd7H8rlPydL75j6
1aGxmseHboWq1VOHx9Bu1saqkRbFbVzm9vUNZ9IMe0nK2JQze4baAHUAj8I0oKfI
nJ7ywDVNEHREVCNgz1WswZwGPosOq4Bjqsf/MmRHr8Z1O03RGDDqd+gQddu7fq7L
X9B3PfYTyBmBnfth4l5JgoJ0B8fLyAZnfQYYq8jk3YT/t4TpVQgakC6fR+elwR9Q
KQKikHyWX2hS2ha5zpW75F/xPuMa4+KD2c9I/wJQNP5+k5vtsYL/OU0/4YlbXzaS
WfxJ1ZaObakYkqyRsz2nPPqHD3TNTpskLBWeJ3W+S2dNj33RYK9isjZBAbsknRhX
mjmTL+r6MjPM4Jo14sC67IMypNc++H6NTXzDDQRnKF61YjlRffm1+Huqjejk1fc6
7tanbUtH+e5lx9altBuvyk0oLB/P0FuLYWD3GZebtAWXRnCpQqPtY2W4rD0K/8Kw
BT2rVaCNDq2wTKg7Oj/Uxxpzf/sOE0TTXolVj5UCV2fh/wXuAttLV+pk4MP4LEag
YBiOcaicla6Z19OLXlYYMkfd1u/0Ya/SZ68U/rv22XBmpJ4TIPDhZ/z5TZB9bf7O
7tcwCLi/GQr3uFTad8APsD+CZZuCYwat1aCSj807hFfuQYBfZZbvsNi9bE6p22MH
Veght5H9/nheh7+0IOvly2IAGN6p+SPylT0AHMJE5FTXQGMD4DwqLLWaU1mo2JBA
+peenyjIoDtCnwqnuc1IDio621MjOR0Fr0dWK008IGGPXhxhPuiEqqX2ula1clUV
7jjTVsXFONBdIhU1ZODAM53kl9QcbhR9q2AB0qUeYBfD9MPcrYL10jDGKk36wNAO
tT4Hj2tiCrF7Z1nesN/mLmAHlLRXUKl79xfmVuCtv31s73a/SMscM1YMr/SJgyc6
Q0DpeV9IE3Ek+p0pW50nvSpQ5hAIbOdES1Lb2eZ1gmz/ASHEDNGLV2ETDRvTJv1k
YsyDIGImi/MuJY8FY1JXJRw/0twifd7XKy5s5Yc0IaVUx3AjlznhDHDwFCyTUhWa
xjE+LYNVibACocon935qNwFasLK9vXd+mIRov+BGmx+T2bJF48IkxQs75n75KPCK
pEuh3zW7Wy9FBrBo+Ldh8rci/Y0qWFbVTf+OHbJ87hx1ScPMo9xT2J5ODWZLemLw
vPd130I23pmZ6Pyt/bYmzQetUwCE8y5r+OmwudaMZyWE6S2ZFT6yOIvusz0qDawN
MMgzxy2O3LGfaPCT0Npm7F0E6GpzwQYk19MnPjwiUa7UIRnWNMo7YVp4kBJYdnw2
qz+VpzWXz11S9Wxtixs21I2sI/uUH9iDw19y34oVoKMQRc4LxiNCaP4sdelzpgkj
w6WP0aWXIGyKZxJemDzOUwuCYljkBVNGd971FFFQAAy8IvgHl6clItnJuL1J/NuX
xcq7/loIRlpQBYMRs01XcgtKwxIq5FyZa0+QapQgW7+gscznKep7prnLYs4rqgQ+
uonthDzB+9bG1XbbHYlm7bf7Mv6wKEhW5uiCNvXZIX8wY+RwsbplqqOkLnGMJv5P
B6zShZ4uY/8jugkGzjeSTjOfq0bIMUQvgiBYvdmL/xKYiPIWhlr9q2k1WeUv6KBo
1RZJ72eY5cEXNw9nc4+Pgm40eXBWqpZ+wqHXSpp55KRf/fRVRxineVEw1acUNmV4
SY2Iy5HKd5U9ewmOB92GT+lpUkwwC4MkGRPMNNLCbr12urIDznT6vnpNSSkki0XP
FdAmKU0Z2Uzd7y7qMxx3p03x8Q4MISXBUmFKCf4YIkUH/o6tp0sAWMx8CrxDKwzC
U0cdaPx/2ZY2LjMW7ceFa3gYJbFsTohn3S3klfxGjWlubQztWlyNOYynTFM4GoNO
WUaHn4AV1QSSR0Gnqre98ovuIU98XhsRdwVADMAiQA5JDJfo+Fj+yLAf1TGkcD+B
tfR35g8uHf0iOnOabXiz5o6tEJgVIU7xouvHmy51bzSrZdgpNHrbrw/2NZdiEC1j
j7SEBV39Y5zKpgKPECCJjWy2/i5YXdZpcsC/u8Ybczwjwsy9drKj+UyA/AErbeyx
xSUeS026LdKexbRK3Pi45A0uGjEt0wrIdTGH1NLtAEQg6+uS9hCS5Rjrfnow3xpF
R3NRiSvn0Sstn/5aEMHqhjhxlvbj/tIDjy0VICh966uhOBXz3f2fxvw2MEE1C5uR
/Aqku/dVDq/e6OpmzfKLA7F5faC5db9NaQpz5TV/TQddOM0af8C20LnXp/LL8+/H
AfGMrLOA5yW9+djwY4pDxADny15uPYHY5W5CkALU/BSJg6ltkqNxxDHJTAr0Y6zx
oDYDdA0k4YImbBVAtfzg1nnyD5o57gDAuO/9HFx9zeHs1ub2I93PyX1q6tGxCrjq
74BqXTYlRlG/alCeYibMUeXfmERo5Es96jENAwqwhZFJyP58dK5SkryNrN/m+4oZ
H3VZ42RT45okBg4oSKvo1UqblUXHoFZPj6/4konedvZwGXsu8bpW1OQi2p3Eia7V
IYcVdAuJl1hvXYgwByDZ72u85nnbDtSPOROujqdEZJXL0aJFi00deKOwiMySTaPx
kCu7gpPnk+wXgvsIYASRvgPr7u1BC2EOfPs8ulmKNV3aNnmiuGEQiIzSKCaDeKZt
BizWZM+8vILDeA2Glilv2VZUHT6tTuNoVMCWvPEbFBfwaCPpI7wTMeBJXumWhHuY
6slvsoJmL771nCvWukiE6rebizBIBIhIEi7doblB/2H5s8UyQfFIeYTekV7XumlH
adGjgyRTbrsGWJZcAMHYId1wSFu6th7ZPHrgEhN1w2tGnkO+qrq3Wz8CQfHKCeWQ
CNpfghnED/jwgqe3YJnE0IwfFxNHZUbnJ7hOx8w4Nv8hqq7Lo85ooPYXSULWTuKY
xI811LQELsGEQzqQozTM7j3/RKPVwdj5PQ3O1/Zs08gNafyA2XdLuaST/rqp7+1O
tLY2T8vAwaXA9+SndfewT8HREEEFjDU822OtTvR/v8OgwpmxD2QRgjiHmFLcvrK6
iFnWSUhA38h8Gs4W29angJoaSvr1D9eTExtmqn6Z3sDvMSgaEb53bxTAy9oM3a+G
EUa57Ru03sxACyjf/rYqmC/1dKqgcRTP+SI9TJBe60Moiy11K1PB4RNHjB8WLsha
7czaKXTV3t9nBMlwqmViQhveh1jzEhs/IcOS9yp+yZsZaJPSdNhkAkltQ+4e/BqC
9mNMjMpRiykLgNBrYR1NipwHY7IjqRDTAXPxZ5v3WG2gQKY/oLJ3NRmTrGA2lVAU
MDc9DSlHxVVAjND2TDgQSMTUg4SqCDnMDBgDlyfz67yyqlHd5LWHljQsDOQJXQGD
cqzi1lJ58jGB/wD+57nMharQBOv/n6Nkp2k93fnDfFtmxeyEYBXIZBEvBYhtTAiF
yKfM339+E10pfHpaJOHa8p7NPCCdN1YGWggvV02xXl+QoUEtuJA/D7V0MY4AX2Xn
MuhVWNq1ErTSYcc6zW+Ri4Eu1k+A4UZ4oZpRC1FbS7Iw2YsF/5FJBASokzV6JEzg
9p9QN+95xIQ6DxP5d0IxQwiYjT0OGc0+BNsHKPxiFlT0xDs0hLexhWmZs6fvxslk
+0bA5GJbT9PFRCKZRt4qXkZ/T3lolP+gnSaSrnbHlPWEw5LWZhL18oRPy6ybL3o9
x7Umemovt9V2sQ7BHB0tg4VVgqaMtiVzcVUvnX8T4WtHn9ZKnGYUDZvlwXaXVhF4
l3PY7AlhZHxWE1R1O3ydIIhvyCV5651ViRYB1p5Wi1Zr698pNxzy9+mM8zEJkC0Y
GXXTsLpQEKyh5hBvRS3cgbhPahyvlu4GXMtS8/UkwHUYwkvpAPJRVQkLDu8NHQ/4
oarfsAqEur2CW3k05/VNo17FOVYTiFMUwFuQispIWjmGWq3j+TdSDR6TKSDGPlXu
2RMFp6VdW7xdP6LgPpPxCWx/11jskUExP7Qo7H5gsxreE7GSWnlIanNl55BnnHL9
/NPV+DZ7lMn9F2o4dSXXvPeEzYPthAYDgvA6OMLMOb13aWtDqyNpS52deN1zwQvo
gjN92TDBE5tgZvNAcPnIPwFcYdeqz3+Flaaeibh94W0cLmSr7hbYznv7L6ERzTwb
ws824xmI24vqBZ8Oyb8fkaxNXkhionrhSquRN8fzNM7BLPhcpRBTtBpL2hLuRuCV
iUTRUYndHz1JLZi7KkN/0/HvwON7CbwFg1c7Z+g0rP49D6nwdy616lo9RW+LkeUq
jBn1wJh5M0U0j5hxWcS8ZnOxakUASh4sInzIgmnu2iD6Gtd3+5WfYvwITl3m5Bkk
dQ3KKaT/LM0sUcmYWThmgEyX4frZxCFiWGqYCjCDDqX+T54IR3ihsei86Iy4lqd5
L4DlrqQ4oDMrRJ6/nn+YVcvmJRB7cPHdX+lovitv7Q/GOxoAtDkCelDpVXC3DtGY
um/U1+HlugycUcbJ8BELzKV7vrPDNv2Q5/xheur9yP1J/+4PTM3UcRsQrDChxPO0
991hTwkWeyz7MqAlgTEZo/6cwqLLHa66KtTQQwP8iNz8eW4Y1cZ3x+VtC3CUSlhQ
AEzlvMjKv/XZ7kCbpfvunVB1l/gau4t+Sa1ElokuuOsJNPQQ58+7PpdZx/TiF6cK
JdDHNas3qThcz/SW2PBkEIYBez49o9074+dZvLjjbDp5CLPuOEXJ2dNzrOZauJCL
kcirEFgtPYaVyIi5LhNxDeVSCbSdut1TBdcd0zbS80JRPqGyZtpIjJT8A7Yirnbo
JfJUfcEKRakQqRSzHvFzABiBRv5h3X/r49QiR4S+hCg6RGM6AKr7F4+CdALzrKGW
IwYgl/0vNda+Q5CSlffxMfgXjhEo8r+xoxwdA4WZJ0MUgIunM8YU9QQfj/uemcB1
wZdkHOqHQOob+MGTOc4wA+k8a090aCQI4SJQBJQyem1l5BKcpcB+KiCwxn49ARNI
/M43jYZfrniVF5v9Ty48EWcH3ut9z6L+bKBrv+JA7XQaJqLOoRCT3OWZy7jFZnOB
DNv16illhZLWcZbVZV1jOqIHU7yr7DerHYu/n52Kmb8pAj2mQbGawE9So+E7T02M
dQoI1q7mjng2yhKHxTg9NqMHM5fWwFQvCCV3HSBLrGL5ekbQ+bgUnwWYt7PK943V
qn2YP0vXPjdI44QT5OPOqpSAxUblBD3rstE2/ts0jPUJCO6JK6lDNUCCJ0Za1g/2
g3gJkc2pfO0TYsdEo6hxC6wG2OmfLmdcDPEmz0s9Hq57Ag0m5SRRc9is1g5sjmcB
XG+2RaFnjd7eRPcw8eB3POz01D4fvIhnQIFXwJ++gHoUDbKnPcduFOzSsaNIWnBJ
7CgPX7NYvDSGZth9uvrAVPBQJChfpbyUZRnJUBfW6fjXfM/BV6IiJR0KywqU0aMt
Qn/Mf0N9ZvtrsqVzeQu12DQOTrsY7FwXdTpSSLhCYIUNWUVihgMo9/ANMBB/GFXU
nAxumvgdsjW6TXz3SgFu/Nf180VJaw5zv7el2PueMWXRcejuMf1nhVuBa3EHouox
F1LC+PqRX76t4vUjKyaiEU4uVgZM8xzWtbdRI1OsoRMZHuITWP2hZZpLlKDGDBeO
94J1jVV8ag3jlwHsYJyrAdDxk0/lvjaDlkJXWsURwxNYuI82VRK2i+8wjM1vH5Lm
lYMkkd/gh0U0lELhh1jd3juUkwZ8YR4rwA7d3c1dimWVmBZbVDf42kxzBvvBy3Yc
B7PMDIosfNUuSDJtQcG+riqD3+BdecNv1sVrPZmB9zAcI0en8oIScU2xQeRc4sK+
K+zsPcPPWPJ+9BFpH7YKHcjVsCnLrZGRpChnawcopSzRQolZumaDh+Ox0IIGyFd1
LYTt1e6d0bhiPRUCy0CQLQtGr2HG07vgFX9euyh6q2CRbQLKqG89swy+y7k8iX6p
LT5TXuOcQBaweAGLhmbqtVbTk07ym09nJlkVHkTumN8dj27eQ1wxNUJO5zWX4cMY
/YIGLNoycqi0qT4NR+wiQBR+t4uMTM1mNEOymsekpuby9dD3spgcmvGtwtQe1wJV
kIPddGXdCjb1HAB3Tz7c5cSsuR++XGGiXZfKC/L4/ZdRoPmdtOPng0dcVs8Q0Wg4
TiZd4MjlMwOxcDUTkYewlPbidNibVNrWNT9KQrXnjZkqsNmuRnYVToiuyMD4cytq
xWzr7+JaW1vRLgNkh+QohW1zpvZoWGyH5ZJDxtxU06VLqnmctrLfY7I7qN/sWlsl
PCtCAHaLAZ0cVileVZFCAREDB27Ez42ec7CaTdgDSl5aknQYW+E0JxVngfWAEe5A
HC73P19chzHlcXJiFMuqqw3ALFlWuUkWUnhTfIEUtb0onp0qOJAQ1cEvEIYmb+ZD
o/Dl1N4azDWz7TWYjfySKVHCHAZwFilL5tFnR43kYvjOCEkCowF+ZZKEEvFEZexF
Z8Dcn9L39nNbYX3A0UNUqVpXlVyekYhR2IA27DWUAbPNl9bpGSaGPWq6Q5ifW3kH
1cOauKG16CkLy31Jv52kpPUptBw/mv/LHqFYenUDPwdZ5zlhNi73WEYfKPIhuY3I
pV4hzjYnDtI6+aWc2sNmBAm49a0QyuoM4lx3Xlz0PBzK4LKY9IKm0RRjzksWHNrC
V0/kH6Xv0sXQRwp1AjHcLYhb10ohj66H47iRM/DnFYOqHUP8HnKtwXp2cU75FCd1
YqGlYV8oaF6jKYNL3ihgAIIZWRehcEQ+21Phe/BLJPy34oSbqng9EZ9NSOZvdt6w
aOqm31XUJc9Hl7EVRtg/jaJeBPZBLhmwr/zIuhefmtMCSU9+/Qrim5vCsMzKZ+wa
cd+sS6//+cUPvyhUxdxhI1VEJ4Q0HUO1kSG27ULPJc06L1jh+aWpUvWO81EZvO0r
D8RkJmTF6DD9N8e++NMbd7ODc7dYSsPXIYBgkCjdDQzDeNJGDDdjR12FB/GG8wty
+zBTb4v++uQgB1cH3YqycCgOYCUuQvCQ0l+nJA8DNSG/cbWlwQ01jiX825ET5sZ8
/bL1olNSyWUyQx59LKgJgHzE3c4KXRdIyh32u+gQovm59i/2TWNznv555vbQi2ZV
CKKRxP8V67pyc3948PM6RMOTMJ7x2OZ3kcp63Z2HMAfRLXYKkaXQiq5tIWS9M02p
cDUs2wvjkOt5Rp67/dwI8bY1kEaMGU377t6l/X5ewpWM+e4dMEkWOOTIe3TQEjwh
nZvt5lvVWqJsjsIdtO8fzltE9LmUCgd17iDPln/oSizv8qJYDNa7XxG0hVykfJ6I
UCTetsvuFB43QGuAMCCaxC1Cja+yuMQ3q2fL0n5hyQQoI0RamOeckxUzG7/o5r0X
G11Pi0kGufTcllfmYm3Kd99x7PXfx9+k3fPQENashjdr46zXHX2lvGoOa1VP4yeU
9ac9oOfgkmNdG0XRqnIiUys35IiPBUqflvQ/M5oagJCZSMYHH1JB/sVb5djjiIoB
KkH+8rYRpcsuTv+O7flfeEvW0lGVwUHyKHYnrJDc8ChXYWx1ymcwvTQDLs2eIgtn
RjqmDhvZmYAeJ+QR8C2Mvr+PwupNeQd/nxoYCthBHAGIBM9iSu5FZUH0HvJfK7cW
4dnE/S4qG71ipvFEM338eKjREEDVVvytBecsj0UJ4sPY83lVQDVIlzqB/TElDgW5
OCjf0NOfjuCwQyvPLrfwQGRrNJtSnIgu3YBpcw33ErG5nAudeStOOhkCfzG3XhCc
SMqh7noSoWf4kdcaeYhIYgk6LOegB+c1+6C9fAvGAVdQ0uhAxfwmWgs81iQwrSwG
fC5xuN4Is4KH6ttOcnmtiSAKX9IpjJXXJ/3dcz2IB9daZFrkRd81Y3e2OvCPMqIv
W6e39OOkzaMhpC4yWVhn9FZiaki+up6AGxyzqMFUDPwRVefMq6Q1ukFUN3m3cVM9
1QDtSHAP5AJFVoQR3L9odXVlOxGBfvMfU1jUX7atdG7NevoPsvljpg5f0Ual1ngM
bPseafqjEKeLCJgIW0e79aVODL4Az9uBS91+TW/yiOWoScbijR+WtDkuuBkRTrjv
OpRBf+HySrtvi8IOyF+jk5gao/DRy6Rjwbi2M8GDvmUTvMt+Qht0HAAFllUj/ZPg
rKxCzZYJ9Jipj/PuQvLJvShYBbgL1fnIWVjVz7bVeH6FTvw5/7mGYUeOmHpfyAPI
0fB67lxZbtIqdEhkq/uOeexEUWBTeykz7zxXxuFXyfJW9XU9MGcqWnxleuOuTGP7
+qhkIy0YoupSnU8r1Sl/9yoNN2qvOomkOg9XLFScVWeoRdjvnhmXVi5TxjZF01g4
g4XZHDd5rG2nK1KEHsQAs8twcEaEg/s+aPozcrTb4OLv36pdCHdid7LNfZgT4RhI
0jnn/PzS5+M90oFW+ftuHl+0Ow6xRMy30tdF4Pb206R695lq6V1jSYTAx8zCnWPV
3JyCn0p1k/6Ulx5dQ4osawMCdY/GJDak1BDJtatJn8YWi10DpQgMIs+VRHXZ75dt
iG7a3JAnavIgYb2taz5A4dW4qgOBPOQhzLWefnTJCeGMltFfmmFHiGsBu+Y7ytU7
IoMT08ySqGqxmd00/PlzC7CQicClCiq3NYFGmvmkMNFJN1xRIho12NsIvtgj++0K
hve2laxuQ60VM1waSmR00VxzNizyIgj+WCSaq4NdspRn+nwiP6ARDJp6iWR9f+df
00bScYw6uHWxMzDBPnJht5spN+vCTCHMJoQLn94J19dXyp3Ot+tN5wHGaZ6PxZVe
c0taCudm3/1qVKs2Cv41FFN2wA7akv/MJLYiDU6GST1BnqrVBFwpSvjeFWqwXz0I
/22zoxBsBBz37u6ObxwwtefluXtFeYvEnNDMyW8d07djqODQl71jF/AD7hI9MdpE
On2cD38+8ZlXVszcKRc1IGfEe2Fj32VhwdX1w8rVbBg0T8GZ4P8RPYKkniNA1wgS
a7IsQyzE152ue2SQOPDMhsCe9VAiVgMSZFfxhsUlMjVgfOjsyhsFOi8TUg1JwFWQ
tgVMNE5sgYB+lKaq/l1BgX8lVqDnXxWrwzdzp0SrurIe+TZuOaWi278fG9Jq0y+k
tjUwTFhG5dm5nwxhvjT8pzcp+EsFl/Z/YlXwKIPZccep/YtBoyUn/9MqfYxnUzvt
15c1eG5E3514An2L7riKqtY7cafGNf/qdSmBTiyZfJ6DzBnVw/aLqIzfqlYtGYiH
7qkOyB7BeW3fVq3maMpm9nQz33/7vVNuns1YJ18mLj+e+EsktNvo0IjbAPvkyMIb
ICVmK+Axz+8ThpNeWVkjSPzSNEdxBqwRiZF+0OBxXRMLyKvp7sJFzyvs24jHJixe
RCnN3ceT/fYpl56IH9Pz+D410FA+kgFLw7NYo4GPrPylQ/A9qY4e1VrgFt3WcvHX
AG1AvVxuzJUmHx5Cdt9CEsK7N9QevxTfDAzKdo35arViQCMh2GEKsLsO87V0kX5i
2JzquFVbWIA9ngQzmnh6dshqd4UbFXJziz814SIGEJDdr+c0QzE2Wc/X9Rh+ysDc
3p86Efs24GBYzl5TBgFW98u/oD9upEp5wzdDc0nKGd7bjysqjemXZJ0IYVVRD4R0
r/EIePeznBjASLNiqU9AUQ7Ou0sLNBr12kkWnogi2/IzCrb8ciy4t304r7tF1fbk
q9SHXVi/94SSTwekjp3WnGBJ++yZoRTIiMAlhaOx5Yhr9Ui5leU+NKs1X2PbaQPX
RsHfrKK9qCTXL3iBKw1h0Yr12OOQIxYRFDDuBs5OG06NKXhiNVL4WuZjznRoHjSe
Oqg2ZSJekA0fyDHwfo6ayOlh1vBkX9yvVG2PkvLD8U7U1+YW599MmZsQwuup+sH7
T38vr907JJSfquDD8BN+ZyI07SbxKfOTkbW5xLzoGkFsOzinf1u3al1giK0SHGLZ
I+G5htnZrBbvh9EYw463vrD1cG6MJ46J1KRIzp8tW3/0m5e96Hxmv2FfT8LtUp2p
XtdKmLxdoy0wRpL/a9Jv6yj/lgxZAzFM/ZbViIR5DjenI+1yXLb80dL3mQmPLp0u
FN6yKpha0K1Vor/lkkpQhnzKBwUGA0NB8531waOkvJimb2Mf0RBcG49kjDDITmO5
L9CgTCWefSf82Z4+/nwoFC1C80vpvOXlWUvLL+iBO7GnX7uLRlPVat9UAzziTVyw
a2hWsuT+O9mQ6z/015S4BU1GV7G6Ah8UHwQEcoeYwvxYSnwfFLedh33iV9Z4ljWr
2HOv5uE2ErH6nWGLrCbJCBb+xPgioTP01qpNGWYzTwsIubrnRJHAp4XCX1SEB0zp
pyQwlRlE6b1RxTbqhkAUo7XJlkQVHnCmrDLALmqcYE0lfYRQoqwnvwMNyw0h367E
yIaiP6hVmOtkAtCnZnhIWQ0aKNLrrNfJSG61BsTHjWf4QI4LRz/sGKnaPQE3BK9v
1Da8ketgjHl+nhGXbQ9wUrAZCThU6hPxKb5N4nggQoYz0lO4H3c1Wi/UOTSN/05Z
maB93Z5m7KoZr1kbnYgI+Ix4OVE0TKufDVDPbgp/Pj4cIXAL/S4v+X/FPRpvBwRD
x5TjJUaSKcP1NJswy2CADQQjxUr7Fno1BamOjcSmfp9JhKHImy4JVTO36Nn7D+tX
bAIhXztFwkROjiY/DiMP7+RLMWXOXFlDgc7/H4lxgsYckteigLDhjLMlnSChffI2
3iF47YxAY8BVuCtglh9RkagCwQWzU/VhwYuGr8omqsb/zV8Q02AZ+YEIFmOMcTd9
JHYFuOwcssFkEx0c7pZkEd4SYfq4GdRJKuzEO03/6SFiwfjGegMfkFrVHEdQ+xZy
5Z0+yGbJT9xLvki8VJFankz8Zg1oaO+ZRKgxcDdGDy2WVRrFUOimjvQ7mtBc6P21
zwpvAYnCRI3obx7M1M74Q+W0c1D9emqkIZepWzi/PFHlpW18Pr+XflTjiLCxBrzS
hrQgvpPZuP6jCcDSn/fqqIeRPIczNcMulDGzptU8c1wMM0d2Fxdw5GcZ6g1m2Iap
Grtn4s7jN1kiUvOQNr5wSgH2Xl8oOxMK9+i/4kBIoZcygyrPvMj7Mm34c5sPomGI
Y7zD7GmE1TwQPoZQvEnOMyHswuiQsZsWK5k5/Pu1/DrcEyRdC9Rp1c2AnzH0+sxv
kMNF4EaPqhO0FaUJkrXaIre3rTlytKAFwcT6JIl6tv+1doOhNbfnH3j1946TAS6d
1ng56IqJdDT0KYQyjuldYCFt3ej+0jAozpVGH5IRfVabKHf+bO6hYnUawmS2qFRJ
RxhiHQ9e46qyvBFkYezbyXPKrmpFMlHDGOSvzjZDsgUHvDIv/m+e9anNyqlGd85C
E9q8kbjo1M9eoJornrNAslG9vOkNNBCrHzyTkRu1q2w+FwqzJjOVnsxqkqUzy8io
WHYq8TI4AEoJ2N1Qt0BwlDDdZPdXjJqI05rWuZpBycgTRWIrAJaXqcHcjcYuwli0
5zZXicRI71wPgvHcZYV6FivbwsAE5gu0kB0aXYfmmSKoIBxucMgtigWU5Wqb0NHO
XjgH+2G92oYDyOjTPP2Nl19yigF9mBOUpyBJcRSdjICnJ422/gTix3UTP16WeXFS
swRBpzJLMORQxloTVyBO71dL8KK3O3YeDJDQikK9PCIAHDmBFb8pfQibIXHWNC56
XJeKqv9uXj43KTnXH+NQDb8BVpJga7JGnICzBi592MkO4tMMHuz86KiXdgkpBf8/
TSJZOuIaawFsNcbfrfa9aBtBoQ90FFoiuPD0QageYRDCQGkjDoloqN9RHEIiLdWr
oS128KYhrL646KrnBvN8jIs68/NnprGgTC7TZizPwOOnk/Ydvh7IURxjQ2sq3AAS
nNYL9Pf4OJKqnWUzgtYS2rt6ZVSvbal6K/OC1o9oGyWhVOm06lAQ41X6st8cZ3aZ
xstgYUZ6ce7sBaESOT4Mf3xVwFD6m5JjY5QU636RWa7iZszlpS7jMGtZnku0fho9
e/cbzPbqzL+ve5hZrnUQ9ukhZD8kTAE0cVua6i1O9Dzu7l9bIcb981uamlyRCXdZ
jDAMMEq8mVhdaY2/sK4+++6M+NkLqzl7kHwifhWVxZqn68LQ31w+YdQb6vXRNVW7
jBPwBlfFQs695AP26guOwueQ+ISv6EU/fn/wkCRLemQRhqloSVPLnZcJiwjWD1GS
/JXYwnRc8yPwzNaG3gg4sSXnpIvTakwZIturBwvO1JwE4gyStR4Ms5iBU9qGdFWT
ZQ2I3hB5i45D10oW9p/PwZCKgAX7fd7CgtHPu29zJBSVQE4fDY3mZ59B4R5QIISB
9putngcyQTmMdO7SDe8pNhgw2LXZzCRN5RXiMHzLMyRC0q3+NOjCtLrVOjxqzwRI
iV66vSHGMr5ICq43ROxAmKEdDHRtiFMJv28bG5eR777koybOswGHjIKuTOf1itHX
FoqRE348ZpMYIhywGj/MvmPwhB2zjpmaLEeTQnMu/66zvj9y5/CYb9/JVxWXEY+V
jzLgQnnez83t5k8uz7csKCYj4MQUnx/EgyUv4crtqoId2WYEOSZWKPUzyXXmI59g
O8HYxmyB49A28EQTbacXCz4dhLy6GXpduBWDY6pfBJjWz2wEBasJXslEenQhu9D8
Hct+F/S6VLWGHYz5Mdua+FCIjd7ymT1/wj9ITz9SnkiKbzvMHH14lpPhXgRP/VD/
FdiepGqBgnc1/iM0BJDfy+nkE9ZMzG9CqBGJ3iZ2+dFD6dePZWQHw3JPDmAyGRTm
WYtBWoVafwkrolbK896G2R+Rpi6wDQCKiU2nK5A0gZGM11pRS4dpao8m8C0s/47q
aTN6HJXA+q5zILRK+80iQthQZCYb3XzB7PcxYOagxLF6FsMZLOch8/llJvQcyY0N
taB2JR/SUGe2U0vjROnysuCputLOWS2K/5Jj0JEJ7kuDTG2xOOkfdokVbLfgvawL
Ie02Jo+lbgRCBitSeMdJelHwWlL7nLtIxx4h9zl+mQn04JirC/DbOwdMSoCfHYmn
geOUfcz5Ep3Sip8mKey7ImA9fussjqqyom93+SQhNX7uoLnR8DPuDhBfjWZ19WQz
YQLrO4/cOhePakWDRlniVL72CvrrQgfTDasme24QUpQjMXY4MrBoOsMl90Rtl/n6
g2wn+5pNorHQ7iez3f63TaLWzQCZ2QJyveCeqC687N2Uq+0JFD/k6GPWx+47JsDZ
qI40dmQuk+gKZh7bf+dB0Ucm78/1JztkvUAjkrmKxMPMlw7WcIN3XO6V0EEMku+D
UZmn9HgmhzWBR0yDdcLZaF4VzcPh3Rjlq0f1ov5jDh3CsBqKFL56lG6uGXbXgZJ4
lquuEUvcKQBQpde3REbDAkv4jkud1PWhlOkxFNbdASaJWYkN3t3LKvvuZgr8b8I2
aFHf2lsSleyPxwWpxkFK5PYRidqlFu0knsGP/v5+4G3bg8av6nPUCqFAgQC48aD9
ht9UBhl2+AjqnAizwGLIraJI8YQHRwweGUR+NDdn9EmkDKgWDJEE45YtpIhhkXIN
/R4g7T2STfe7g21B2rpfL/AtCEkCRnjDm9STE1pQntt+D+VMrU3cOunJtVDkzm45
7K/adghxj9pJ899ogC/QIiiqNfxARaegdr1vByZgODZy530YAeGUPna0umYZJ599
2aMisxTiQYCK7NlYgYyqFWZp+cDFnSzjFrkzXptyVlZxg9Tmf3KM6pDvC5fXAy8X
ahCULtuX6tuebYXb6blAsKDvQXnHJXs4qT2WNbSlh1AO/OIx4N/k5gx3ks6wAI3F
f9k6s1lz1/tInIcmTsjOp7ap941sfWjHi5VcF/LJmCKU0WVSHfWllbc0deGMrvgj
pb7O8cbuPm/MDQ0S6qBRn061khCPZElAQAq6zXDwzfcwyOSRm8NFL3mLAQIX1Ati
PEVBHvKhEshzzxkFGu8UcxfLW244O6xwTdWAjJlqz0MBa4s2vzIlYseiCoXHJ2i5
kmzoUCju9/9z8CslpF3jKTCIOy3/4vkizLx5ScdMSDHdvCCA+rq8mTSkmHI7lm7G
qSDwDwS2F8V2TQ8cR8zmp858GJ+s6dWCMNmV0kbbIjGtQ4x8zELjWWrg7hoIH5nq
0c+SufeWAaYOn3kwLBe9XebCqQwqCdoIclJX9hOY3Ww5HkgtPezN1JJqwEDZ4YcC
ROsXA8Z2jW6j7HIKkzh5Md+QVGwsFWB9l5hawVAw7IzqR9ClT+uv5NlhL4d2M+CR
D87SzS6kT+0VdjNifC3js13B15rXXc0aMBjT2Y1TL8ZUCKm/Eg3JbDDSZJvVjDi/
k2qBK5+9AykpUtDKrdo2vqtbXF/nhX0GPw1qHMsTjWUka7tnStzvSR8nsTG/YNhR
7lVG/PriH+A6s0hh5d8hNe/OYJeOJUUhAP1duiO90zPkcuu0R7TVBxVDWek2+BbI
XM2nZjz360FbJ/jNDBSeugo6UAgIIj3ua5F2LLw0+ZvrnU5cZmFUqIBSwBCnR9Fb
7Qf8Lap3gHED1HrbCKg2CgLaJG0uosEQdGMQh9JrZ0BKqUUemrbg6mPoPpBHVXN0
Z2E8BGxIIt4616Zmt0TD3GKzZHQmyBOnbWLJgxbt9Q4U8cd1BM1ipGTDg6pkq01m
yTuEl9R8o7K6zZ9gr2iHfn9JxioZhis/UEWx6AKB3CK1H3kb6dTVgGgHrfp/swfN
3SQzSDtmJc4mZTDHMAFUq5KKV5JOaHgL/8hfXIWHj8fAGH3iO1HTxwV2se6WI6Di
1c1dtUBOMsGlmGLlLOMsniQwivCiKAYSj6/amm3pDZor0XY9YzqhrKzscAVohV7d
oLPHFfAlxL35aAcpSO57KiVq2L3uvCE05sHdhHvJaWzknhHhKTM9phNvXy/w9fVC
QVHVbPhUYK49YwdUY97BZIyF+JCBuC+L4tFB+XNh0wG6arUjbVOHfU4T1piBAyna
3OQOIQ2GNeN4lR9esYp4Y+FEwp5jcCvK7kpIJqJGNu0pygtQV+fA8Lj3GHRCAYik
LGp2vIf8ynG7Jn59bBl7wGvnV1lG1tJPiOvEoMZEC4jORGDwcHuxq8tazOyvCSD/
6givrnCKH6NFEETB7ScC7P41ZndbEjVuhTA0AvhbkBxnHGdtTwZPPw0qSuMwtP2G
zDBGz/eZf4C+x1x1oSyOmhaGFUyiZkYJAEsvl22VeeCRNgeXX2k6kVl1qoZT6p/P
QHqErZqbBvNCbzJc2naIig7+Scdbq9Zm7NKyKir4rD01LE8q2wrJlifxf1kAV+8t
sqm91fM0Id92n99IjVGZulLn2d7CR2558KS4abJExRt0j6/oYX8C3gxTBaWdZvB/
08Qj2XcvD1QFzTvKq3yH2RgFIcjcNWY+MV2VZg4FJc3/W2shXeyUCj/8M8GwCJRc
4mT04alI1qUqBS/aBcWxDXyo+az4BGEOIVjiBA9ZjSfGca/v0eor80xjbHBRVYL0
d341Nz+dRvbsvkrJ3zaVD0t/Oka8EJW6pVk9lawhA0PvfYbOkXN/hJwCXUdkZ9p+
Vg5wxuxGU5bH3cULy84oQvnhzI8HEGP6/f6F+DOhUX7PNmQBII3PqA+sEfW+buuR
qO3Jh+ztitl0emmAggFeERVZp3mXIEykyCH9j6o4br64g1B+BvPl2rPXMrHuncqc
Ea1wO1c3QxPsfk8bxp0yHoG68KPyawVahIyRWLRl93G6cJfRxh8Hd1U6DJWbN2Dl
QQy42Kge0UpKH63Shcy8UBMF+QyIEeeOqGdXvoancBq/VbYLGvq0pLjCRMxyQTBO
gg9u9nFkaPj9D6Cs72C3QejTpmcpJaUg+xS9Xy3jcTgHhjr31rm7+GcrjjT33F42
T/l0x/et76GBlfDfVCHhWijAR0Wt0GKOc/7a2+ixD6G9V5jiFEuJmckzvU88fHnT
zY0Wwq60H1UMqKz4gjiOMxYAaIhYECOUw9Gizt9CoqzQW0t15JLmp/g7imx2YrqI
5WL7mjGiiOM3vv5ECPme/BU96btzDLqS1D4DlMIvXv5oRf/rDQftSPhvcSreZabt
jfRTcZMkzYEBGn0H1lhQ2eqN/bQ2jGaI/NejWR7mfUEO/YB3hz1d4g1QjiYqq88g
HVaT7J3bUQB6mZBz45cLWoMdwP2yudm1zRX8wTtvr+eXr4fQTTpFgr4PZlRg2vIN
dT353FVBRsOl2ZUN+qtpPhDDx4+IQjH1xf3glA1WsbKdxxxeTDnsho7Ve0G9Edbx
2S8fnrhEKkqGJA1G/tbYMcxiIlwmyg1s9x7P5//VNvKuFX0dgBcFZ3htJuCrLkWF
D9V7z8CIiQ8SPWQ0RidAWfv2rnQERa1dPCA/0BtJwhnwbwqfAinSpAIFiwZguIMw
F3r7qzsaZoKsiKSbHk78Ww0ejRwZ9DnpI5jclBJnrkF7U3PEfmnMmbqqcznOdO9/
jIZD4Uj7bvRG5Ly+whbwNhgcS0sFRtIgNULadnS6Ld3qOp1Pf4dadGQxNdpy3Qvr
VWcPtjCE/6L1o01sFxDLocbulWJoFT2yCS1Bi0XErUGtCsmxaxq3XSkuMVzrGPrj
AuAw30zKc2FHrftCjUnqTKNUr4mPOBh5++xyV1Z8ax1txGrBz4x0bDKGTS6Jydwp
c4aG5kzcuVQtFs/TUl6MlTmSeyusuyQGUYc7nTI0vnzkkXBbSXYf/swiUArWg2so
dH4nxjSCtvcl1ZNkagYrCiYq3l1KR1GC6k+VvVozIMyNGcaw3qjs4w/F1u3zxjAv
QrYfodqMPLv3JPg24OFi06/Szs2QSjoa3UrtdP0Gwy3iWnhrMRkB6CkWvD/zgCpx
qOHBCBK0MKJXD5uBMUdN0R1FEgTjX6Z9FED0TGmtJwdXmmrReMd4X85cwhtJ9rHs
oRbgYf/QWncE6ndJYgVKhF9Tot9aJ29W6XNPflysmCBW4muVktH0uW9vRL1VvE/8
Z1BFXj2TcfyzBI84FqAPP/O7wxYFS8ta4Wy9Qb307MijTeDKWJB4HkQp4vuaz4p8
cGaA51dEGkECFb/7tE0DRj/2G6qcQZmxSwBYOvjsoSsyrbXJDxnAOkGrXUBdzh7g
n2mJuj1O3GAU+79T0NgTSuz2rnch57MO2KN4mhgkSSuQPhlHTs95o6kappW8X13Z
lQFLpJozYGzVyYiTeFuKuRB+jlYYdT+KLtFcJmseGgT8tFk2Uq0boURPAR4EFVyt
oP0In3RlG49G+CilSQik1+C624oSwnf6QM+SFQxqXKgpEXZ49ad4AJuiDeUHP4i/
RV9MDWa4fClXvBa86itAoXQntThbD3El9eHnR4026qivW7OV4E4WHVFLbPKlzoYj
7sKjHtxqyskREctkzDMQ9twcxI55ONcp+y+uCAcJFdeqlJsO+S1HhkoBMb5Cft+b
SGMlNhSwMgwQoTgerMzeiEkY9AORTigFYvHc27C4g56S24dc04GTLAnXi5RbOo/e
Na3jQ+2XLNRl1ih5OhnhRSQdvQRasCI9H1KsbzLiUBt2gsx8pzkz0PsPtfgxtr5U
5sN9WvciSUyoHlJ9wYAJPV6UuTK8g/74J1qiqSYGU9YPpmRIu2kisyimbLA9z+4Y
MYM7UhlqjBgsvB8NHON969pzMKa8sNhdstx40oOr9i6eYG6w6PCs3KPplGQYNoUN
TtvQs3ID0Xhj34rNN4SYGQh7ClHW9m8jqtMQ/ZW70AD7JcyU5vWLNWDmkCjemA1N
YT8inPDTr2dbeDhniiXlwMqh/Tgy4PJAWVWPpu55bZWErgyIDNJA2RPUGbpkz1DJ
W9A6SixjDiyGO/KdKTspiyTJNTarH3mv9VjNcn3e2gEZt4Gqu2/0mygteVuQ51kx
UR8Es/kGVy/zSyXgIUdg/KJIeYhgt9IoofCourven8KO0XCVfvNv7w89bAe+RYMB
HAHzJ3IMLa+wcvDH5BqNIyu+t2msiC0qWpvqaJpv1C07C4ViBubMkfg/HKF/X+m/
A4UNpD4yhVfIGTbPp/EpE6OSbxfFgDTBhqkcIykf0dup1p9cG9F5lR67xBy4qvHF
9wZVSmWV1+FV15B6VnzjI/B0ybHIDTDcwr0NyYkESzBYJ07DwjMKcQtIGCdgmpY1
dIZ6GNcY9JkcgnzwkcIjFIvr2DEvAFg/QkQB6YNUwq1fLzU2FrNLMP94POniXtOq
e7PgSCFhtkRmc3eV7rSyKwKcMHLZhRTGfedTATGQf4WLmjlsheO0J3b5rKR6mqTW
q4K8CgJi0ZxKuwbGD+SJMruTC9nQU/rvpBELnu9xGYljUSPN79HvsJh9w++BcxsU
Z8FUS1/4qYOmqC7BiHsEyhjItWduMaH9zoPKhctld1SIJGT17vYma1JK7TG48rAx
8GUtv5ptfSpPbDRUu6/eAIg6omB7zD4jLaNbZe+X72KIhpS5LBA/bPLf1U7anws2
FIvUWajSMjMcHrkQ9BmQwXkQkheqmhwi/7se1rQJsrTjs2TR6FRfYzd11eMCZIFG
IvtlkRY0A86jBT4QrYd1RnhtYs4CtPFDAHlHWROngU2mAffAG3nCvRhljGB/idnQ
O9uZORqQZzl7lhKV+Ph6wi6J3dzxvDk8zyQAtR8eEUtB0mKHmUJabZ4EMSXOsySZ
NjjXgcAOi5ITi45p5UQ6FH3S2r4SNT1ZVTCqMIrRvfX7jujoldM7hyiPdjRmoDm4
R78cbRGFzhNAJb2rgJl+KadrIYJiI5dzyseBdNMP4ZzmzFiHftp/xqvdoR9sqFl2
Lo1mTKBYY4tyGq2D6BlWonUxVunyPx/Mq/qZwSF3nN7a2yvTWBzmf5S/6fVhzjuA
JZgga0dr3DzWJGeUCPcQ+RqybNUQfHV2tx66ohuGmeDPTBnFRFJr7IcsW6fCY957
indPeboPD9+B6ciutE8GcqygSNCst9cpU96u3dpb84BzOtfkaMp5X2ZogbAP8S5Q
S6Mr7fIih027TdJnaihs0Trw1TSdnr3N2iyrKE7qR2GYi2vtQEt/aNwZjReYKvjN
fq5LLtSbsWFPbqXeQbjT7HPP81WsErR7OQXAMPFwG9kIfHB2ldIG8CmNQC1iFk4j
ik8CGfCrdj/1A2gEYAMBT69FcrbKnzBi5vGF6Ulxy66PzPSOgsuqysCK44+exM33
mgxWSa8AS361tAlu/GoYfbESEd+NxImDq0ItCFsgGSJrQtDD76F/znbCm/9HFGTR
GKLAkL1airM06wCEpN8HWyRPAKBVwz1mHg5GfFviv3eRoVhBgVVlJy9Zw7B0ws31
D/hhzY7XBcFOzUBWYukgoS0XXdAXbhjEuI0mRnUzRurlZqyuZC3KuNM6pegjjDfb
/Zm0W3KFi2W+Tez3El+TFIeG2peZ+TBblU2FZ5hm3cFLdc+Q0ti5o8UxmPkSK/re
NMFuKMWQXa4KKCxWAm9RzjuDJWdteNMNSeX8YhLcZA7t+j5rwOckBFPDbuE7xKj0
Tch7TerP9NztamAASaO/9uliW0SpJbuKN8myyBPaPyfNev8MknN7ACi8zkQNrJLN
hat2RgybVXBBgWZJzmLfGwuFe+Hg7Kwx808WlGd8bK8Qjthu/+tKXnpbwVLShTJe
6YctJ29upGunb4Mt1hssJ/ZTdY+G3IS6yZNE04knmKVLnTwd/DWwkANm9LlHkRrz
I83oK8rPY6sgEKpDzLg3HJvhqx/1JToayrrP4hsf2Dm8AInmLphnMHx4qYL2fg4a
F88GjF3knY+g1TEdBM3r9HZp0MXDUISDVH0YNu3QGzDTE8dVNzOOiVyIio7jB+2B
ps17NrUmjzuVbVSGeVCzdVkqmArGZanu7X4kFCquJWFINdq4lDUmYl8+mQ+z5aSJ
q9fqfvFaJXZxbSi9Xw13CqjzMN7FQodbG5xdnCgdQGtV/3RYvJMim2Lb9EllX+9c
+zy5czrbxUW8ScV8VtaNbBezve0qSFTJQdBz0bwqvj6lKY2O+GYSBOINI/9ReWjx
rdpA3N35jjBzbsUB3KVNZ1JKYJfDGUg8YBVsLdLf0EyiOz9OWSL5KPPLqpL4aKSb
sVGri+biCK48Ra2U15QK6HbkRySp8Ww/in729n9jI32MfwnmPBV+ZBfFLjo8QGq9
Sv0pYd4Rm/dR00kOWP/txt3UH9R5kldd5Rrc/q1aHtbofI4p526hHns2fUTPFhtv
7zxKhGMtcfPavg5A2kFVt+s0UkJsc5IV4HypDNG2BbWma47ygF02jxU2b4lomtEK
8DW1wzPzUvuV/3ZHysmwyhenVORvUhXDVJsYdYFd6ih/8+MdVkqQ6CVB1aAwBpFa
pJXRs/ETFCHI49h3FyxYFNz+gjvamKDBWNjHtUvyj5TKSgKXWmTvWHPGfoA2zBU5
7MwysL0AuDKFzbOQU14BFuj8uTfgRs9/Sy9qNEtg0BkxbAIQWx7jCvbY7PRaAu+n
Gd9+9rZBpxuf0J0mwMGPNsMJt346/41XS/zZlq5sfmaEfg8R4tbTyMT/1vIC4LuN
YgFo0YoiQQqmKoDwOwnymGLmo+LStKr8Ts2/YnxSFhgay1cXNsR4vH4cAZgXdB3l
PYs3iCqtHZbq0AQ644kNy/MW2dHTQ9cDs1VvzXDrwTGXBoBPiW50ThI5hcpYmssZ
tEt/+u4WUrz8Pcq1kTGUeLOjIKz3nC+8WLV10DHpDFizoeFt7MoDdPY3N3wEXqa3
inuBBOrMj5PIb4z8fR0VzR7T8J1rZk+AXRm4/1+21I0qHQVQP8OKOMDsnYkW8IH4
UpvXmijHYt6Uh4i3gDzCjkCl9BKok6D+WtvcPpyzfwSLWS+1emKLHe7N9vyWwnnZ
Bk6u5s42BJydYu/piwA+/KGajAQ7T44/d4gzgjGY58ik32/XTkU6nG8vUCPPCG/m
YPykurZUD0eUUILSUTrNlyYfHYZ0RW3hbgfb6r88nSNFH2ZRSJtU8xhvTwOk7q1B
uzWZsMrH9VuoDln5TprJwOGju4O46jJ1uzP425Xxa8ZVxte9/rFYApw2O/9IbqX4
SPCSSB/fow9R7e80mEZIHs20cVr/qv9HGdXM2uy1OXaLSu4zn61Y8FJjsjoQRnAi
/YRgy3NQEWcHiffdHiNFaOof4jeVYnTBhBlkK1caKrZgtW+NyYeGAltrevAkuAAG
0qRpAPM/ah86HuW1sY6yybntG54k/E1EhUPzPnu4OjO4vCZVtRHl9SwRGmQIrinE
k3YmOPSSCDHkWacw+swIEhVxMog3mcgSFFKqfmIb/C5KXrJ5MfGVlrkTTIZpYcWe
USFOlvIpncC4HXZpIuY/uN9ZuIc4D/WSGS6ZfOSqejZMvMKvP8aAYxj39qm4Zbqz
vvtY5i2yJU2nst5d8TYHu1OPVfmO//2ka6yqA41r7VbPgYU3GE7XYZSjS/Ht37mj
q3JMzd8e9DDFYoF08Ovh5riOHtJnZe80HNCnUfUCfzznrBmosB109E8XRVi+h/XN
bMXDHwQ9QhFISE64CiuShsKJI2THIp1ixCnZ1J6rFERwjcrWSGGdvYryzW4536Kr
k13eIcY18EOrVpCOOHRKFSkVYW3rqIDWEWAjfTF+nzrgDGSR0Nr04XJdoAbcNRtG
DOjoqv6BD+gxPvGYhpxQXGQeGyvE4G4Oijx447PLGd4d2a2sOLyPT5ksQ6IkYdWg
4p2COwwGP4UomVq3WHT3vFG/3i4f8343A/Lytrs9Hcu0SWLFZCc5X0hSRhfMevXp
jIzhq7dyS0sVNwLJ9OLc1KQNLKk+X4SgDfM2Aktwbb9CDxHCD1kVzH9AMrLCQDvZ
wvi6Ap9LQTX+2seHNGDvO3r0P0vFaZxO0Wjd189ntrqbPsWddKX18V64tgN9x0Iz
wb92o3IlVxRXtwNagSF2+9l45FXAYcvrZlcDStI0bkrhSohgO8yRWDMn7O+SZrzv
uHp9DnNO0sjprk5f6uly9frxnCEEX+VmVGtjN7nKoz8WfApnbXFW+7rjO5QoNv1M
hTp3ohj+ibkZ4xe7uKns1opFdZLQotCyMexn1LAai1J9eZJQxlYdbBqBjhDSceXU
xg52JVEoSpp2LbBJC2WlRPkzTp/jFHV6BuRYR1hHv0Oh5qfwykUnAJeyCxtCXtmn
0k8ktf5g1yFHhL7nHbY+LO0hqR4Dbs7q96w6bNRySX//WSiuMNgji31X3l89Cr9E
1x2P/F8yXDrhi3jVJNNtlnX0qoZIokUePgPNcLNsw+GUFq+NBny7TKJphvjfMjYF
++3pzW3bgYYpZZW1jSyG+2qncb1rCZ03akLTrhUgh/wXx0XQRDurSNm/DMvFMPy5
oaC1hVa7tXT2lJOwaqWHLM8+SCXwfPhWVkdH2qcTI1pO6Reu3+kRV7rSFBSGUGsa
XFyKvJQY35uWQhOGKP0BzCMk5Zby3G9wL8vWMSh80hITOYtusB7n8X9tz8cCihiy
6zy+GjPkoX5jIfAYkNGeBGjIddCPvjF1CkIU4pkZjOXL5iy8kDof8uaqAygu7pN8
oOI0TpRER2vuRMdW+IkdSf9ZO+SEqWqDE8oGPBRlRRIv8FWbQdBUY/JlFCoUFQEH
R+rdxfbaodM+xCEk2aOqnmLygONLvPx4bcUnqvM2a8cO7bfLNUER89irhwoWJh6G
8gBfQc5HXidRMn8EifR+SC3w0w5k5fPAIjC0rWDdLuTA8OMva1adwCcAUEZUnslh
cnRsEZ60gwpQAsGZwItotX9FHqNT524wcBlOXMOkneWl3zWFD5Iz4ELCBhnTSVdD
FsiQEah9wxpYAYbLGnufRKsxWML96Oo94FCk36I1F3wOhAUpsfJBqaVwOLMvFb0I
t/TDWow8F4LMpNQsHwVUZxonece/FcwCMmdsxsFLHJNN8Infvdze104Noo15zKi1
5WF4PbKVrwB6ras9zCBeQv2MQz1FzWWVeGms/EFJWU5r7CA5ZEIgeQ24NaB2zF2a
1S7+XGaB7BQ8CntiNzNnOeVvRs0fP1n/95WtzNqh12xZUFwdhbtXfMIBInVOz9k0
JxOuP6gwuiahFcgxosr7dF8u6oSh2aXivZJYrMDHEOXBVoAain6FUixevDqelnXD
Ak7CqOlrM1o6OS+BwJy4Ghwghi6wRIbyilEQeUZMNNp+U8DkATEVNLAO3ZEi43gx
CvbkVzs5+a4k67tVflnkCwvs61NdRCMqICVzG0H2NEFlEg9JL9/SdZ0qXeallAw+
rtrILjLTEWq5eKeLxOg8WKsL3jxCcZn0uLaoIbjT6agPzKWYv1W10J8wrzw3Ynvl
6iLHNmkN9xN37hjdtY80fR19EGzyZ/aLl7QGW3s42cTn37Tg9WsMFw8tZ/utOeno
EeOU6fpwDkEe3sn4633mO9dGLZmUBt+Y5yG3HQ1jsGOVKv9dO5JWbgy6wL+XSqbb
+7SOfaOIsGUvpZdXJTinp9/HJ9sPi928mEz2scKGEm+nlsqqxOgehslsxWK2d+79
0Q8YgXvmVmoZdnNt/yMr5QS9kmzPhb0isU7oJGYezmK9toXz0Up7t+jHbuHoDXS8
PP1in+JDZS32EEH/Cu2t5SqzIJjoiR1tYv7/JsgX4zSEtLZUilApOmFyp0SjZ38n
Cy2rNWl1dfdqsPIrELtW21H7L6VhU8nZbZJZ0TFy3J7T2O65rlO9wHmioMhATfJ+
puVDqth7I/GN/QrG8fie1UXTWN52hAtYUNbBsCQ8DWjLPZyHK7CtEWyZKknNJmdS
kCHZNGCV96Nz6gSXI5tEBB3qd1bXq4UJa/IfXpnWUg9thJcDEt6u7aC5XD0VPbzR
tDbRtAXjPI3ucsup0bbPBQGDYSM+SabnJcxZppNzv2XPERs1g53Ia6exXTSi3dbA
YqjwX8X4xO3qI3vYyT1XL72esckvDHWmuBJPY3R0JBikSM6ZveH8/v2oEnNP54R6
D6lTKZJJ24Yr+Bi8l+IGIC+aybxjWb0wUUX8MZAgcKY3h6BxDF/uN+CtzGmMDP7y
zSspoudMZCtZCYzC4AcQP5/ateww1JFn35NHzwGG0z2dwYVymAb+XO1ZShjGgsoq
442UCjLuYVLal6JcerspwSsVCdBNEynzzoyXl1ByBmy460/qUOLfWThjjf8kwN7Y
cUCbGnNzTS0uORS9lJENX1An7s+j0Jm5Odp9yaPzSQmaUcAXnS7LWJQKU3IG9sZ1
xYa2Z540eDIUpWsc8TPMUQFBDykbfwK9h0W+7SxPnnOg/uUbw/Q7bb8xAQN8a2/A
1RQmQ0kY/I2kBNmsOmudMYfeLPJ7QxoBsBZVltVBU9btPvYo4trx9FFyTxmQumAb
c86zWMefoY2yAoo3JADG+r/tmdicunvy0lrYZgk/isNFKI9pEUAoAYjl+oP7lxz9
kNi4+k6dZHlc876xZN773KPbmNeogD620EyWtMtZkWjTqmY3PP2Ryp2r0hXnkFkx
BQamjxhX6a6awCw6Y2TinNyMxHazJIvaBMIsh4VdDWTV3Z8uJhxDKrTgWiQE6+wT
VI09f4lgz4/DTb5QzCnkMjvZOeC5H49+6H9pM1wXfJTVWO5eNlF4lVcZ0MLvb2Fu
oc/aDnrR8aFw5M0HScL76JW5/DJlaeaAWQBytD1C44zpo3Ez9au2e/zz0N7T0L47
OpfwOJlz7hvEL4ml3vcA2P377b7nb6B+IYiaTlcZGA+VT8nlVxmGpSu8B9NIfjrT
oOcT3Y9fZVMvR0KtKcKIAxRD1KyF+CVeA1if1v9q5YC2yZ+trnEV4T1gmOYQmRiV
SbRSnacrMrh5b3SuAYIPMyeEgCHNvKorE+GGGo6GaH+VPYjdZNFpx8eBe2rssEl8
CdBoBLU1ACyIuKTFGFVWiqoTsyyI91us1OcTG06fBgYSeBg3FHM0ZB8ay3AKzrlh
9Ft6K56nvmy1lTeThkez4oMhiI6YN7/K15yOO4Seh/tpEOPYoROcd/muHL3X3d1i
EWNkO1EUyqqffn2ynPg9m9+sJW6tIcDR1lZ78l21Uve+VhrssdWxjpg6BVBsDh1+
+gP2E4dDfuRJwIJjuh1pCo1yX70XTk6HNTlQdo9yG0xtZ7DgtCYGch2rnzmpCMW/
fhV4a+mV2GVaIwHik1dy7fIoDngtBEAbON6ft8iF1GmFf6Mg1vU11VyfF0Q5cnY6
890i0BE2aIr9YUI1xT1YesaE/I17LexwEbGLBy1cjSeGKWeMq+G/QgY/S8352YEk
YfHhwEcSFyyP/kzWO0jjTgvo0Jpxio9Xn4aoip7qLOMAkhDKlrHU//3eSj+qzlko
9S9ADvMGtJH5tRHjf+fI5ovb5uEABAsFimK+y5j04r4t5zuDO8RMK7QYnFF7UyLi
/+DeWd8TvIx8A2EL/Y3jjYtc1wCgVk71MlON/JYbZ7+4Wrr9ZRA5MAKUAVza/yHu
4LxRCjJCfSsQr7IMyR4WZ8gQGt9dv1NOk7ktmxzbI7ys55XsJ4MwbWbI66W46ZAg
YWSvUM2vtCXQsblYlvUHwkbWVvsbLLtRaE2a6fDbOuP+NB1MxIA7zF1OpJkIGuDV
FbwZpqOLyV604JVM6l5HxYNsYtqWl+3NbVU+llrxAYFjZOsf2LfOmZuzXDWWSxby
AYjrxBjUSXGt9evYjLr0YpkyqO/XXiPn27/4i1DWvK+j8/W+6zx9cBGqyoPupIuG
AifpJUg+CbupbQbAcHpGZUc1EgBwqqIxGDR9wvxJOqvqDoyrBW9Z3gZ1qDC9umWt
q3PjN6rYrVT/NjTPBurh7SGRb0/ObfmMArXtPXj8cB6T8mh5C66mt7sxVsFz2atW
gTC0bF6lcfnTIzSA0B8AOLZ9XU1eb/ZD6hgAMM8DIkt2wctOIdEmOv/314ewCaSR
cM7HQXpKL8nVHoTKJBzrpVzxfksnsTfA+BtDsnIZeXyHDFohvle6zA1geRg9ew+i
VMS2NHmq0B5ZpIACxBdOUrmg9BQjJEZNGTw1PGe26F349pVXCt/RZkASnoHjstqg
rSk+yBZf+wpqn49HvDe/SLk06gs3aGUhB91WbVM+6J2iXehNm+KYqwLHxuBtXeia
Lx9mrYviALt9V4FUC5H1ymHLgUQX1kWPhAi3l4ioXvtJd8Api5J6eMkfhcSbeU8l
xOFq0Zel8bd832c94r6JmP8PzJCWDJ48ROsQO7Lo+9Gt9lqQPRJfJf55ZIZh4mYY
t1jyFUMNQfYHj3CBASRpb8ZRnGMAtGJL/lCLAoU5JULHCkCnjYn5kenuzSJhCJlL
sFCbv8eM2ksTw0/1ewLDxa3yMUT3LkWYXoWEnLnqqZIAoIxe3pUbKbxIDjMYb3Ut
f4ucGNpFXI3pSigSmxpV8kQXp6SM2jTq+8ETySMd2GKSXIhwRjLzN+wQfFBfaqbe
/yf9ogYnvgarvLREGh1CGy3ZJPIn9gkzkJOvlLffNexyXjD7/FwpTWhxTpYJ0oja
9Az57Cw9L+YCazdWrsuvSuEH0jD/lRTgn+JdwPq2A1Rur6Al+p47GFtAM4eXmsQz
mDp7gktxHijFo5IjQRgeysyDIdqNX+HmstcqrRZ7MBb+zXnCg3DfuaTZXjHhBwFL
QnKaumIqBHHMIO9gLhLMYQsOpkc7u5hV9ykEEA6t59VtatPX0AM0+Ey8fzmEcT9u
wR8R/hQRvgM5b3+m07kTULkcSG+6Vi2su/lyTijNIhiaXXLGo0rLDqIToJ5tMsmI
HnjYmiGobtef5gFkubv7Er1NiV3qnnmC6xYvniAWoD4zWMmksojgybhP/n0dbNgY
K6w14yUrylsykKWpYe5XNbzszAYBANaf63xHAnY3dRk5FkavWOksd2VZiuH1J3QT
a1Mf8S8i4dSQ6bU3o8BxjOI6ILdOIGIkkdClyvT72PDkR5FRWhX6J9sxuX6J8/Re
rnlBIj6krC0Kh2J1cSYjghBNO/VJqwidUWcsw1laetubK1t8lOdXMs4m5nm0Ln8p
2UH6XkrviNZzdfwbOPfeSlyCbw5+OdZoh5U/tQmHg8w1RVu0ornyYcwNVwgJSuKJ
EIrZ/hGV0243swpNuSHlsZol8gDC4UPenu4l81z4mqfZ9mQNoAf3GxGr3qE0z9an
j0AHH5yXKuq7qZkEjFSgT8L71IcIhfSKWfyevGBzGrKz5qZOnzymztPU2gtrIo7z
xBaS2EbkhM8tWdCJD76JqQeAmptsmj31jCKUVXliBUEDXFDaNPrTj/hZvJOqoHr4
7MJimEkl1d4HdnOOSvVeVp9Xq7cOZdZ2lvkjTxPd7K55wa3A1+DpneO11VKqHsB7
k1QcqRb5HN1OlBNMGTfB+pG8ekD0EXEzukDlb6w69t38K+x2wlE8imiE5dT5CJ+K
LkMwlVoRz7WcAWvScjR1M+SwqJCyvUfTxX8ah5dzqvxYL3fJY+4jTqA9jxFA2GfE
11sYmfJdWRvL5YpDi+KS9Ga1t0IrRAyTal2Dke8leQ3gQfZaMXCOZBqzW4qsEMdh
ILRIG+EyLCCnO5iYAfv6BRqEA3lmm5YxpwlkLMpr9OlITqAar0EWDZf72BdnmxfJ
sMEWJYISIa1Tcg7b/NyQ0hSrWuNo2GFnScl8VT++zg8lO0TcL4tkfLO0THqWfFx3
UwbNQD6DIdpoUDlslyVxij6KA4thoxTIziLOjl8ppepVOBgz/GmdqY8lRhG/O76D
F/WaO9BmiMHTZYz27Qyi5Ccv6DOAuCYqTj4UZ2XBVXIp0ZymM3m93jpQ7xznjwFs
c00oNqGJoe1ehf5zyJM4wJTFPbWLF+MFBNDwhb2ZLBxSKKwi0lRZwrEoXpEJ6vXB
YSFe+OH1SUoIH1rF6WwltXKb1pyA32oK0633l8+ucr65TqVrSMf5CIxEVslOx6B7
M4406nniXFEJ0xNJq0JTqo8wZrlb/YIGsncGDEOwuqFJjFX2nMgdTUhSS2326ILJ
/GAh2KV4uYK1agEVqlgfhIIrPQvCukXy2Yx2MJ4PAk/ara0O0mcg2D92GPLnnX5M
zeSNGCdpem9pn1qQvMadpcO3VeQPh91htPQ0W0mmRvfErhobbzWr7fSFDKOUu4gN
H7IYPH7iJneADyM/amw1tGvTots4DfXlxHNZgwL19A39+XM8p5t/5Xvkcp8rGH0w
QHKUivg4hO4UGbBy57TlH5QJCGgbcuHmlDTkH2D8F6vuU74T17gkoIzo16Vxlu2C
mwhn3usNCcl0x6RAyvUfqXrPzp0GLZ2tgqWqbtSTtze+MAhFTklYpPhJum1qp56o
zKMwYVoL6rygNyVFmwP74w8Nkg49+VCVfaX1UJdMEKe61DmH/BjLexQoPU08GoBf
EYl7Abql/vh/X8cL/zYRBod+36EGlZRNint8qvClOdXOL76ngqzcHmmtgTxCn4of
qz3TklB8gq/5u83DSJP8GAm2GD7SrvQQ/j6o7zcN3XutSzHxatEELofs4w8/wktu
W6eVwadEeCT+luYfF3bGLX5wkCycj2+p0DW6K+8mwZSDdnZaSUUER19VTs0dUYhv
veFGv9XwFQ9T+MHxeV6df3a9B3YacPEVuqJMZtJXqK26OQNIZFhw6amOjHNj6glE
VroMDIsopi7xlik80vNrHhElxjfz6+O+aQcMUv6xjO4OfByWzjKSZ6+gWunHLXSK
M8Ce+z7hzuUaitjujCJV6MYhymzwG98JMTFY1X82Wr3kb2p5k1+VDjfKnSEdBlIj
EVS60AxGaH8f8ZR6sovElDZZri3CkmoL2yaCXCI8F194sltjkUclG6F7BBSwcw9I
aNKKgaEHxS0JCfRQIbUjVBBHPn5FOf619+bAwwW2MkgTVQMmTf6Xk0IKHPnOEwwd
YcrATkQX9w6KER8dQdNCpoft39BChcB+3LU7nvf+V43KJ0748REfQR9hebt7ve3/
2V3dGf34hVWSchtKkW/ckd0OeXWJxRxkVurUD6f/Bs7shlG9ttkkw2Mww+TsIcaA
WW0JYUG51v4SsqZXvBABQxfp9+/RZUXaI4+7+2L+/6JaUi5eCCOoryaG8nhug7St
J6o2N9RRLlCwBHN3u3Ab9R89s0ReW9Dwt7YyxYonjnA0pm40IH2EU+ndv6IIiock
qJPs98p+nSF0RIOr94IRBYJCXuqGPuQEt0D+pP/Vx4wiwq+vCKbM4dsF0Si4phPR
cQ6IyPi24se38ir4gWzWXFDvERaEMy8yUvwMH38fi/PAppVvDxYw9wLBc1G56qfA
wmjXK5yxGKOubitXEOuxPFAEpDQcwMdV6rYMVBT/+uSHkjPpHvOkrFk/S+7RfF99
mYA0nyw/p5eXrdhJ6p+QmduMxc5l/bR2fu+f6VkEMfIknWP2kzYHvS0KFBj0cRdY
y9uwaj4D2Xa/1IX8OjPmPN8qPbdR+Zd7hrncSJ8TsNMd/jSsA4wpHi02G+Ckn6pQ
rdx9vRt3VMPa/68wKemrnitENHeyADJeiRjj0OGY+pYTvFMqtyz2Dhfuh6oKeSaO
a2HHi+Qc/3CU9KGwHbQLlnG2Eim5aHs8V+zQWg76+juo+kOxERzNPZUTVZ39V3Nu
vkwkP2QjR48IUU9yQf3EJrlGEkSWIZzcDNss7+tjjnym/Ar3sxNO++QGSMSiS37A
LszzVw3c39a++nwIkCtd3JN+vn7tY0ORZgOVBz89XRJA1UUZJA+9uUtFMW5Btgle
0+mMN2jYPt/HOAb2+JX3dj0wb44/Xutu8Fe6zMzIFHApnIAk+PD3WBBYZe02BgSz
JF1yuTwpQyTUJJuQFEmo0im2uVNbilyaUwYDslJC3m1HuusVgJMeEbYSqhLf++xh
UnaozC3kWUgQmga+9fw4uiKfJJvVC5ZvPgy4leOaxJ4Yo2OPTnhz95c1ueIpwzls
SEGHTpAeJtpndojRf7WasOqDVSoWtryqhWHXlK/I/zR9uF9V8AGIhwRm6JXJQXsC
wuRLv7QJfNnSHmHDj3kd1uZsX+jB3CwzqqqOgAPkG5JJcL15fR1iRyGx+wWueb7x
lGDPE3rqK/KsWHuLBk0fzeWh8kh4sECruUknnNXs+OfChhPZc0z1//JuDPQ2FNZ1
r6jFUpDbWqxr7Fyi9NqVQ6z+e6wMWAWARJS9aN1NqOB0ktUKe5H/v707jpqAItTw
4lKq8SPic6oKCyOM3mUjhyaMvtJggs6J+P323HSigU9++pqXPgkUpxtacutfZe/J
zPaBhp4wZwYEa3C9ja/ckkjeEVGIOMZCQ0BK8bVhNPMrwNvJQMslLVAcSVNJOs0S
+yiHIxjPZCM660SSGEku7cv69+LonLUtJKfdhk6nGJAGTrU+WO+nENdK4VMimySu
ofmgpTyFTnYbeY7jTj8iIp87eVg/H7d/u+wptaY0i/ZB6h2RWKxJBeVG8dQ8DyVy
pvj9aOCAiRaa9l96noD5bHo0SWJlE35PlwNAqynR5s6FQvpfQwv3xwA+2jBAaC43
pg2XwySLuLdtsD1JragX3HTFjDwTK0/7c4taEo9aPlxwf5L3IWW4nHdJZjgUPubG
D8KM3qvGW+o5DeXmiuchGozKlgmLP/sUAbFVnciZavhm2evGEDuREQyo5sVRGTYo
cv9w5EJdI0t9pm658GU/OxAHOwayepzqNBKgdLvmFb0eP5hKNR7v76y3fkLpZDsF
nppc/RU4d1+TMeVb3/+E7P+ouRbdeekSEzCVazdFdhuQ2VLrsgoXkq776UyB8uiF
ayROgCZ0j5JoWqnI8WpJueMTyhXpFYC57HrJKUQLChCa5z2Ofm1SjnT5gk8nAP2S
a4ZuVPqkAeLZKiBe3bqYwvGIwhgjL+kfzR5PlBTnSDuw2zCcBwexo/9EmG+3Z6I0
ISxHlNshEAcukdB1silbn+8D7k4mN6Cj74Nh+8LUXWnN07HCU2KDarBE3YkY1gNp
AWU6zQW7vJrT6S5G8apTzNwyfNQrDVqc3FFaqTXjxpbTPafZdw5OF+lFUaxSQynh
GKsOXwJqpiJitIglLUk4rX+4W+1jq6ATI1EdDGpOi4zjZGsaPZA/D1azk5g6koRf
9mt1QP3Xwb81Ph+ynT0enOgT6il+OaXDrKx9CXpWzogFTI7zY+wW9WS+JzjLsHIM
X2YgKWKtGjITGcDAufu78sw28X3Be0ploJrFB61H2KO+VwP4XPIvctPCzI+dhbKM
/eZffCNh/oHRSGKLqxAnh41tboBilyvMovglCzP3WlHETvFlutIOZUiO4KFOIMtL
CAnYJfD4CXFhaHQ7eIpRmlTJO0rcvCCNP+9H0kYK00p+1Nq5cAfXaR51kS2GCGri
pwAOb/EXHweGm7DSLTKYspZo1SdMXX4mljo7QrxDih3Df3OCn+zYGnT9K1/gqHEF
dSkoW/FM82epYRuqCXtAOiEeywXbv11bAHzLRqUPIQEGEDtizsaqaLqe6QwIfEe1
g3yPw6vyeypg3vN+NS3mHqUlw0uqn8j/r/jti2m4Vqtp8n4HF2O4hAnvJrKZ5qwc
g5pEaILBQBkrrT3tKYHWmtWxxwE5LMw5aXRDNqF1ZUcHa61Ba86pnSRoQ+puM/PY
/9PCwcRr/4EsLYpDj3yohZYLn2skWoX4PzsZEZuvS6OZU0Z0d56WF/tH6yHOkLDj
pabpRIkNqHwtxzemIgeU7XVrrW4KxcDgyhfGSQtvqE+fU6D26iVLqU/UCRZ87GW+
ayVZOHaJiRd5ZKfVOBEAoyzjZaiBhF6fODff2sJUSvERfTFF9b71mf4t3avC7+pV
ouZF3DjI6gu/Xypcn9KvZMSeMl61xBXIE/XqMKKLkpiKC24k0aeX7DyDt/UMKHVh
pLw/VZ4EY8F4tnTB0JftXQkvJjsOoFn/0lNOGvbaUORlzhWADr1C2dKqygVVq2lV
cDiYjid7s4XL0sA7KoKeNY/XFgG2p2GtTbv014SSab5XzGQBLf8JJStuhJoRArZs
zmnPLi2ukFGzdfaa0YhE0cfxR68GE3XFjqZTeaVP85KOiATbh5jmSOZ3XXwTduYR
vfwT9HdpaleGqJ1OKmiuJPrwJO43Ey5n7NZ2iY9CK/OZkPsHs7Yji7F0V7xdKCjj
o/wqeDTrBq9lGEivaVOwLlX1QLEQ3RsK5AYr4BDbPjFwgUU7uI7ynwuT7IjbY/pZ
lklhodVZB7OiwbQ0ChMbHGmG/y1IN0Q994erbftlx331cg5u2jZnOsZQNmv+e/5f
xEQ5+bM7qk5y9KERTBaih/jH3VDRolkbQvS/zSUtSS2SeAPtbHsz7i2m2YB4lQKr
CUploKSazqh1R5iNm2gzdNqkfT3SollGx1HEVz9MBujEE6FTMG754IElPqE0QPj+
8qI9MHiNmHuZqd6nnlhKtTXTwvaJd4MSM7LH353kSEFDnAp8yPLIEWytrMSBZqxL
w/zxx3Zmek3NrdUsmFoNwKz7pJr9MXp5lx612p/zLxkKh8eZeLqrt0PUijLuAd4+
BrpjxjYZZsUhLpSVniHZA+NGmlKIYwGHKhToOTxOaFSf6xIrVcNzkxXSLfJiPI6d
i65Fg02C3eO5vNWKx60bkqqJzt3LxA8O/FQcG/E5LgaDyx6QsWT+CHZP1jNawozr
ZOYBirsJbsdDw+MZAkkcYkgQErIL1lIv+D/REkVAHpGpdMjCuKoCaMUVht+vWIjB
Y8CUajmwaVbhtDRnQ6sBy6GW55O3MSduxR0JOC4copYtERqPxIOJLLV3Oqo6jPBt
ZcwBisIW0gwJ4eAvmOCofAlhWYuhlehGfJf4cghTL90EK+s7nqZejjkyj23IY8qF
OfIOWkAtDtGKGDyNxCZIogFbXZUyxXJ0Spr734M3b1PEgGjbvcmjVCfdC1awisIj
GJyXrqUC3O3hng7kj3e6BDXvFk72TIGYFCODcG59x0nBQNzjwR2nR2ffHB7h1qm7
3ZDQL+8jK0/VYXJ9EIL2SDMPi5rv8Yvr/B/TOaA+3WaJ4yEbwBNg8cfmqsdJmScd
2tOgg6JzJ9jP+C5/l1baEC3H+GSGzgStzM+UxnpxbLND3eaQllupSRxG2m+oCLv7
wPf/rOiwZlJ7jpUvLGQsJh+nmLw/0bvk8XohaoX2DqcpZ1PbY0Vr4M/gJM7wneM2
HT1WRdkjVPTz0pnEjSaryrDp6vLyLQR6pqjdMUEnI1N/mzJdzOVs4KL8TGIPHpim
J46/MFk3FbNymZ0bwbhJqjDj79gS0XPAFJrbUSnWoBBeTYDj0Sgc06kWMKWyVu0E
o1N27Yw0MUBKCTtISej3Xl4iNVr2EvQsW0diLPBQdlc+BbklufoLirm2VppOaJEV
AopXC37dX0AYlmzRAPlqtjdt0tZwIK81AqkhLAyr1LDJJASCRLkzKHeUuw1MT9A4
MQDEcos5kEsOUYDZrtMD2WWYumEjUTU9NNRa8ndrQAdWDIXURxHk+0ASfzK9xA0N
hEorLH49ghfaR2U9lawS8Ur4PBONRXLRvCLUPnqci5S9akDXOAERqf9GQ9mF9sFS
dCBiPfeVj3PQIiksr85hxAD4WQYGoLtxNFSUwFlkALgkYxqQjzFrN02xd8qkfg5X
YU2ejO+TxWEGFOwajuJtNBPUpnrBilqxnhLNsA6aorxas9D+9h9rHXJSMVt7hkPC
8nema3ZF25mLM3vuGx6pcWbJZg6caDV4KPt6zWElFEIX5Gsx+2VhpwZEpKkC4oEK
6MxWAyvRoNlCPlmdxGwblLJ9ARi2RdJ6yctmCkCrcej5pIJq0psmzd64s6SNsFKU
UJyyhNRnXVEKDIDQaMQTYVjkR00o7dLBTS94UPDiJg9Epsc+n147Xf0Oe/0NwKbP
bLVJXHZmAGGgqnHE8Gedx0B4FDPUKpcV6ZxpUFr2lU0Z2TG+//AZ0z28h+HnCv+1
zwsXNyE4jZ+pZlLymvhbDavD1w/1a1MoPPob6pxkNLqju6mhL0MnXqwlNOL444w/
jpCiytEsV0ObJ1S8LhIncHVO+gxU49BW5AuXLLTGaz0moxPfmVv4U7vTSLlT6P8S
4J0mZ+91q6vXgI54S2rvNBHknXEkKur8VY4ObewypTwiVL8YZ7eehSm3/WnnSM/C
HvAGISrpBnL+ffi8Wov9o6ItJcL34Pv26GEOsLXdvjRZ+kAiSqkcQD+aHC5UUeQf
IzmdiCIo9pzpmxDdkLK+iFrWIgbBdlp4h2h87HyevB1FBcpM2B9l3MaWBJnvZaDu
yldK0+erpjo5v5652+iHhcodjKGzRNoSrckKjOWikvH5bzld4FWFWNR0Hlqhs51T
w7FHAqaQ22ZppwSWTSLz6amagthpfTJA14xSxQiP2ASeLJ4ISI9r3auRqtiXDIit
NTBBnjUMMVlJjoRHs1XcU1Sz3hXAALhX1OmNZq2o63YXMlUeY306nVw7pWxxxPmu
vqm5/rAMwltKTm3ETfYkn2fcuNshjTrSMDg7Q4RF4iCGy+1XnFGkAL/09rKkzvXm
SlSVrVyFqeAuE9g0vhcTfWMKz6hF3i3ZcU5i+PUV1jbCW901WdwlX/ppioaRfNwo
wWe52t8oCPZP9q6DFXBASGnYFmUCVAHrZTZHLEm1v+Ape1n5KDtNqFzB+ctxy+jU
xqZrq6ZBOw4qS2XNm1x0dlqeKKJEYN2jcRmbpLWBeHSPpiWtOVKeeyyBycBhs3Z7
KTh+gcp6EWhiE3NoZChQUEA0H0ftGCmpxLC7RIeXD5MJ6zAJRvtPxrjvrT7psId9
kDzFhGHVprG9ivj+LrVE8mlB1tMjgx5fwXiPCkj4NwLNpK8ad0c+rqdPYPIqMIhY
dd3hk6zKoLiXZ6CbV4jlek2/JcKFEQToQQN3McMgT1AccICqJu3sPdliN7G3pBt3
zYRuXkkPkrKoxN/wzLGMzhPGVAWDFlghXGUh66auWrGXR1hpjm9EjNNM22oFGPlB
Is4CCZI6ty8eeGoCie2rF6wxZ21eudDssWs3yLrM9hTHPtncdD6hmEFV8LEPpw1E
gTZ7G7BABwDb0KJscycN7d+di4eOURHMtHM4H7bSnRdiasCdEFSTgxylP+KUGvsg
FBd6Uj9ICLNozHmxfhdXbFSYCZbrg3PpXoPAxeO0sH9iTQMAh0eY8La/jo43lXo1
T/mljOU/DBpXXGjs0e+FXHlZB0RjETVcn/fhqPiQH6Q9X8nGlJltwPbN7hZvWcTx
9GASOUGCJXKjJfYCWZBj+FM3sGjNZPG4wbQsZMu/XetBvwolNwrnb0LSb3sZ5dO0
5E0jhhdAzTbPQtHRxLEIa/ORuTin4IZl4iClYKtTg/cimZGVuQMeWuy0QANCimmt
dh68csDt7mgJ6hjAnmQlL//PnxL0X65tndUoXVuEZsYtNqNgT7Eew4xiJNxJJFV9
Ju/fumaSFqGXfW9YypaJrhftAUuFc+jrmpIhMdZQx5y5n5ENmiKw8su0p4xcwsvr
vBxFicpgIEMXTVTYg1RdPZ9kVXNjObUqMrhJB4cmVqhZPnOD9KTlr/csbGDemVQK
dFQFo+FoeL3vj6mxWolND0HQaynx28F/4M4SxkXlIxkLrFmZBFZzRL19YSxXMTR+
gjE9HGLAOFjYHDK3M0ibtaESAi6SMW8pNVK9BRgd16neYpFu0uoFBhCd6r77pZ1I
y6C8QZaT3T+itdLLzB/gxGvKm4uHH+zQ7hT74+hqY8jHqDSzTjNOh8MmGa/KrTfD
rMFRtZJYG0FL7u/YKIbzVreVEUGvpLHh8TQ20MnHNzuGn2MO99WKBHHiJ90dEHM9
06SI5cHpVJVIPmN2aZRzRwDQekoHcz4pBuUEJYb22Os6Os02EK/hOGLJRPBUP+Gr
LhbvjoF2vP/6Atrpf0PB7wlYvVDJn6ElDQL6RZHUatXLATQ50WNHDn/NaGJR3dc3
QP4CsqId6Ls3zsjfWOCVrTc9mU24j1fa1yQDHecoqJam3lCpk1T6mCJwvI3atPq3
D6u7OChODk9LnN6dVyFEwtPSjc8MbQzTWqUqRGJ7nZGpXAkMzkkg6t/7PICnX7XW
4mMMlYL1og/cve8xjqkYMavkQhN6kPzxq+MzrGJJCysJirKUJaXxwLB0ZHGqsmSO
qcY6HFWENF+s4esvOWrtQ3g2jacjxbPlg7w7hNZXEeeXWUbtFdTm9AgdRfyL+2fs
1/8lXJk26U10ZX1JyF4wTCbPyF+U4xRNGFIRnW8DN3A90b8vMRq63DlWmBqvyYh0
JBgKJcJyqPi4g1ha9ur3aICccWPDZwoQcxAkVHB6TP/l6ytRwOw8LkBCl5DyXl3+
M6gVIqUGlleV6Xwv8tpWJdL/uJoePr/W7boBU1EYJnlwFuDaz7Jvo6IOcYFI7YCF
+MU7Ua0QUaxYquTXGpU1HItR4du8bjQqUgzrgusOvyJ7YG5pOCxkpaFNeY4+aF3W
NiUD2C+kHISBHUHM3YxDLOflm3mRqFEQJ375nH4y4tfjNWjL/xG5fTEOzmGBnU67
xDva+L1wVeeJjJT0+/I506auLNpNabxpn2Lc94n7049k/u22cWa7+hNGz9dfCVt5
0MiiTKX9KA1Q0DyH48a32R4I7vC2CVrBoVnKXLJYEKnkdKtSnR/iM/kAEsseng5R
McfqKRr34M+oXx7A635aeVVdC6e589QgifXQDZ7eOfUSFW7pLdhq3RZ2kOHO0djh
Ehw7wq5fQMPWQQ0DusatpQ3UFGJt3ArCbVm7GbIFLFcmMNwQlHbySWqa8ptJKsmG
LgsWdjB7bwPnX/Bf+Y9RJd+kGVbUGhvwC6SIKZkhRUnG5MwjiKd90w/1RqipVFwL
cby79wEHawTPNS8RcehbCHe+6fEertF/0qA/iZelMe9l367F4tlTsYgivEOG3uYc
Nt1VAgYpfaPo81cNuDqYtA7mO7QBBlD/X/JTk5imqlK8VaUbCh/UyIAjzJe2tnT2
QyzOMckVNCWjUTjPgZXvEv5YXkUr8jm4lBCkrzH7gUFKDKWPeOj2H9R0CSPT/hz5
lGGY1v/PL4g3QXINzyJ36Cl/SI5zm9sK6ytGbvIREO3V/VMRFBz0EUHyBh994RCn
2qC0Bnd6OaiHTdGhHyygqu8T0yPHYmwwJRTjOo5fxJ8ObYH9MiyLgsuSdJjna9ZJ
2SwqhxNL78HMDcW9e7yTaOhLPJSLQvIsLof16C9rLbNXdn5U8BlOx52FPcgggRVp
zxFN2HZOUzq4xd//zjjdCe7tWIlsH+/x6+avRBlOsyx4Norq6H8HfLRPUTx28FsC
yBdLYR/Xycybf1LOH5nuy05b8KYzBIZ812qN77GNKD7fk0XIlQZxQYGz10eFMQao
mT9MsbXUVUNLHl5oesoQl7BY7eQm+Tik9celX8oJzv7N+gx3n7EcZCiEFkEZWRPE
oMFrrtXluILHU5AE5sEVYeHCstk6H4OY6kivgQomCqcX0yLQaAgv4K+ffsZlvYeq
z+5Zap9kAIH+8/YycrYpG7E+rdRnvAPEgVmKYQewb3m2hU+W0/znQXo+jPN7gnx6
I9HwPyeZjQka8X4u4wz51NS8mCkIwOhr3HGNFYabdAhji1IRzwR6erfP75tTezPW
S19J9uNidCTCI+9BY5H7nzg8/iMUK8Mb1cXpu1dbyt8Y4I7MaFAQq/leDU337ex4
i9RoRVBY/b/jJENcf/bPjFTDHA+iOikAvlnWYyLbP4RrO5tN1GYS4WU/e300X9cC
E5krmA23dYwqnNiFAdGGlyxADRmVAiLX9/5NmCP0aG0AI6UGtoExKTESBizXZsxF
hrZSFDkgC+NYgRT2+JuZO/k5HYw2xrxTUhP2GFoJddyNJRpUmCtNISn4LS/BOkKd
cjisJoRLzOMumNdTCdXiT2qehPypcduksLiSL5kjSCA3cuiobJjtjUJJ9e3oAf4+
7psTZyrriNb6PRz2Uzr1Lv2N3XZIlB8I/dAMS12CMQwBb0CWShPUTwBnUtU8ZY53
Zj4asiujbYpsd3We69p2pNq5GjZKzIe9PKILkKrKw4ERKCz1QWRGbr8SjZvRRKA2
qO9EGs7MxdYEkVWBM4fzF3Jt5wsyraCu0j+ZUJJcuAX/OGg1qO8S74tjrOFV7Amy
A3kgq+R0djRXzhZza+c/jx1f/wA78V4Wv1qBpUeyQBUnTGMLyPADDkmZ103UGSlm
/9P7tzjGcZjJQfKvn+cLFDU959+N111AVT4BLkTJGkBtFqCjFL3xBJUlsUojZbzP
ClEeUnU24Q4IPep5OaqTXXiEj2y4Ofarfes2TfeKZsrc6b9UaXdnce7eRY4/8PSg
DAssP9GnzIbkIlwORxxqSYVnasiuDZTvSRDXN/HJVdFv7lcNvuWkqg75S5XA6kWN
QioAt4i7nb/aLFcbomaNjxwTKm5g3HPGK+KPqJgteuSt2U1ZTW0AEc9C7s3CdMsf
2F0et+Ol+ZUuSti2nk7QM84nXg9z5uL0ZyanKZWBf4XWMyQrv1hdHufvP5vJR/3V
/k/QWKQE2C0XHKr5UekCaU8Lk1cf1FRVuqXhp63T4SGzMgkLGFWncjX0G6Zo7btH
qdDcZQm6tdU9cIy9TqKFhEICV++TS5yy/Tkjcjma6NUMTxG5BbYGk1sc1M1TJD7Y
TAA7MMyw11JVqj++36XFtZQuXXtUJMBpYTckDLpW9arczHjRRrPiK0caJaLrDDZu
GWPlOgjgJhl3JsQi6MYz9CtHvZJ0ksruwBiOUba3ABPUa89qhIOk0XsHoxteJaum
c4xnZUvhTZip3SDKxpTFiaVWSRRj17V9DSe2bSPF31jYW3xBbMd9dgj3kNgAtg8c
W7f1aO1U5NGzqzSKX4keC/CNvACtREGC20I7EmhIvTMdGcidRaYk/ffmQSTMAZ6F
INIdqU7YpMeYdqlHOw7aIjb8cA6r1NABrumE51VGk61mleoM2GEUEOzyXcmzxNwE
ALP/mnon91EZ2f0QqmR4d4oP8q2eALhGr+PGuwkW0yzWSbGQKcSxB+tkEW2DGaX1
Ny9KGKmPlBjBO3KLQp9kd//Rt/Uc0jhpD0EIsikp6qQOd7KRFxcBNlgG12TEE06Y
laX9rlsuqng/H7fQCY/5QfX610haLlOGhid5TthECAmIY67kERrEa45gEIXh/RDK
MWqn4wf7XCiy3wCmLfumUZQe+odLSLUbCT9uyTdbm4fqxdxahOH3uablFVTaIiPM
yXa6LSGu+SqHkDcniIlBgNwdft1MhoDA4mx4T3tMiDwaoOnQ3w6w+s8JWNtikPjm
cA8qKR//Suv38NiECT3JzuX2UGTlnJJtYlQXrTujdPcxbEnFhxKu/UEWdpdo+0ZT
JVhsz2JbpuQaKfEKUHQuSKrD3ljoHZg1e+EQcmEDoa572LXAs279jFLMhk9QcwL2
NEZOdTTPa1OyEKbs+jDTDZMV7N9gi+ZNtgFBhSdtCpB473AWC/RmPIZxRZD0aKbs
B+XFTxm4ddi18bver+i7UWWKFwH7FDL8nVEjO/urjNESPIe17CucnPSmQecXNJqD
deeluV047nRoExLekM1owDLxGpwBaPKYPpWwTB9zuvZFMdUT6fA6FP890RJgXGAp
h6A0sPRuwrAkViCOq4YavP5apmqNn4FqcVgIx/JFNjIES07iPNB6WXIqHUiXTp8M
oFZdTjulVeWBFdhPABRwQueTlz0Z19zlVVztRpLzkSESe0Opd9E/rq72mE2tU/LK
yhgm+wE2IvFQNtTYhHhIacEuJ5RlYQrPymtOBUb8yv4MTS2QHGfLQPRJN8VKQBzk
UYRkqIWfvzurOSPLc7vP23z068gYtN/kcyKFhE5rOFiXUmPE5fyXZkiAuS3eI7G3
fNehscW0hqninxIpHfmz7vU+GJJZkMf5PpTGbePDTZMufy5MU7O18rNp6MaFLnAd
dUP2yCY1PXIAi9457RVWVyzh6AI8XFehzmu1VQQSuonHaa33A40qoW9aQzRQKI/d
YEH0Crekz5LpAsYJarxCZDlUndBxPA6+lG+vaXjAyJ+Ru5wzk4BhAegpxn0HFXPI
uoZxltg6EcS/Zhag1ZMtM7LRj+9DoJ89IXXJ/sHeS4JZOXVhIZJzQuP4bCpkhxkx
DaxdDPclCYj0pu/4KVJiZqhRASkXvGwTupzoAEWoRQMqi0T/uO6CjRRcYJg/L4cD
+7WJb5zXzluB8zTtPONA0fUvnJG168f2VT1mawTSXjR3q+HFSM7P4zZlYU8jI7x+
/2QP3jiso7RZIU3zgqasvuxs2eXcXhgIR8+bQGOR+gXjRmFTBK/CJJcbnBX22FEZ
qH1Q1hGKoVBhryZE9acCgetZnGzBQxajb6amLDHhV+mkR/gP78R0SMMpvnZmIuPN
YjzKm8CuEF8+z1NX3yHpY7zfGFRA0+VuB0qqpYI20bGnaoKmu8lFK8AUcE0l7LG+
Xg54wV/pHfxBhj4vlspO6ZtMpMweA888DCoJ+hcYxIPwStCCj5qF217fmOyIYsPY
+00W/xrYmUwXbjtTEzQG39H5Gk8d2raW2mARdnclef/aHlLDcrKEXDw+9F91Yxqv
q0DsTeyoLVLs1KmeKLN8cY6HhHZd2B6IAb97i5T00hmhlJqsBD9AB2WURH6CQ3qY
rCzfe1B60I8Onnmpvoay5Smj8lYab5Lucuyn6s7clrsDY002a/mwOWvtLrRMneUw
csZya6PPD6fPmuxhGSeujGPEF0bzjfFWcmdl/p97CsRNOhg05mSBeJR4iWhr+HLw
lwg+tq52LXV+bveK/QwBUh4nh2DnMNy2eUq39sJjnv0acLeL9Yk8/gmMPJsUCAh+
Ji4ludSSIOsiFYLoEAcpPC0zqEPL+uUDavX94BGwCzyCZbkk2H/7nBnHSjIA9+cT
TaW+Ce0pBCcbZ77ffR4yPmyxyGUFiF2b74A6YA9wMArPE8IRsETAj9HOOHZPTboy
n5+lblGOAL4PZT2FcOGJKi5MUP8nmrv9U+XiZSCUqPXYzvBsb5/hf88eFtl1zehR
50/zOoRNx97qGZOeBF8ei/trWykTybTf9lPZULS8qA7ndu/WCAt/aMgBRvNBU9bC
pmAmPMhdXKa/5HBMiM/hcEKBH4BhULzuaVDsIgnaz89E68gjdgELZVYQsvcHzjnt
kFDT5G/N54UXzFNMNNrdw0NgVh7CQ20MlnukgYU5o2tjh4HkHqGzu4/mef7+kMVm
7BKnY/9SeRhfCSuuXXKHIj7wB1N0wAPhf4UfxYs5VD67EuwaBCBKIrIUpEEh9Iif
iua/xpiLEZWaYyu7ZQc+cB+6J6GgNCCzpINTCpo18/Z4whhMO38VPrkp9v6TlGpv
IYbaL+BVtaZV4Q0xzwmM+Xwj6Ipp2aRUKhRcw7B2xgVWbBb349uGgVQbM2KQlASf
QZNMmDNtPrxuz/kp5sSXvDq7D824E5bKXrsiQoToNe9xHpa2zpMytufIhWdo+IYr
4cyBvJbXs314KsY8MzPuWQYf2nupxXbwK4luMPSUi+KaJfQ1YDJY3rNIUlqn7T3E
aEaIrhTRzFgRpBZ4KFHW2pLQNPVx7DESzxf4U7h5czqH9ZsIlh+caDc75hBkv7wQ
5XtCYza/GwwFmyPUGjduetC+ENJPAn0ulgRz65IaltZNvvZLrIFU8dm+KVvw9q9l
0dZKOPtaqhcwmmv+uKHxhjZiP+enamIIEYB170/2+fHn6LRkhSr86s16BGGX7cE9
K0Qg/b8UynJOTtDBn7WjekhbjcbNTvFQhxBVYUiycycdIotVOqjHi1hSzv5Xt5+v
QOJafwmtdtLcCpAT78mHWX9TgRDQiHQSIwFf9Bqx4d8f+YjqNMYf/Sucwb7I8oaV
OnoRbyTy6R2w/Z3JgqkHR2o3vsh2gI5015hPHtpttVLazMFeFnV4xVxGamUBkVTa
sp5zrFqpOCOzG1u94wF8GwJ9F96Q0rb7YriQOI7nhdiyZjA6ZjkpvhSwFLYFV//C
60I0dWEPBEHK8tEw/GW5ZWKwcMhiOraqMvGhaHPujuuk6kwCh+sTiOhuZfN8YTbn
2Z/w3C8IgJdjQSm88Hnkkqj+MVHIVF6uTSEPbzH7j2dTeHLptImp2BiuFunqvWC1
3dFeqFGDTnWQ1sa0CUWDKqotZIl2LyIoaeDbczj9JO2xqn7Kt7AoDKYfg6MipWhw
/ppvqi3oflJokgA1XeGyjy8nkc6ml6KdLBGVEZOCVO/Ngw+XlK7haoAAE/jHRQPM
3sQU4Jx54A1yzkTN9DSDFbuMxdorO7NY2BgXjIpTPomapjodC+1ruD8VhlLZ+Y0e
4ZkQt91h8mvibxuhDazENDZrrObju2iJn3KmW69MJuotnlYbJ19w6RRCg6UHKCA5
UA1eWiLr1bdJLmW6to9nl7n2XVPOiV3FxUqmVikunN8CfRiRtypsUigJmZC7+URO
vUWA7Y/3abaSh3wnZPrXFVangQWij9RUIie+zLFc8YD6BxgTe44YubYtlhu7D9Fi
KrENNWXZlQCM9FgtWqyx+O2kDG2VDPMeIzCCfBfdfy0rrsDWGXP+R1JiOJG03juj
HUEhWpNCQGc7MVolW2O3sCREMpjsy5a6Zd7bSWBloxRPN6xAB3l3W8wh83pYz0/z
1ddwxa0oepUkuoxlKtKNcVsVe3/Dp+GWll3gnkPushJb4sGxjqYnEh4uu1x5Rk+S
uc3dSiqz3UUpwRlpzFVz/ZeCqbnq9pwqjbcyLWl0+JsWnY4IXsgAQdcr/ipwdHc7
a6LUPA/pFj1ookYEr7dqfPfU3Lk+6ZtvfyRk5uKkL6bHpL02lIAfeW5xaPQwZhvp
tX/6h7n3jTWX5hm3NIAeK7mp29ok8OMGKQ+soCsJxc54MFpLVTq0fTFH9GwFueZW
eQ4hf5imEMDwgPnfRKHBe78kB2ScNvRAo89Rq9FSEGGP87bKAzxfydQnUtRzF8Jj
Z4R0yfrNl8lpRfAEiQ+bzVqj9zLVwjZHlKYsdhPEhV5MQ75Z5uTpa9xVrWuv6At+
s1jTxwMFPazM4G9ANZ1KY5/Q6e1hrLdCFXX7tgcUbyWaB62w/dX9j9kPTMZ/0Rx2
mn+I66h0shG57fWstoxL1pNYk856x2J0/EC14yA619m0jHfhbzZPVXF57vZZ6h8e
aVAQ44ieQMhNClEiwK+FqyIprcA8iL3vf1uJxqUiWtcwdZByUaeeBUHvggLMKomQ
y7PUOp5NB37+xiy+6pEw6lei0BH+PyODco8XvbxNLqJVRT8F6+q/mXmhtc8FStd/
2J10Dq4bubKmPIxKiVL1qh8nbq90Ltgw/0ndsTC4THQE5BAjiDZNI9CR5RyevsDB
L/VLR7fW2iEgVpEAqGC+IjVjgykQbYH55AkZgGmhlQRjV9Bo7voRJ4ObPk5fNY7w
OO0T0t+U62PrGCd+ZvmvUDBOdpgscS0FOKoTixc6A3cdadUYlSxU6u7YvWxd417C
IAOVKj8RHd5DAGmEkhehU2uTG3fztu/JQsB4F4WhmL5lue+v6yeR4n5Pec+2TO0M
TcsrkOEaUCZwohh7cNqcMWfaH164LALufdCd7V2QRbmcoDiMci/eq6rxKMfHb6EE
nbAihvHNHJOh86xs24MfN5jyaw8uGHqSHurf93vpahDNHE4H2xjdwyLA+9pm7VTh
wpY8uyCDhptUko0AFR/8GQqSQzxsqTS9wvDvAS8wE946l3bytGD8fadWL3hzIQsM
n3S2ysn8elALDBrM9nhY4SPk3iwdF4ioHEBCWEUIxTioyBbPampLeOy3VyVMxmCl
cU2YN7e/IASSehfhurwpLqsJP4dIAOv9+LS015GpmpvM8zb5KOT6iiEkUKxQd+rb
Ow7bz5mg0h44ShhNaODfOL+DB3I55RYxjQHC7pplloMXv9sjNmuytfGH2a/V+/aZ
kp5tnH988ljVvqF48QB8csPSus9FQySwrhVA+cUCypaR1ZoHkVZKga2Er/w0QeOd
3ga3FYmX79ue7cD/oOBLlX9TaD3mo7tFCntq5IhYcfrZzD7UgUI1el2g30AJhkOt
rmAB87ItYdOZtxet1/54ZxYAox5a4h+C2G0E4VsM3uk6c6262J3NNN0kZPzgUfLz
ilBrqoTO850jioLHnYqm8g9Uu+TLBgRhrVsfnd40gB3tdwGgjKdeyors/P8iG3AE
QIQ0Q5ag0lGvyomKDUvcsss+lsNC8XdAou3bKahdZ1fDqO8vtnIj8ZInNJLH1GRy
Dmh4ldndwDMaUDXQHPybBdIW+s+MgqfvniD349zXwQKaaLFBwkGZe+GQn/R5/fX3
xfaT5leaZnr2t4UOtS9vlz3KFJIT1BcqpI4T4mR3UlPu6BZOWNknrFquvgPMltTE
hdKes/t6Uxgw94LPRYEln8CGFkU8J2k2IsMENzYCmA6+qMPtXKzKF9uIr40q8M/X
ujwlztGTYDkbdMoI3xYSCBuI7E2sbczW//nbT3q66PCWDYdORfk1z5Hd+BSZrK0y
PLlSxZK4NwsCTlycyWguTIPLfJs097pL8UqdnRrGHF7i4FL3mSZEthbdwfW3hzrI
Pzrn5JA7YCeZ/zDKohHbP2SbFNinOdr1UvWyK7LIuLJRyOU+tz/wfiN+5+E6e6Ss
oyrFQD//UDC4FSvHEVHJOwXC1Kh39rPzpDdMXZBSTUhajBphdi62WuajgzfNrIBK
dASU4HLatnBy/w1Wg9tCi7Zzul8M9E8KHx3DWPQIVUjYtOPdgQ+rkfinjC/XH+Gs
GBe9JcC/ItcexTdAwxVXzBg6Na6LlpLWyQXm2H70A9xMIuBzpxBymWl6w7FTg91K
9yQ2udsTLDYldzRYGex1zdah9wxlQdQ3qFKvmLfiqv7dnE0/Jx/OcSC0DrQ4Msaa
iYll7vbc/uEp59+/Qdhi2uLeToZQr+WXWZeuQA+OqlZUMTk8fEfc4bPaMxCAwyuN
tBuL/F7JwVSDtl4Xr3Apcv/J0xks/AXKfL7rIVLL6rqP4Vaicg0UyLvybpZIB/Oc
YIDzzBwAXRmSrhlMwjKuIZmmf7Iz6T5LJotUeNTUmnFvaFJs3fO5zlYb0HQaq5qo
EdXbGCUylCLdR7FyNrnHxDVlff1f4EUAq0O+P8U9IThj+w1opmn9d864wgvBIFoh
oZio6nPY5qOeRlkfIvjztlOksmKL9qxiWfba6+Ig3GEmcMhZDmtwWsx4vzpQMH7z
pv7l+juVAbioclJax1ZEY2MzHZcAbX1roRXzNVKu5haJ/mqYlGxBHogFmaWrVHQr
qXc00aAzq0eSAYqUKUd2PIB46xh7Rm4XDKBUcOD6cNVCNSJB9p7FdgQ8XCa9jhpS
dwefs9XFev33+OG0p2Pnb0XE8T95hUwwvFqcEjKQBAkBX87iqwZ0knTjb79BgfWi
H07hdc82qYMQASgmpkEe4zwZjqq0+JKgUY6HbVgXS6QUJmhKh59l/2rmMk6groyv
WcfWjyOrSblx5EYsr6s8HklYg3v7+/NyTy1/dDVkN0R8syy+I9RTo9TmJU0LPZzr
d7q3ZSw8zqtZKCBaaqI7WYqfy9w/gYgLcv79FUT6QDYW60S6tMl+oQ+rb6/GaYak
pkpp48YULGkBPyds4P1npAzwY1pU080KKbPd4P2mxxatDiVj8d456eX1mz9o7XSs
Ynkn3MAMV2nOXv+PVa2atU0E1qb4Evm+AY6BsU4ogF3NEyrEbUFuWMbFO4pVggNV
Cf6lgJ2zakNE9T0YfdvSAeDQSUZ4jnaRO2Q8v9vNoxh3fI/fXAKdYmzJflrENxb+
GZB2mmqf8z9BdJnz7aB/LkUVapDLeGZJz0yw5otmcKCchKgImCioCyt1dQy26kNy
cDuACL0tZ3Up0+eC8rDeHT4qTZG34kJ0XuFKztvMH/GQUN3uxbvUvknbar283ocH
Nj40ZRhNNsGA3njUrbJ8kB4zjkISRxxAerJZ8irpbrCb5Du360KS+m9TJ4snoxFW
BQj4bD/8Say5QHX1CgeO29KDygNld6UHddoMN5kqgAmXtay3DZgPIU5FKjkgMxRI
GkILG4Xp7lraVPVu/o81HECuEOYDQwZ8VpdIe7evSPHMEJBrh9j2YH23DbtPq83H
1FEQOCVoDI4d3nK2jUwjEx4SwAZQ/26xbyFiITb9ma/oWS8rN/Xn4uflI1A66SsV
xIb8RqbJY4g9yBxOT+Ie6NFSUvv06s0zD/rdDQJouuDnKdiXZxnLn12nwcl/Hn5E
e7gCpPwK5pN0wGoWotq8HROp84ITVVP9As0Fsk8zpK+HoJGw4Nk0w4p6WkfkXKNn
ORw86nqEDJ6GyIU0RpBNEwjkmj50X8hlbLetKKeWcXhz+EEkAFVPyQrUPffZx020
AhRp0nz9b1izzz//BqjyOexjwz+piGdKdfKfTCJHK8i2dUEA091ie1wy+4VXdPiD
AwS8qiwKFptwXUBZpWnVr+LJH5TK2/eJd2P35NKw/Lf1vW9uWba0UItAAjMGFBU5
CwSQypfLDJ1mhHXvEkuOLdRRYz3k3fVZBaWqbnfIz+u4WUYBJKHl9kmiqnJtXJpO
Nmiq51Jdr63QOs7Dimz8qoZrAfUMyCCuoQI2QtZ0g3bMdg7RdJPnz38BGD1jrTf4
uZrpCp6MAq0Jgj3oBKwHnD7BeSu6rmMmAko3GYWwPvNedxJtT7m5XIyCorjsrlPI
XDn0+/jxoQ3yISoOksDt+ZfpKMBW2D7zscpJjbP5iftbIVqLyNfeVq9IlRzQ/d6d
p8wdi1g5sgVrRziBsmFHqp1l6s6AqwEvUH1q0cclpXYLSqj8iEIaN49pwxiiWMbY
wJmSnSPMd6pCZncl9seMmFR5/LHqB7MacSeMG9utO1Uw2S3auNyU1c5qT73WWFMA
/VULG+ylgqj+a3dWKJLHsS+52S6tJfwiRHWoCm/wfpyKDAfx9cpKnlq2BxDtI47A
JlbKsrcUJ791JP2qI8o/q2fzGwbQlK/qy2LpQfPBVUDXiGVe9PEsMOiKxoCW+OUI
eOGgKbqbDkXn79Cn5U7WjXI04VlVZlRc89Iyz7W8kTtcJtHERyl84zi7zKNKz7tr
YzEE7IZoLlhoEXjPOVPsKL0fy3xt6UXp+r8VWkRWh5cZKZYtCz40uUg4Yz3NYviQ
j6381jOULWy6vlAuAoC1Z4bXAU6KHprluCyrJTSTl7xS3rrsExgLeoryr614XjJo
P/4LpGXPMfg4LKjsY/BblCAv3AoeecSNGP0SKZFmx502jmzvJgiwKYmRkAGn8RvU
fskKeOAiCvom1X5PPJsR1AvSdPTYub2JUjV+XPuD0d/+vyOTxFn8HH/qStPGmRFE
nxY0/cE7zoAYQNaCw9N0xCy85xn72AvEi3HaI0GuSYy892mQ7CxokBk4UzwhgOZp
MuDl47OsYLkDsUfetWKKyPevNL3x3zPJGplmtynRdw6v5WAgMvoAEYBvMRhCEMe+
eMTNsxK6LcaWvehrNRDMhjtxlLSOIZkBfPi2V23gNt5S2Yi2bjexrfBGVDBCVpWQ
ughwx1He4DmkU2Ew6F1/Pv8tdw7sJG1Yo4BWRPSufEALdQKOuxShEewlyOtvB8J1
LM4NgrOe8AMdQDP/eh5xWB/Oc+9n66y4GiEiuRF+qYyIMudmDj7oyz++OF35jywd
et8KoTMevDKq/DN3Xu0bsfSLPVFDGPYfqGha876MWeWp/wKBZgwVG3/EXZ5bh6fG
YuIrDOg5X37AqFYXw2mKB/ztX0ckbehBJP8U00ZWHhdYTG5DoAE2BzJHWisi3Ors
fVJnxWHL+7ZlcdgZH+Nsb4rnVArl0lsIbKSwBTlnKRFpo+uvQm/5vN7QZ71bp6ok
mljCJIhTA1I4EHV8dpcnkSGJP+7BWWQdzMjVRbSNQAFKSGFrSLcBk1DjmGO6lmRD
xH5wBXIU9YW3SKPilGczP+H4SXW4s8B/44X+phQYaCjsnNCEccV1baX1VHpaNxTJ
isW6gIDtiBXAXC0CzrM7jH3F+mRpm76lcyISS+XNPyKvHATNp0bf9S5WwHeVqhRG
N5PQK4C3Mwbkhn1kW3BtLnQb8FZPoX6mbh+2M7jI+Xrjt4i+BO1XLtWRunwnzJup
ILn+ZQ+PI8XaZeb3/ziW27UDKqjYVWhBj8YtdOm/5mvQUtckOHT2zRuBRKWXcMl4
6XAleo5TagLey+GAyJ9CXB65PQ2PAA0R0LYG+ZNS9VNt3JiBhX6e+ZPeD1GiYsrO
/dgaJtGXjh2NtXV0pp8CB0Pq7IKqAl2fsmaYVabezUYWyx4hDT1H/6/0ABwyPgbt
Fgzby1nLrMeJxhGPUoCNJGD7OnpFmWn8ph9p0Q6RoapGpxBDjv4Be9ysxbHt6bGD
dsjhMfD6gJxpLruRXFwr4+14Ae0Ne+spVJyFtvy74ljqWq+PFrXro0B8F28ntNyW
TBkP8vdYPjGsboWHzLAnUQkywNRHYQca4FhzDjHt6BLjqj+Sli/thJX5WRkoe5k5
R0SeZtGnP6mtWM+rm1C6hkFxkRGBpiw4A3Owbl269Ud9xM6qHVcm7Rc+44E3gXWd
xAEsZDMcLDGRA8w4lr/wMl/zBMZ33+PTFc8zpxKziHni+9J8yDwA8g4hWKxYEc0N
dFvU2dj0UsYm42GqRb0mVkV0IGB+aRiv9spp3bKqJ7m3CqU3aSuC8ux/16Vkl6in
Es/lpuM5ZRnKfhlHSVH+ZWovfNgKZGjE7pX33D2bm/iphXO3B9IgTw5S1EObkRkP
dZ2KTeYMGrIxSwEK0yXlellWCthhSisWSprYmZmF84c3YiqH3FwkP30MmAGS+xlU
L6FkHqeP9W3ry/JkkNHTN7v1FW8i8O0aU5q4z3pZTNo3LSpuQX2EK0K4gFK+mYrU
fo3rbyxqoGuDYe4F4m4BgUrB1D1siobrncPKz0zwzgCP5sCmP8RaDLCVw1qdsOER
YievjcZgeLQQmOw7JtRBeQ1t/R7z7m9Nc7vnQ2msiZDr9WLFSGpvvXMY1tRhrXUf
vGvoV8jlONdQcA1pBYdpCqsT9krz3i71vDc6YuFds+vjD9vW7z8EuZ2gMiHsIo5q
iJOtHKPqYNyU2EQhg6fy3TEjKCV6TQm0vM43RqFl2Feu3q8Ipi54Nukh08jWMGiY
/eI4JgMYzIefOhPEsCdttKt6lTFS1ZUX8i2y55MkuXhSQyRSzZsppVimeAqoPNev
FTn9nX/2hh0MUzKHM9dnY8n0nh258HxajW1idte5KNGkBb16pPevovzEEhRBx+Xm
9aIhvn5YuRrwWvKkMZJSFRPlkI+Oenr5WYsz8NphIZgwmSUbgcimuQz0SXMpN8AW
sXsECtHTEf/osdafNh9ocZkagyVql5ogYYAc/ypJhKo9HBttNSLj54JGChh0Mdpv
ZhM8sZgmDSDo0Mi+/r4CrneaY2kl5j9x64RREYiOqKFOeKDO/IxUCGcRpgt75QY6
GRyogkVguk7nr/5T+rYrVCAuwv1hxJcyYXkycqnYxTpl03bXmrafeZJNE8UMLd36
03lPHdOEY9hKcreOXhVQp8SwaMaN1s8BDQkagsQKS/cO9uwyRN14NbekVfHY0ide
YODxgtYVuUtGEL47eyzzjlJAS8t4Hl5aRkfiYD+MXADeJ8SiHbe5y/WZdwbLw3IY
eBfaGZVn57Zsslkg7ec2D4VOt94icbCmKpjzO1jLRXtFGvwhi6ocN48E+JIimEX2
10z5O01Q2e6Y3vy2klNmLWnIhfSO4WglRhZnEvk7oGk6uwbkxKgnEjQmeepi/lTp
1A7MfnzqGbIUt3aErcWA9xQdvTaDQ8hX3oMX17CyQShvB1Sls59LdZvydVpK+U0/
yT0FDldNKG+zVUAxv4xC2K8+Qdgz9ExYwZR7BEj33JlG0MM33z3pNy6OX76wXX7h
fvz0aRec0ejpLDrdi/ERo8VynNTXqNKgMKzBm/YPUucLQhFj9RpPxXJxRpu+m7AW
UjN28KF53z0EPUJ86X6pHxeGSG2wa8UCnQ5cEPLgo4ujyYfvAtp0Ob1Bc9b+4NfF
GuZrqo2RoPfCPwE6pKDWAls52xtfAZNEWRiqTvBODDUZmYdDkh3dwXGD/11NZ3EG
uYfKd+7sLYK9atadDoNw6wyI/Hc55W4Gs6gYlNblja6Ubi9/nHSnSm8IIHwBKojs
aVUvsVPijwm85NBic9uLUoAJ9JDorQTOuQ+JbSflmNG/hyE5cj29nWmeSQKxVc6N
hkxKbWIMkKkW44rktBpTyk0EZJsN6RSqbxy5IdQmfX2pzH+D+wDJDbocTbAdi1Ud
/2x5DooNhNR97ek3487pDK0mV/MySGkUrcqS+MX8qKjdd0YG0MB+R4fE6i2DXlnM
xHcIPxCk5izcjI8SU/UQCLplSSzC3lidha8CuO5q/xB1eybvYkrjDSFPULh5C5r8
8eQl3L8AGYEf3rz916B7F4wRAVdnmg8WqqGkP6OJAFue5xdnasuEfVV9/F4SGCIP
cDD62PC/L4iWoP0SDaqaSgh1TCCdOBXJC26Dc3JcIhEfuT+NXqPExb1Yb8BYJN3G
MAT7wBVzOMdcKrETD3Yh7s5z42EBvnsBroE9KexG949MyyBPVHQ+YR/UyCyIaMAE
NFTvzUODpVXE6vC6lzEwaaFAIgEoiQio6G+/0XafQVyIRnfNvA3cnTqKeYFZxygY
mD8yqQ2Qk+T2F3v2s0R+SFmKXIeZaNZdSA6wcs++5fLAHTuMdOSPIO858aXbTGc/
XYkF9rHwVL54uOfuLp5hm+1O4VgB9wHEp12xbfY/d6f2v8kPbP7fB/GZ7CSoSV/5
khtLn+O5B8fZuQ7+QgaOJS4IQmp9ttVDrsjrsbi/SfxvkZ8ecDPDI8qg0mJfihy3
WTXwwbHwuPExZM1b0RbzQIrU/OYJab8aqmgiwbGYYXCyGgD2fBFoehsA2oJNBj7e
qL3T2/Ojdmudm0dUfohWeyycAqJ6DrbKWGDN1MUuxkF9PrGsr8Eo/7bMzSJhMtvX
lzBLs17FIVU1Cu+9WLL+ANpEnDWsE1ywWVM1pMohv5QL9WupL+U+tC71lfv5L/Hg
zGo28EymL3NuyaVvG54/Qp3xt7vexEu3S7+5e3xIAqMQrJeQLGDvkkyl9hbQo1Gw
KkFtmaDcqGMmunvMcZf3uh2sPK8buXNKTElbLyH7JM1Shz1jBxZdLktB9gxZuoE6
NEvc1zTpqxgZTl0tSJ+Mh9yGdXni3LaHJ4eI1c5Rc9W4xfD3QCgKz5pCEZvMkHVm
qI90fb+W/iF/oplug91nt9ntjusx9Mo/DiCqWLymPJFuaNQf2IlxpOsWFiRwfgiQ
jKP+M0C4bCgSaPdASPWFUnQreq7qSORQBWL6K9ubimj9HSyQfxP1grU3U3mQB6Bv
v/eTtCGGgQDh/lHzKh6+USew8Cd7ZBT+NnS/exK00cb5IxLc4EfdRY56rkamxcga
W3rRIbPgSrHGGCTxJUhpmbdVNynd8Ok7srf9KGkb2/ZohPG7++Ulz9yA+QMK4UHB
Vjnr2Aq4eexkNlg8P1CJthfoc1HCFkF2rUIunqzytmyyH9gEvH9rV3u+IRitagPU
HUpDYzOgD9lo1ORk+dAxHbT0njVJdpSGMJZ4njKXnx0MFVJmSJzzQZ8HHVt28ZQJ
ibzsN7rUlJ48/D3KzZH20Q7V0HfvuKjUE2exLZNFDkpQUwCNG7rPOnT2go08AiHN
CC1SMmDFOakQFu1YhhfP7TgtQfMG85Ud+rrGZFsxrwiyrCCVVI4KuU/cQI/HkBKb
xogRthY9j2d84HmsHFBvR1KNTHhrehwQq/VQAm106dmrZ8J2IM4FEtnqzIUHZ6pM
26DQv9BT6iyQnX2W7rbgmjqP5xB+XZVzCdI+Dw73gB734vHIytYDzjepsPA6RwTA
ANF23pCcW7Yl3LmpoZ91RwIyqijJ32itbGHjbQdEHO88hmmle8nn/FUeAwh/kkLn
lvGadCFF+9/Mg960uiVjfg6c4BoGWH9l40COAPeRMR3tRZDQ+3svlnzEqxNiBjOQ
sZbtijrj1K86gMJcXkusySpvsVb2lv6JuMEpl+tD0UihX93pgjJTGTYXBy3dzMBt
Xj4PFUd9bZgdCHU5fgZrbwDdU1UF3UmN+vaWQACh5uYcmiAM3fSyyPpHDgd7qHXx
LuEVznZP2HU+Ptwoey75Q9+Gmt/JRrSWmfh7CzXCu5yCEWuhbIIc0tN02NahxRGv
g9NddRGkuDT4pbGcYcBiqUx5aTy1x/Hv1xMQHgVhK/2vAoTIpZ0DO9Y0Xuljca4R
AZ5+W+x9u1nViSSCUUcnybNkE4V4E/NEZzfzposI81EWaWNqoaCKd93V+14nhEt9
p/O0UiO9IYpL7+F9lZRguk4kcfV0OFj6GD87YjJpFTOwJcer0RwgspsSBIIehds7
YVJKdjDPlviVGRbUC0+LmHORwIcHuNCbodDRnNaIw/7K9tYNPeO+u+yExqdvKt/g
HrUfNgYNGaiDBhSjKrdwZGypjT6aequ7iSIzQSGRRI0U1IaIRXSpyO/2L3iLozDW
8LMNh3jBhd94tFpuQX37b2nKSoNxBXC8HuNZVTjHkNMncdZphgJqGJQegGkAKdoo
tYuem0BHyNqdps49/zos1o9UxGtWqxWtYhnPEISgTqeqNHQJN4cr1yC4tta0AMKd
0mIKlGEBnHyjbYL1BadWCd/mhl96hsfb7gYXTitIYTvnbKfty3ZuXFpKHWQGqXrU
IzCFTreUFVN5QkzJcUOCGze6IabPs6WyuFh1QvQerY8/itHJglnaVzEmFc4NyC8f
49PCwnEnaBkd4gn9GUkzLOi0Ajj7REWG2WHoH2cElpt84xmtzCE9dAixASOFk7wV
8CAuU+ECYwONaNPhjRhs4QDF4tnfxlLWn97P5be3WRxYO13mq+gY4A3R34uJWLJc
cOmr3mL+RzoIuPTCUnZCfNYJRZce9pAOqXSsqQS+9Hrb2/UGtaWQ6qiVeoUGQ+B/
8rUM4t97L/hGK+pxO8x1S8qfFNo7KpZgB32Cxcm/WFItvui1DAHxCywvU5tLWsNV
5+IytXub9F6kyPgOyxreWK2g8ZLkXc4hEpbz6q2b/DNLPotuo2xPS67nixETAfbC
5kROSLAhcgq5OsPViF4ohublYOSHO3QX1VoG75FpFyr4/UJ5pQneg0Svxo3RdUOz
rTOFww6zos+JDRnZNZuSKJJRLN9h0iqmQhTtOfU2ZUrWkHQncqhQD2qeEYV//L+k
8nolGvx/ew47GSU19c5PFhPy22fWJ5uBNb5tjjVi20XtCko/2tFE2Ipub4Cav7Sm
IS+rLw/8uQiy7q1CPdieXVpWXILYyCKzmMg0w6rR5zrVJyF/KJ1YrXpSOXygnMYc
zV/q6+b+Cx6Y+U+3l7n+0EXxO363iwPiDNe3kSC6tn6y4PolCWSCN9DT6H8DgDlR
A5jFVy3f36K+PVm4mgwQm/yN6HawIBgKCT4Ap6IKnuvegJRh9yDw+TTFke5F/UnM
ga3j69DHNXEpsJL6e+Pz4AHj87SEakR4EVxNgmZhMyE0Jdi9/lelpCjh/xn186et
YenhTsoOUmHo8T03HPy/p2QtfUKjkdYQ58Z+0BFyG2GMzxOWXziDNoAASWkLR0CI
JTLQZd3G4XqPdJSya7o4Og9mJE0kTHjgllRG48W8rhMrt0E6XX/qyKTm7pptPj8d
Tqi+sPl53TlSA+lRgdDeT87RdZ/ixiDh+FZxkENgEO+fkLXswBtHIHiKCAXnWdxg
WRn291lziqUJ3HBo0VS7ogQ9CnChsd2wLexn7qIGncyYfDjeTjw7mPKc3otXu+ND
8NA0fiQQAASVzBgnkLiCoR/htWlzlZOqKdpVc0MKyfo9klYfbtfYeKUNkoeA3CPM
7TV4YHoif2w/+wqhAv+sRiGbr8hLsZnn6ur+xjvAQWofjnUU5qpW2dIi8EUs3iq9
ee3uBQ5UhC7Q5mMZlD1k7ON7EQ3QyJiCkXSqSBcb0KfYAQkYve0qeW74fvqTAhhN
MVVlWVzWY7JVc/8OGexlk4AlW1UqU0ohHblRFfNVRTLh2gr4DSBwjQpn/SIcIzqh
GcdUoQjXOsmV6MnThN1DmzITwiA8vSZD01O1XHIJtb/vb5yQgmUwDunpSf8TVpJ7
z+Lv/Vzq+X1mi8TWcW0vE7F2HdiRQ8mSNZ/X40G16KFi4p1UWElnDnNGQ/WRPmDD
3tmkuEGVZOJjwgvlCuvTCeCz1GL6wsFC1wvBKUXhl68iTTzsDDJxYUHrRVNVxxvR
MfCTgKsPKldYFIo2kYinje2gQOSDbT0BKgYNGYe7ln5bDbEhDlKyNtgV8NjTAYxb
o4E7CNFYFwNpIRNR5ZvvmXSAgTKztcCB+9MyrNDbAlolftJ4ZIN4dfFaH3GjZN4q
p63Vn5jR91V8YAXUmkA8w/cE7iWtehm8LTwPf84iHsZrEwiMA1mMhZa7kifD2of6
+aYBdPAdDDPX6b0Nyutn0y+xRmquPNjZzq/L/2h+SbfaZNmXbgove8T0sdmKEH8o
uVGMPT/gle5k/NW3VlJcnrY/crEmb3J3F+uFlCIK6bd328sXF9/EpZgKMBfohY5q
4TRUX4lHOr+HMf5AC36enqYMOPPvF8ux6qvg5bZxNnI2i0eCLBW57Nsv6L2lmQVX
+sLCw3y5D9o49WK0kJUc5m10Tb6FCiuD1XEjA8o+4S17klfscS4GSLXqXJf42MM5
NR6+poe5YA7gUY/NVgxQ27JYUBr8sWeXLcOKakVLqjQ8C46VzVE8aB7fx8mWzmHk
kFff1/XIFzsr3QLVTrNf0QmKKVAdhghLbhvAB0z99RAkbGTB4bN64rYK0Pkq6ubH
oqcZCGetE4/vOTuNO9FnKZbr6zkOv/ZzbJbTPBdC9WFsgTdsWmV3T8tFPesOjYRY
b+QTvmhcwya1l3YCMeVHpsTRn1tTVO07nc+XTzyCzVbb2iLH5BT2TLX0WPc1cJP+
0K32DuurP0hQif0PxsF3RqjVB+6RscFrdD8zSemliBOG1cpdMz5mAj7Sh9xNYucv
z5G2mKOSMGmhk5qtmrZQ6y3+A+v/w1nqkJjyVR4dRKybKHHCIDv30vRGkJXTb85j
/yf9dhwXkZ4Eb3JrLGTUOkb+HcLfYjyXMCphinKZ04S2/lGx7lrQlTEa6w0pCBwZ
KdmEiz4y+HUd8JYbTxwrxP4nbJ0gqolYj9851Bn6ZGbiMhzCzds3c3zibgbawAx0
TK78qnzeCI82WBfZG/gUYcSEL0qlqWF6NFk9agjuoN3e73bw/eUl46MgACOJdoOW
IVLxWb2qzagQgwTqhK9u75r5Bd3GgjnfHAs8G7Nb65OgUZLax/o44ANeHFNot5Ix
j6g5VcCrtYzihNpd3J3C04ZHMwwzuF9B7FXkI45/W4anwbw01wfRcR4MJzYVnAt4
I3IrPHRZaUzqCssmd2JlubZ4js8P+IjviTfyNDYVyOJG0JzrzNk+N7yZEOxQysRO
VciMSmGobFlnmIA0iYtWVYm5Y/liyML7KetIPbAyQ5MSyF8TFPMaOnLJNXDuOFVj
pZhx1cdxEC1Rt4XzA0bLWEaaeulrjNkLk4uC7XwfkessVKsW3l+W6dQZf6FiaIUr
RahDPxe4MSLM8BCAvO2YXl6qnTzz0LDiKURUxWIkPJt+RG7HZCJQZUiAKdeYcNNq
GWTbMZ850li+dm7ZxO8dWFCnkUQH+l28xCcuGkTYNDv3qIXDGKTjFGHYTuT0F4Fg
HAuhxoOmc39j/WIz+oDtnDdHX+6bJw1hAxVM08nHotl61IRHy2c6TUay0ghKGl7Z
I/TShBHAx8BWSMn1HX7pPKvxhIM/DmFHodKJuost4M6EMyI63wikenB+9i2MacPc
wpD2hEI597XbbvGIWVOq+FFSobuV3cbPFJVp9FqweTySr4S2wKhsyOfhxYedUCaw
q+YDIzWPk53tEjIqrXsiDW/C3wD0BRAwUGz4aT44m5rEO4ncMWTOYD1jZ+k8l9KT
8jm9rcNPQlzp04w9Lq+znl7/UrOzIoY39jDTIa7UDzU5ipCn/CQeZHbtAzmfb1L5
QRII/AgQICdUPqDzrXoyiEQsR3G0ZpdC4wNQxPddmC7mi28MXSS4oI61s9kjPL/M
JZwI3KP+ZC/bnhg0KAuEKw0u9Jv3PzP4zT5Sl70rsRAoYnjS+MxVJ/1kcNTFgA9M
jBuQ+JfGJv2BGhCBPgSu1b1Pm6eruUaOItiDrrAbwZGWafWz+0rttPvlOdcUHayD
TqC5w3hcPZ2Hj7zm23kF88R2v2xEARJydCdZJVPtZuAeIBhh9HYlLT3Posy/u+0I
NaWwk0UPHXbndBajhojKjEJrnh7AC+Ny46qRVE8M2QKbArb3+ImWs/JP7sqZCJvj
EnLuh/U7IH8tnkVk1Uvhrj8TANs1V9zxqMc0vLO43bINHoVB2mvOc38JrSHIzRYu
5mOS50l2ViwnesG14bc7excAyJ3tejaiPDKnmSnlvxQ9mf4IwcfZND9IoB//l+rl
8zus0c9WQaV/hvh6kFDOWY9UI5+H6HCYzttDS17y3UlIjNCmvL1LUAZmBODI6QbD
jCfKBoKJowIlvXeKqoh9QKOEY1qohSgJMr1WJcl+gF4ZS5TnIgA/oAfp1vUlaXB6
Lc8DFSjRdsd1aR6NOCg2RYsJ74gctfD8ZF1Vt1iQx0mhho942RCTrXZRa2dIkSSr
gp2334VJ0wfoI2K1X2/JAiRxNNl1IoVfZS7+IqAcoYBjj4YB37Qc0CUzYqX6hBW/
UR2zbjxtZ32Lb9f1jzM06HLa0h5gLu90Sqai/BJ/9uejm2tp0YwM9+LHHrReJCBM
/p6F1J4JUlPlSu5UApykaVSGLClsLhNImQKcuDK/RGrpVsNDey1+hZyeIaEim/Ny
SGjmZ7tDByVTmk4clWeB6U/QFjC909HSLzWsPWPMY4S9QkbSgTp22lo0tpi1q+mx
C1CjegWWqw1F0ahJ2v3EaAw344f5yfOElEXLkGSgou31ASnDr3DfCBiZTYN3vZIJ
ULgZPEwqpua2b5tRDG1ExHttbX37OnllSm8l9+aRkbP7tri1ga3pFAayTP+PoVnr
BzcutXxEJ7GUbBFz/ru8wGYmlL+a6twDS4pkGq7nNjtrkN5p0pk9QdnrrGq/8u5i
9WOxGdLqGt4Qp9K1W0+nmO97KjCD9BvJuCucUNlRFGCGx+qCP3eIWtl0t0yzGYTc
y3UBclWTFSS7e9+u4Vdcs7lTP5ojCV4zPwfaDOAEWli9caxRbsTewRPHQZkg45S4
AK4dtMKOW7jNMlaV27FxPvO/00LlLodts2KQomulHcYuymdb4/zottC+TOa4hSN9
O5sarBCVsmPkEWOXi9YmMLhVwaNUE3cs6PjLUwQBLjqhNTRh3CnVm1GaSUSlozh7
lI0iTduJlaqZpkHlrabf+FQyRXXZ2yhJfXLH2BUdATm1k00Q63BYxUStX5UWz1JS
4Z/Mpi/ZgiitBu8LoBweutwqfvECdTiuqNXDYE57AGQKBkjDITOpRiNEMTyMv0B6
HxbyalWaYsKlsvzanqeC0kpWGHLI5FBIE4BsSEc6G4a5yZpqMNuyINplsG1+iQTy
e0ZR4Pm9QvIniyqxE/AOVC930tp9IigRv7yB+8EQBDRzH7Kx4pPymy3/JCJBFKhR
o2h13WcATvv8CE72DmTOW3Nodxwr4nYtxaTG1eaCPJT2bbYJVVda+T9CK2agIyki
+waiws1rPJX8CeWKCO0Qc3jI8QbAcv1RlyVkNSEIokve4FznuCKoVob/AswdUylZ
atg+dH2XDmcsWzxm6CJMA75rwpTjLvE49qHqpmGaoX3TRY+FMeXsj72axUMoYIKa
WNycSHC+Nc1q7MUUBXhBG4EeMXvJkQ42WW9GKya9EnNTWwm0CSQxM7deXhi2lFl8
o4P0ZL6h6VGL0ACO0zXQhM/oyg0fhStYB1KisaRz9NfWZIY8txtEvHaDojY4A1pv
oRfYBhmYokCgcktkO7a094eS1qX8pErrRvLhyZUgg+0IgwdmsxqqEwblgH2oe8UE
+AmsPk9zCIoMjNbZ/2QRu082V+nFyJbxl1kel83cl/CzUURH/bDG8kyrvhpEvsRg
BU2iRmeXQiXIBIRSQILVnPYVR0l7Sp44Bt2ozx2ve44yNkErRgNhgDSpP+px4jwi
9wn77xYxpQdGbSEBxpbkGjhGhS+uZ1wQNeNfQ6mo1OD5izoXf01thd8dY9lFe/Jv
Y2H3jWVGdqRe92mAJTeAk0cZTEJxqDLv4Ose+nu9Xpri9BCTExoZFsZJiDiRDng3
kuChlbL2RXdm3sPGeSerDv0OHdrTlRXqfbWBgvHJvR7ulBSVY6yWk0WhzEvKB05L
Lhlcb9fCynDRiFib7ktqM/hotHPgnBv3PQ4sKQwCy5K0h3BhAlnT7LkQyRRJSqKA
IIGVOXW2OcdYL7MEl6zenFBJxP9MJurgjkXxFjWktpU7I7LxATP3kBQsD8s0UMGK
zZMK4a8VAeKYwZTpmzdjyLmNLkZkWdzijdKXl2RfcS54Piao90VUA0pN3X7RTzeQ
ngKlRNxB3+sLrzmrlOteU07SSAxv9Xhqc76XSaI10sg3fDWzkdqmw/fG+4lEwpiI
+WZvZOAQI/wgvTr3KepMGRwVyYH32KdzTIyLRk6fDT3SxxsRiQC2Q+Hi38C51Kh3
DhczFUEcWqdzOhGVTRRaB/gGFRl350g6w1gy/7er226Kc9fSlUHKp9k5HSil85BV
FD6GWW5okC/yPwCsgKNQpOq49xgB504KcXotXUPq32qPLZ7ucga2POlApaYTleG+
MdO7/xEkSPQRqWZt1xR8tCsSPBQALKGa1UJQnFS+hj+GChQvk4dOg7mvOXQ+kYbC
/9N2CiaQzWRFJAkzC7iww2JT2F7Us0NSa4wL19F0oueVqlUdQdqMFuGgXt/QSjn0
MONb8HplDD5on3SSNwWGrYR4Y7FKf+oWI+L9gYkf9c8lK9Z51KFHC4Dgy76JCeyE
o0FfRKKU3Tag3Q3pIclPSYf430v8CqYT4NtM8JTd1yU7wcadi18oT9aUzEn0pi+2
rHhlhWt2OXCiEj9CPNsaWksl1wTdO8dSeoN+iHUagU3Jo6RofMclZNYBsShlMwY4
8GQrxeHoTld05wOhigju5jec1ij7x43/zJ4VSeGvrjs3zY16z3sjXX9I8j7q08ZJ
v0Y6VkaBIoA+c3Bcqc0vkl6W6nYnkBG4usDj3o4jo6uKB8JZ0vcJTRj/9ywLiUp2
xlY/YywcArTP4nNF171HXUG9E6Xrc9aKg5n59Q/owYuBXGRew19uQjOvVGYCZlpN
rAotQHXNWnnDK0WplEHcQSl7d0O8rM7oOSLaqHvS1XV7a1tMIK7NrK0QpkaSGF9a
mqaVs0bZdkM8SSjQcG1Q7a8m/3fLd9kAXvf/t+BkNZi1FIVeVawbZvf9mEhDCT5p
odrbA4MND86odOyK2BueHGK2vNVn1OoBjx0DmDBVQ+p+zVylDJXddtQTJn0qp2rl
AI5YmJKyGsGi8QOesyx2qbmYWtx3GAmbwHmLoUzcUsbCbykRXTvT596eMEysrrwo
bjUrQOKY5JprbqQ9TzEzPclTf3YlQi54WqVtgjcY6WklumwVT43C/1MHSaSxfEQA
j+jg1f4W2xayQwWtJcXZSQAz+ZXpaWSAGKdMtyJCvg+D+toHNHQBck3biQ+Ocg9A
8BP0i2I4IV4rKwfVV43KV3YgcYpzkGwPnNhZmPRsxYAW/AB80Av9HCgjCMatSiM2
LBohJNhj09MUvqmjuRLHp5QDx9Ogpjj8fOAnAlqeyIiCuCdqZAv3UncbuMEzDPT9
ZyHYZJjV5C50otkak50702bfOLHyqXHfmYFuQhZNvLtZ0bRSzSrw3WNK4FFnbyRn
Z+lzSYDBQVYOfywdr4GLFT1TYiPq8OFoVErqZMfjBi7j8maq2xHYhWj4bV676Whc
PXHS1Ocj1EIMVJ+bBj/FrzDUGxFgvB6QavBhQ9mXkPAY1X7szwqyCeRBqLt3VXdo
JN3BWYSQTtSS9gdogyH5+XB69sLlrzlPLUEzU/yuu3q2QaMIi7vdpcP2I57K6Xg+
t/EAUbPkSbuxdSBLZCxIIucGMy5z1ptQsfsqXdRh8UFk8rKOGFRlF6KJUyNZpVle
gg14njrQyz1gaezkK7qG2O9Vt43IWPy/8YGCNyAbQgNDYbuhvEjgocvWLKQ0xJlD
e8u18bu5m31yIuSpLlNauRofFI/inCeEUmbmDpypOZaIgoObC6vDqTDaOvr3Nw+b
q7Ebtkazz7HBaVYBOyXU9K/lFBclaLCCydKOVIhBect6Os0m2Lad76OdalQP2UAk
IGbD70RmgYsv95XoiOq/UTRIGbMxMQCWyb29uIom23Lf3rBW3525Z1RUzYH9o3Gy
PvzENgihiEWwf7S+rHVUjZmGU9gGkLAUtVE+gi+dqxAc9S5cTdPzYaxyjSByLL1Q
3vVprg8kkXz37w66bfI1jiD9ZlVFSxUJgSjIhVbtDZrF8/1gdLDgtsNHISC5xDlL
zqhd37CFTGpYMx3ih9O+pdMO468iandpW4CY2nQTd88Wfhx34jJ2iftkhNt/O83t
6kClqCIIIpb5hAYhppLwvckV9gHSAmMJCt6A36UbsC1YopITVJrGsbcRl3t+/B+a
rBFpQ5S2GtrkYTmep5MvwJ3Eml27/SweuZ8Z+SoYvgcMHGF32Rd1Z+orGx38TG6q
wwudpRAqUKCtzbBEFGwh1Ud6YyAimSmWFafAMaeBG4kF9PafGbdeWCj19zB+MZHl
O2r+be5oYyi183WdpHQiECLx6hNxzjUYLJ+C0rRNxhqG2l2TNA8GYCivMV4HHUKA
36qAHJTaYx7ZmMR+QQ5HuTbuM8CVJnkRqCikeMAEOXI/68vXE1QFV+cU5afOCyB7
bgq/RVzA2cTrDKLaUjLCjcZDAtmnLNHrA9etWHyE7HLIYO4/Xske0krQH5Nzb6h2
Q7QR0bP5cL5bW581mgG4PHh8AoLXn/3972t3VJx7kysjO85PPXm/vFGL19CQglyB
T4rQ6D2QggqMzoIcYLteNt+zMK4AL8twNimjKD0fvBHit+tn7Ro6qhICSJNqo2tc
aXiPe59FmJQ3DxScm9CS+T/9HDpqb66cuS0EaTGgExwNHLayuyGUnWRLyxtRFdV/
pCcMHEufOE7AaTvpK2i4rUeuP2+b+wEstPNtXyDh5xNmXyG52MLwPamxtHRNE01a
j5zeLVZkNhwWkyc+sKoC90rhJXZVAQ8ForrOyZSMA7GujNDDYb2MLwcbFfP5pKyv
6j7WJXIwD4gZXWKETIaPF3jl0xoJohjPn6cG9UYAcLGwJQwkM8lMo+IhDInrmi2H
hd/B9vdOsM9Kx+Ze8k/NF0tdCw36H4D8H4cPhRomKd6/6fFINnf5nA30EUWfSnZD
v9R+sCNb60o6rNG40DGyc7xJS9pARPGI02/i8A8KX/sgBXFgx/9pUFBNEQoonz3V
X5xvd7fgeLIrRuScLKO5P7Kj1mKFSUybJAtvEcjP2T1CVezmUM3Pc3P5ijnZncEU
NMhpsa5cZz4G/d4wFMl6/+QFZwWrzbtyl5JpYlWzWneMoccjz44W/ksxAKPse7Be
FGz1ZJJvqFLb0OcXwjJsPhhf1gX9pMNBvNzDsnhuh4Y+3F2Cm4PIQ11Iam5ohx4s
lB9sV4RoL2eAY/cswxIF9ID7RBR6U+sP3DnX9q2Sp7yRZ43lV7DSPnahPlyr7A1j
IN3MwvXd1LpLX2dLgIJUe2awwFJMeVe0I3z0O+i18PX4m6Zb3ZcfgisKCjHnWt/u
xllMqdH3ZvuqgstNa5PaFZ7vPm+aVL6wK4Eqtk2zQVgDkcv8VXJ5XLzQ66W2+pml
nsVhYdTby3toGp99gjJczkhbP++28xfhrqpMsBq72GHrJvEYQbd0GtuDAckCN1ru
uuc9Xg54Wn34e9+TF3XmHPmM4A+UXVWwgz8DD9jDbrNSWj4ckjl0yDPCC+09Z4wA
1NVx+gqRxPc1Mdq2A00mEfI5NfdODMVZ1Q639SRsqb+eDpZ49zOrYK5nTWrdrIGi
cDS7jhtGpif6Xfzu2bOgmd8klEXP0UgRojvGtI0+Ll+hPA0NTfw+h5zLSm08cYK9
HmcvbEQK/UDdu2Sb7cA5xtTm5SmNFOIwa4pccGS7WV9kgedE5IjUIO4L3UGATvPU
HkOEOlios16C4HLNOX/ix02ieT0uhzo7BsHyf/E3RE3L2rD/R3PhXihZGJMNmEMa
kj67H6St/QJrPmTopcbUx4rSgkkS02vVMtC+mNnxum+b9zi35yKOPBsiSLbUBa+2
lleges9NWfw8rbwcw0XrsAho+dYU+Web6mCcidFQuWPVM58FbUZetNP0nRP8Qxcv
8AU1kqz77NkSvrTxy4qCh9U0HjY/ArJdsjdgCOcRfVI5LL8igvPe53KNcTNN+GX7
wl7BzM/ZoF4QVMfUygBRw5PFYPt0/PrH4QRIFuWrZfA40GDJv3XRHjSxdKn+dzYX
yDGPGEgBUsMGJakJVS6nhTS82OinHxVYs6JF6pfVMKJUmpdvx+n8WitfHmWcRXR6
PBNmJcBft1Lg7qwH4LOum1cCwLHijzJmSEWdk4QfG6+ecjWNN4YyAH5iKl1aizwe
YH3sCgHirRk27h2wXbMqPlpvJih5fIZP651JDybHMVfMhIzI0V/nxV/FGD3qsSnb
EAlzUcke4J0Nr2ASdEeIqtrPOk3sCdqH9y2ALi5tl2FARlBY7s29EkCCel/eYePp
9l5seVcFq9NL5qxIdRoA/B78Kk7/nM+Z81ec/pfyd7pbl1C9GBqh8YnsdgU5B0yr
dTltJmH27Ocs3g67RdiXbNHqtvlNEhB63WA0cWwhYc1gaB8iJgTWdTBJUJoCU24P
3IT9ChaNHQCjFgUvl1Mk6TfO0J4Vp09aZssUUb4ABFtonXeTOEm1Wh0RakWYK5xw
XrL/iQIYBn2RvnNOGzPGkGcPq8X2QtoUJfadg/D/pZdgpB0nXt2JiBGUWSTOh8lI
6Z16fuGt/bB9LkqBseo+Rj+XEKKXctvQ9XAJOesCA6m3XfvO9zWvwoijzN8SCPN4
aFMPWipDNZYtSW0yAh5HXfUo35zKPDK48vpiUvR36mxjCru7kAtOwE/jvfVR3oH9
lq2FmtB+98CK+qZ+pZS/eeHPkEGbND3Sqo3fbHSbo1jaou3a+780lsg9BKO0J0uG
OnIUyNT997kXaaCtQ4niy+VoZJxKmlY5QGYKFIGW2uO9AcU2wqTT3vw0f2wKaMuf
XZpcR6XyBnu+Y7xSMQVt2nVn/xnkFSFeiThS/FJC9MrVkIYDNjhehG4oREOJjFOs
xm/kpsnvOalVOsT41hoXOfL6qYQSqChpHRgoQO+LjukTe5wJ/G01iXhMxqvcW/0y
qgqbMXeig3Hq+Hvz2cJq2kw0D3BR5AebJHQeCxmMv3qJqbR1D+Iz9li2hPMjNeuT
jNYWE0k/642KL6pNfcpDRsElGI4uV/xiV040OmKRtfJdbyP1bMeD4iLR8xF4IB90
sDaWY/3N/NZ1otn7qEo8R0d1OpBrtXbAxXv0SA1LJhp10yQNkelYBNj4QvHvkyvP
xf89SS1DQpzAJWqqVghlQQhqiV7bEk5cBg+TmJtBgcdzQBHxG5gjmNvq1673Eed4
1y4lObN1BNRmMIzMVG52ZlYwyuNo44JeMeBiIgy/8eoiG/46ZYzGP0ukUIJSpQ6p
BtNEkw8lcRXSY2XCUqBJVTAciVQkkFFkOjaYh0OQbFcsfExY8Fx/gNb2nm65sa9z
Bpn3Ld5P8LC+gl+/an2Othw4iJDu8ijEWfEPFwg2AtXVB4AcbUpQvypWoOgA7cG+
fiLgSlLzKg+OQGIpQb0bbzOHPIPuYcDhX5+YtMBzHi1+o41qE0FIZJIYfpNO7Sgu
xli6NC+mVhAlkz5jRa6u7j+oW6KN2W5VaHoA2EOPinyvGN7H0Fk1zFriGhNXuJzj
pu/HjwncQDka1Q4DaLYf6XHwq6IU4NannNkxWzu7dqiNi3+qqJ2k2apaplchzSzW
UIbJtKESY7wDveMFrGvBuqm0KGwVouRzMzlapZIn8bk1PwhGp6CqqEMU7rKiKNC0
MPVSbT2jU3SUX6k4MTHJTjKZV3RfZZ0o5rJ1uaIhfNQOv6c0+y+w2AsQWUXzB0yL
Vd+gHVIzTYix1W1hvoNyysR/V1dgBEsV/URoW5SbeuQin+r30KhKPaKmHc4LQU5k
UWtuHL5J1Yi/LdzEB0fLGY5rnbTkcW418NwLO7v2n4BnXE6Iunlm4LOGoFfqhFkt
6WcXJorisy5wNjsVNFC94s+Hvit51QznSMNjnPJvMM347Ht1Cv3SPLpnQ72PWESc
Sd6bL+chPHePUvc4T5vV8BB1ScKLhrRoPUjpZlzHMORw5q1Mh+ZfFBPGFvlTZ6jp
cxQa7+7gatt4MZSIfqpIMR7tmMkg4cIu+eVQ3MC8O7VnD+l61wqF/FPzvm3G8Lv8
7P6q9k8d7qtpqK3WV1mZUn1ZYFmxXEArMlCBDUv0nTEeQPW6zWHDtWXR+CxFfUoc
KASL+nGQfWA9/GQdYnPJc8GAxvQ50IBGIfqk1+v+1iawG/6Ynul123tASVjry75w
6qwDB3RKrhps1nW3KxdtF4M/R1Hbo+q26J/hIo8TNz+wSVqI2C323F5S/f2qnvcY
2cU+VaGqjzZlORU/ic+FyJr8Wztbg4XLkvgrDIT7R4j/RasdBcUdYsCC1NmOkQl1
CNtWxv2jq+uxjSP96bim+LbAaYxKxwu7XJZrGPJRxumbkDbQQ0FL2ljbr+E+wJhv
/A+RT1wroabAMN8yruA61w+Z7ahTDSv4VJpJ+xyKySjjqvmYRkDh6mt4GgqbvEw1
XTd+qmUgCalv3AzFu6r6YKTE3VsUDcANgp1Xu8oNQoJWoT1mgOYwBxpeT5NUTI/L
voP8I3AfJH6FWSdyxTCZyRzYyMeSNAYfA/etryiIZOEXkMzRJjHDFGxA3uErjjc6
AfL87l2IswWCrWIhmXme1hYgk8TvV3ATh6j0iBsXkmKLDafzu0aZLUU65yjQjCj6
RQGfjiohBtx52oVlOuRLdvXV+fObx3kHjHU2uGakrjBaUByBdTXMPVJ6MmRV42PJ
13aqX8pf7OcF+NzvfzSLu6r/NUbUgl/nHC3vlKU5yOtXZFHD3q2JE3w1pRSJvKFc
xJ4CXGL54qpD+l9KTbehl4yBvzhhWXmxW6zABHVuVg/0RClFiP6fNxopK0FPZZIL
SW5VG2EiaarZE+HGSYkhXF0ovh1ctL/qclMhP1dugSA+iClUsvBkS8uu9427E3M8
yhbGNvSE4L5b0PBBsjPRhGFKMHJctXrN1aHNBg1T/KdlDwbuGlgSV22qkbZVd9gv
sfiZD8DNChM1Qxx1/OHzVvsIHRbb9/t7Y6UfgATRLaGJUVhq+qJVrYcuKugDx/D9
7TKOOoghyi1VqIjadpNmgRr0cLOgpAHLHRonCPc/Xvg0Bm1zQuHjSJ2jFfjTKyD5
KNEGXmmU1a69FcYAy14mS55vKCxv6RhFPqoCd9Ht6rp1drq6HYn8+aOTipLAuK+t
+3ApS0f0dZN+fpUtNuWQZC3XuBjMs9X9QPZVbFUP7dG0KPtt6qV1A70YRH5bkhjU
jlvs0+n26HYMIEGlonUbLsWlK8r0BQtedPHQkY1MsQz8OW1/mBlDfWb/yVZk2vUy
1KeISc63elfoX0jVmyu7TkGX08RSPNQDA8+HLtBI4bs0zvDs1K0u5T97179IU9AD
QQ/ouRNomGv4qkQ2zAwbRRklos4NU0g6JL7gh7gvah2T0bn80QJZiXrW2geJX/3d
gAVB8YDvjmh7JLTdpEMXtWllsPhrlXeI7Ff8+NcqjuESK2tr4PItuAZfbYLtXaBa
f0WAuGw41UeB8DDhT7VNhKDQxLavBLe4S2w3bSi7B8FaWr4M/vxRtFdRN6lLgggk
i26snO6d9VYOqQk4xq4cH+iRSWVoN0gS0cDYsPZNEwtHLSYlK4s/6mTlg01CGRwO
5IpAtqajNJYUSp+VeyKRJextSW/bUnxUu2sbGqmhrUxgqonBYdvOd6jv1lvytFYg
fcS3QK927PbfZmUi6gY4zQNjXXhvFVTC7AN4DCJk6Ja7fHKI7ZJjNEYhF9RqGCfv
vJH5ksU9/OB3/vYxCJdKLPc5QFVvF3rzlb04c1CziuXmfZExvRlMdg1EwCVr1MND
+5aNNqdnSjZ1/2bdQFS/W4xNx8rK9gVRhhTvr6SWsf7oautDLYb17cZQaMtepHy6
AfYGlY6Cp1T92ALhWkV8CwkGRQBwOomTJWgfAHqVpWHhF4s1cFDoi5q4+cogtlpD
bbu7qyKU2OesTNO946srNA0TfI3dF3ldKD98QLoGvjRlcWa8xvV+T1NzpWShTXHK
CVLjBsxgf5r36UpzO0BYdljK1Xdo36CTm1LsXtrV3fPdRszde/oWdZqU5c+5njlb
LPeV2jW2lN+0vjhW77+M6/iaBSyIGkb8sgsQJjjQYh2CUIwhgBXEoeiB8OL5Qeiu
2NXp93z6TN5ixoJPf076c1Xjyg0OJDWoorM/CaSo0XOgixwXveAE4owBUAkb5IB+
5bHh6BIp2BoxU/n2/5SBKIjpeunvqdFnHCdhp3Z2XlNmxG2az0rNCfXHm6zsyNsa
S6t6iVwJq/TlSzxV/XUCF/TfQsv6a4RkEaTYyA/DINTxnUGA/RUNODgfoCK7AnFE
C/eXRUO8Loexp01iUJy/uaSCylXvZ9Rd60CzQfpSMNNxqfH8umEQA7sKiXnhtbif
Eo4DMqrMt530hYChFrOgq80/dErZSyzqMMHilausZbCiL1Ksznu/8x4FLfvnd1QL
/jz5a217T+ROKMd7X2zl8Mq4pnec7PQfbBDLJDq7W888ycc2vj0rRU7d9DcibfPS
zyI82OCru4K5tM0SCYwptbKc2pFJoJCWrkafv8Vt6qbMthk2F9N/Nvisyfcve6mP
PFD9yD8Yy4MBvv1STdnZH1ih95n0z8ovTDIU1fj8zF8Z4RhMBcWygYHpWzd4i0qV
+CBrvjhhvzzRRKUp16sluKQD2z5gwTwuszaW2jqA1Iub3UZSDPKmFQtvP1qWZ6VA
AT0iyHBP0H8P8h/rtH/g6zRIyaeYlBw7G9j1WcxjfyxX36mHj5ZmmsgghJQAR/Yd
/VXIKXlhtYaqB80kmRNMdJ4yglLNK/q8lbOZh/m1lOvINrc6QM6bFHPqDSrb/iMt
pBiJ4LU4MPairppG/rHRZ8kN2FUPdmGZOI65TtsXXLbS/BGAUBY4P5n1cBLXjQoC
kEiDhLDSyNrggEkqjTQk5JmqsWEMCarjpwT/BkQNCs9v+ICwDuzPA2Xom0e0rwFj
+89OrdpdmGNl/zPhWjJit3vC186BNwXZJ5reP13Ngby1bvhM8Nb10we1Un4ctD2J
NVHueucWqQaOEVzA7u40aGH8Xg8cqw4RPEHO+qubMYerSSLOp0TpMyqlNG7FAtol
7N4WsvNOSBOxqXuSbDSOOem+kDxlJOyYDOEt93NrHApH5Qu/9u+GWuo2jGV6XEYf
zaCDCfGdNWSUbLXdPuODqJashQc3VsxkpZWFZylttYlh0zGP1UfZqQRBnSzYuZ5n
tJXOeHvnPQhERo4Q+oGzezHarbx38/OHLybVXOX3Z66uYKrTuANkjAPh2XgqeiQC
Tt4pJBL9q5KPA2iLqmqgvYFjs6r0/qaxgal1rnWUN2G/gEkBW85NLnYyNj97Mrpv
IxCukT3JSOlnZVrNo9J7IFTCTCENGiM/ijl4uEwCDK1tOzpRQumGeQPGTRZ+BM9/
fUmU5Rs1Gcl4EAnkRRy+4ZLNLt4/2o+ogupp9WKC332bhw98+LOPGqELCm+La5vo
xT/P+hGNCHywVqlL7Ni20vj+6NeKwIQqUt3fWhGi/hSMEkd1gTOvDwzYwgL8cOnS
XlAIRgv+BGwyNScQF1M7v0fkAJ7yQJqDVPyAz++zqq/WNeC/Ey0WB78femm7onB7
riZtQ+cYhH6vrYVCg160mZ7OxC0dYqMGFPI9Yn2VUIa3uFdtHZfum+n6wQxyx6fE
YCxv1LXqvaEefwlosEiWylsrlHNGziiq1kOGNIOonwCKkx+/yHU8w29MrGJFOHHi
Atw0NNgxAsU81YAPjz5x46Kkb6XayF6RTAJNecSUV1DmajNcJSaGkOQiSu5C19n2
srdb2WyujRNJsS51YRitsnowcrMEBiIjkLZzBENAgC6vO7ppKyy1LRqtb3jSBLjK
2zw9JSqiYPfthCM3xNHikxE6umha45LQ7O3iTGGLHwvofpOiyjMF+y5zRQFCquKh
tn7gtuVr1cdQ+OUlm/EJapxI799FCWUR/BHD5E1rFkYR4uW0NKCVIcP3ujLVe8bJ
S742WpD1xd5DX+LFusrZ0gm2k4R0jwN4PkYnfHF6zqE/H6+d3NbUNqBh/fCLhuQW
C7GtTrMxTRMzHh9DGX0cBNB0AgqJ+CiKjx6pptRdxN1YtZ29KgfhKGcIceMvB916
pY9BecUwnwkQl+moxSYHcdfA3nKDyZjy/K81pSt6h/lqlJWzkWXxLosCmrT2Io5V
RImrbsucwTvmsduCPFMiRS4KxzMwy/4FYk0sUH1rls/1sE52d/PrNa/ocgwjFSf4
LYuRZDpsGTKS0cM0IWB7OjagVi06a8mSvcmKlbYGJAkEsNuigjdfDPB6oRc9nt9N
1j1q4PqEgfSkxVUfKD8Z/0OR473cIKuojUzrUhQ9S5AcyEI/uaVi6g0sjrE2gZk8
Xrabh0u0JD3wjNdsJGkQMSzE6AaDwvI6N2ZRHrD3bSdXGz42PQZYbqjN35ZQAXVK
VoM031gxFDz6N1kJ0lc8Neduuf1bOncrS0DYvnIW/bzQy2kJEUaEwfY/C/5egZzH
qABMCc5MytwvfskPPXmWnSIHxjmdpBoyz4J3tKwBoDc9cs7nsLtPZvpsIERbBxeZ
tHwbtri9ANuFi6UbA56j6wYHON/on3kguOA6nwqHygzvETIhhZj93GvVJmUOdiJd
KW2f63hKIfdKGsJYxHnY23TiPP936ioTmdXvE44yk5yr9hNQTZMpnQd6737jNFGp
9WNACoKuIru02WA35tkNmxU3si5KpcuVJ92pmQN12x0s0EhZ/0X4SLGY08QWztVC
YUaK+51qs95FZ5LXrITY5T91G+5itJcDZceok8wbt7HFOLMEpsTZiviREMT91tSP
3lQ8ZsVmdx6lSM+DLiOsidmfkVpX1cu8Bj5bthsxSMU3kcEKmZAQldZTNAZJCh1b
jq8IL8fYF9flTveknQ/9ckEqRMH3crjQM6kYSOIlizQE/yDm7Q2rOBUJbyyBwXZT
ZQ+6L74oLm5IcVdMDa3mXLK7++rAt0Pblh0DHfT/RWNLxDmF/egenc8U7tnK2Kpi
XJwGf5EZq/wwARYEocIFGcDlQ+Dc0E3e1V6pPlqLJj1Yb1FOrG9ZNoGmJS93ejjS
PrSQDLKEte70pqdCxV8Td3e23YhtSoAO39FwWelvFcp99f3zc2z4mBkLk8XcgbGQ
MRmcb9dalzdupVGUWZbbyHQZmtLKTQvJ9WSzU1ONyLvBoR+yBLKagBbIVloprKU/
oPK58wENYCOqQX2FmL3SzcqJ5zslEAqjWM9qRWbEip3X5WDt1WF/d826kXsS4x/r
IM02Uafk2ApPeRz2y9Mgg4sumprW8oAJZ5WjPlYb2v4ly/WZkoDfATc39AoKgN/H
ujRPVdQX7F0epzWuStcajnkTagsL8RJ6nUpGut1Xc3E1owjPR9yVwyHEVvbfnd3y
FrC7A2mp62M6FQE9B0Y3o1hBMA7n8w/DUxQ825XssYdqTKHNT8ma/g7PI4abFcFw
fgAsJRREnu6yR0qquqTulTfwSY9SmmSE84bPbbhw3nUOKXgIIHgStPMFib7gdx14
zxNTDaZDMZIWRKbeKzb0ITSYyDvDae/BsgS3LOo9QJbM1CQ2PQk48KNcH63wIT4S
qmgXzU1GMHKuTfT25rvJ210AyFOxXpfAe3i03qxcUp86MdclsXYPNjw467sQEdh0
Zx2QClu7vleMOF0LeyE+zcHzkqTZa31erKdmxqwDaMtYkn121JMqVXax/4G54mr2
2167B/kVjICfGuULZaXw7rrcCYkwfCbt6x3oZt8ybv4/1fY3v13CQ5nP30utouVu
mBBaVrRJqOo2zjLo113ggJH1Z22mlYjNTcLT5RfeBrRyNi7BGBG/+KPUly5B8dJk
sAYy5PDqkRHymMw5Q8izc8mBnSBIliN+1AQLVg/EVUPhFClgug9PbS4uI572OnPb
nEgL++BKXlxyaPOLGjq5mJOjXqvZkshWCovKrI7YhpWmDCiNKWxVWMVnnKaLTqKh
Q3osM7dfx4MMLrzliHKZx5lypj+8MJoPdGy4/+MBl1jVkTOKvj1qnxFZzOOfkf29
z+xug5HFgUYJBZnhUnBM5rRV8SULXOVXPz3b8Vm3wR9VrYVkR6zPkdqFU6eeSq0X
Tzfp1b+iy1bFHNdHxIyPS9qsHQ+7e/VWanlHmaDW1EspGcaRCIHWEDSAFXG2qZeT
g71ugcatDRyM+eZ2SzJbe7nuTE7Ic7+jLAN+/FGaRyWuX+3STVbv/AehRDSQ5koL
3c7hPB9hgu+d3jqC1IFPg77J5e0HjgxqJSJM7L+ZtdG11uBXRfukhCtFRKU7qtcq
aA1DsmXkSioXzNzWyj4U83eL2mJ2rQBU3dwregxK4X2jCzdGZzsntrM+bZV6oXJP
5pL7h2ZCWy83qDWG1OcuesScPK80hbM+I3QVQWbOSnhvIDbDH55b+6D/31ORurkf
qCysDRhecopgukRfHWQqAVodJdRs7B9cxFSxe0m8smmqwhrG3pIq/1Q1XDx0vkPz
1TGxcpz1QeshojQ5MHmaHu23SSbBAdRUEY1Sgi8i9lw0r/lOCKcJcFBUXbAIQLe1
ZVvoRapHpYqIts4fUFWQ04XiQhJkcLkZJRnBBSEmdkG+uwt2MmMnzS5nXWu7+fQd
6NsuMYLAZ7Oe79xCqkTaA1IYKG93Cq9+3703t9Lg8f2v0vj0G4znM+0eCy9SCDKD
7i148jL5/wOgytB7CVNeff65blJ8P5uovyWad5i8pNdoNuYTZqXtPXxd7COWWPr9
9ILqh8wd9PCuiHx6UC38DJu3gyJPcp1snS+MmqQQMQvbDlNwWUDSkEASUhQspBO+
IjkymGrndpld7++t8iZIO4+CGJYPCqrgC2f9JGKEqWJ7tYCbxh3qNXQL1DgWb8Ys
yts1S6yT6DwX/yeWR9ZjVwHxRCViewwOn92zbc4U7gtSVHpHFohrto6eZTEM6Gr6
9437rz7WHZyuNWnTEgEG0VPSR8ltkeeAdL2MGoyKrhhM9SAka+cpCIyZNwJ71cRl
rfvJdrtawO0TpsIIXOD578Rlm4zcUBPyFkoA49iuPfUgXqhew7NfLPqzDndn6W5K
uKXoTKLFDuGJhf3P5oHrjGpQFaY4/L0Mgdq1MUasi6UnA+VY23ZJyfONgnMnKixS
fwM0FTJOn5vEh/4iUPY2lFziRi/6wxBlZHPwBMeNYe3QZZ3X8wTHn5RJ8/ic9fME
Jin7ofKFCx7ohXXr3FPVwoLqGJiGqim3YeqcsS7KmQYOk9DSqUNW6A8JDa5AFKGu
4NS9ZdBPEoFqLR7UwINXnzCKQBVXsYLp1fGP66N1q31J0edAyAqf43+7PC9tjvAQ
AOoQfAY+TUGQ97akUGMefeFcjvwbkCOiOCXWrnV8m5QH59Gwhpu6V8Aau1Z1MbaL
SEr+jZjGpqQtANDbSUjExKfmg01NJcf46twraGx3No/slB5KQzLhmbUT3WE9KBr0
AS1v2EyQFdMWV3MCtkIhzA7mrchg8DTfhSWRKQssnamYl1nPZElpv98VGvdXIucA
2XQGkuMNntCKYaOR6gqHwBW1NayJUfvjutd6AotaMYb4DwraBGycaOxtzemmKQB2
3Rxaqe+BF9iG0NoGPYAUSYFpX8zyZ9mOfKfw3QMvUiV77nF9NnNaKR6yvFB9AlV/
ki8nzr75+aqD0P5YwAkPJ9aL27Mx4nIy8ejKTlTgxFuL7x5aUiem8DR1slvkCrU4
FClQ8Vsygw2eUMA2r8HPBdfQB9+BLMpyHyBMKsivYhRNpcTElMX2tPZrlb98K3Co
6t5NvkwZh01B5C118BT09P55tU69KPuAlUvdh5gZiylnXXGNWU7NTYiOnbWyuF3Q
6kCxc+kGhCagRuOIL0ZV+M0gRK4dwlmf4n9ZWLgAoqayfKOSN5nE2cqZjZEEdOPQ
5bm+o0hcXItqUpwQZJXJnNHyJ8CkKoDsQGTtq1qEg0eH/Amd9NzZgXvy9XJJ6Zg+
PPRIY5xEO/orXmAbOoWZ5Kr7qkK7Ce/uQpgAkxQIei/1fOwfTVbwKHkMZZdlNQWt
Z4PA3DTLX0/pMCukg5jkuIq449I9E2SER/i5gTqrFiMTnzoplkL8PKH6v64aLkR4
PPQpNO46mJM78i4aY8nrAg/GJkXzPYcZncwYJkh9kVvUEcGC+q+kG0vLij1Id8hJ
jf1aFcB5THx1csHHu0THO7IDPvbQd9dX6Z7Rtua86RcpcJvwcpAvRi+d0QkyUHQ7
dtbZUwnu5D8563W92BBGkTPFMI9HG28hX7s21ntAZcbPI7nT/2l38Qu82jESlhgv
V4EkAZWlNLxFo52lxdZep2HCjtVWPp9YjMWc9CKLly31X3x+aFJqeRqYYgSI+JV1
oNJ/rfFS34246Ljvd/pfPQO5Gt7vqFBgQ4P7ubi6CI0oWjJWjgbolP/4o/9fe9UP
cH4e9kHhABr70fzb2/4rOni6fmqVmtyvM0/NRXoD0pmq5zDozWJbUqWPCrRNguXd
6Ryh51XSk5Mzg+JjCyk/WF4dtrJzPzT102Nl8TnHT9HqlDsC8NGuDojEBtXD1rPr
KSRZZFIZGpZmR1It0dLPOkMbA3v35OSS7DRNzChPIG1SPIXwtLgY1i2q+iFYK0g2
/fj6wSoEBp4NYxVsp3Hmf4v6EM7asFlHXYGFAySJeiUEUO9QJD/lrkUXW4433bsx
9CJT6rBQxmMwP8+2/DpcIeFEBFnn4Oozmc3oue7eHaUIoCU82hqfZTzeXRSNhWrB
V+FKi9BPquBHynOE8Z7EcioHtellfY09aqJEh6ULUyk/Z7FDNUvUbr+oXPEgeK0D
z2zt1MzYTExbApoLjbl4aQl4dgwtMPpadHhkEsH+1a4jX9PGdh1lq4FszLSklW9p
9NUGi8aO6Y9fboCL6IsWMMdPN+B+FgPctC4up8mscbr03PDlVS4RhsDyGJdyTpIu
5jt7g416GioMf3Ph7LStLWehTf1MmQg4adO9VwL/Mb1xQ5656PuyrRsV7Mycfm6A
XD/5hCAfCkHpSCRRv+WmxqjcAeIMGpwnLcN3ySKoyWSBUTxGFBT1OSKSwqgHmzHy
Agji5iPislp+TugD1erAbziayAJ15hb/32yAsqaDMV9hpyVWyVEskFmCgHXYjDsS
FGrsSnZL6UrvjCdxjOoKnw2GGAhbFAKeOAttggbNbDdiRoonxO5BD81juwE/j1Tg
dpIlVFvztPn+HB4DJVcfXHip/6SUHHZbrm2sMF1WttmrqbKkRrT9d78x2r8OLYdj
lq6Yo2Pd8rc9nSpcOEss5s37EdU+dIZX35mNcMGWANQjx1OhExWeRQPMsjVcW7c9
0yuPatY5vgQKQ/TU9VD8Z+H1e4mNxEFtQEiCd8RJpy33NJa0Ox2zv8a6TsMR1vJ6
VB63jYFJzyrOxSePMVtC2OkVn93penUoQW4C95d2qdLgBWDNNskdmn3GjxSrfnCe
oaFkTIfKUs+cZMtPoSxRL59wXssvlnQI8SNbcoHs0t3ifrkFO7jFoM/4RAucdAYi
GPEWZrbPR2jpI+FQ+a0n/5cC8oiXXi3VROTU+IVfbuNUFlcmlLnNKtphtkRhtUFx
5rTAQh23HhSb4cUoMAQSeup3mW1WQzwrvi9h47JCcRLekFwHO5OTVQeU2yhkgp4A
Lh3MkTrArilso6fkHPfJf/JU9CIyUFY94oJ9mikAu7KX2vEbWlqLoMWCpIgGYKpN
0TJPk4vAuhZeHnmXKs/byf6AYU1CGvZoRcKoFseSMyXK3ePNSroRlxHv6MGs9D6i
YkQHJ3Fy08tn7HmfzxpYFlaoUbX1V1EL5LT2QfccCjn8xmSIJD4+WlZcsbDhPH0l
Wq6WCjYezQU2fep0x4P8+oQvIr1o18L7zET6VioX4LnK1iwbMVH1sksBFSj708xF
hdk+jdFgsGYkk5gBgaEcMiwqGa0G6PZtLqzhfGiB4AFWvTS7kNA+VENUdNeukoUe
A3J6QPYBaJwWkp55Ah9ChBxDqpa3VvPaEyCmcEaCWeRs7EoJyYuxFwWsPlkCW2dS
fbziDl79ghxb99Lkv2jEv3q9XKv+eE+kuRAUfoa6ohb+a+MItimDfFNgE4QUG4jE
quDSyJ9HlMSplUXK1oTM9CwgxrT7fXIvPzbDdG1sCud1qyfX8biDW50dBkbcv89A
gWZ3lVT6z7HkEs44sLttR3pqoTe8vqpm1PZALf1EtauyZ6xMsIOu02bQWx4O3n6+
xEfaZDji7RHTYeshRDDs/oYW3h+9MXQwyFU4GllCyXhIyYRkptwV7UqECvXKBL5m
8v3CV6UPG+1oJdktytlp+RWotVchNa1Oes8MOX8dJ+KysJ9tIY6dLlk8B/GqqlNs
FYhQjClEY6aKwsNTOswtCGzZkj9YGJUrq482+gobIB8s/4y1qka5yfPdtrHJalHy
ZKkTWYijQPJ4WWcg8YZ7Jj9gUOICgMGKX5ro5pbQOxsHPTb4y7KC56//y/ZDhxi8
hw+Z8G6UWlvsgnUJ23kvNHLoY/sI4UBZdyy0pfdH8GjHnXsl6TnnibeFZ4XdLWNh
T7O1LzYqn48XYaJqVoK/tL7wwWdvt35g1fmjrXu7FkhqALfmv2cwyD8eOqG1aMS9
9BqdMS0cJZpM6H1xGDIB/jDmVckqokszY1fXHmjb8R5/8Xxd821RMP0oef8H1NpP
ObSd2QDiTB39ZDTKW0X40COzwrxcAt3IuGKTqGGFEG/UHvkCfp1CVLHpRoqXfbTk
PjGyxULoGmdn87i4HCiUQ7dH7AN8symlDPCDSJGPxqAVk8TBxpf5QPQz2N5f4+Le
viXFmd+FJ0gSbo4UDjF7mU/HmgvxA5Ikn+t95Ps5OJ9o7gAqxtcm7FgmO6dl9uZf
F1Vjqax8gc/VHDIRDBRjDTigGiHmNPkwpygVsHYN26kkR4XxA4pWgiscFG93Veqg
TySNLn0SmXQBPWBrNm7ZC7a691+5ILLEQQ0rwuYvpM+B6byjBlPBedQWT3zwaFPB
BJBO60nD78h2NoHd/pKkQobH8lnDBua7My9K/s+YxtA+98l3CYNNQeCnR62qvuav
ki/U22J5UnxvoHOi6/pw0E9lBmtmDFyTox/gQ42rjUf0FC5ufYFqIUB3RH/OXs+Z
Mcnkb7wy9XKkY6GCbk0z41eC3pYWkF5K2g52H13gF/OhSvFeYmIUf3nC1N4++PKP
87L6cPPQCuNcp4eqP85Q7yrXzHVrwbvdL9CMPrC3/bGbZPEG88QXXbhGcWnWlM21
sky+EF96B1C1xpwskMDs1KvOilyA6HU+eLPAo74RWTvo5VG21qbR/cp4YrMbrRaW
pKSNSqspg1W34pZ1EAX16bwex4/eV+hQoJ9AuN7e1WGupX1twrefWyuWqRkINbe5
v2eJCzkw6Dyc3CjQLJKGUulVXkrxRcwL6w7aXaVZbfvU8PN89/c0Fzgkl/hKpSBB
5pUw9GwHBqNOlRPFZSyhipoImxJHkvhvuO4dxddjjKwa6lUgFAG2iCUx0TskeThz
GjgSJfa1zJmLqaUPj1Ap6e/3RsmaTw6uz6KxUsF0t8iNNW0jmc7StTiA7TgpxfU+
zeWn5knyzgMUH+hG0aDYlxC8cmsl439BRak2iNqILsiB+JWqkTqxYnLIPFOcMdu6
LCyxF/S7TaSpIVjrzygcfRnIHezgnkum5+/pKgJKS5EnyS7JU2VjWLMi1Q5B2EOi
tW0lESooxW0dGYcxE/o7SvaGwNxA2ake9LfEl5+xGSqpGQyWuuArmQHVQkhtGVe4
qrkMs8L2WYC/vlBcqFGCLQj556LQGZti0XojMa4OZASqnXVYMXr2PMNvqfL6unT1
DDBZmYu47hWfuxPe3wTqxc6R6pP2bIlK4trnzem5cB3DH5f63dxuumyupwPGoDOj
8/UD8OW3tmb6OvmAQIxDKECXhJNstP8PYh2sZYHTmskbMxsmOcXpOTrLI8BFLL5f
J0HcnfRV8DHlNqc1QXqbExNc4pC3qmcff7JnxYJDUeL6Y3FxL+UgVRXEoBeBkTvR
V2NvXymE5wjar8TRvb3lWcpUQDMsOODJwVvYV+Z5RQ2TqB+gJaycPijc05ilLdGv
EbJf2ZIxFzJ9Ah25Zxv4GcCIqySmDwambXPTYBkzGQ5hHbCpB4XPiyhVBD+Q54MW
FdDGfwTawcp0VKAhQPxOwWcwPjOylhomUHJlE9b3DHVOuFknITJTjn6KjloDpMog
cdd5LN98NoX7+FsZ97yufP2LoKYRW0tGlhmpW/Awvu5rPwfdk5PAEgPDSqvbzTsT
U5nvMe1aiR2vkbxwi3QxYQ97GwQUjk0kWK9Ff9cOBX7NFRl7Tw6Ivd+orhRXm0bH
xdXPP+Y9wrZkopPzwofojdAE2ECXBeS8Yl5EpLm0kMi+pC0pR8xJvqS0J+D4t/jp
K0DtFjfpiePaFHsrmZeO2Sf5u0+q/INaxOwMbB507twf9ZFk1at3eWyiM8pmSRSv
X+Awbx/EmiO8UNQ0moZSh99Tc1rDEa6370rGMPZHmM4gRp3k04ooV/VsqX8kjU3f
BI+G6l4+2902f0kNA1b3BZRItuCgrUU4syRMTEclzrQ547Unv53q5h+Awxel5MK1
Vt1V3Snsqi9LKRT6MICE66G7ehmlbt8shLN9iKlyTHKJ6hxVc//POqpiAe4MdAg+
z4EkV9nQozT7M/niPPbvWbEKz1ib8hMttosSG4U5h4hZSg2/oNITsyCRoq6z2Snl
Tn7n8P2bCBlAIkxQ5SWi625WK7VpZzBgH15CsTuEiT8S/GhYwddISktEAYHMctMO
9pVUPlgH48DZy4yh21lGE04fp0SkPzLlRwLdmq6UFxojk38EsAeqCIyqWOQ/Ih5u
Wc4X6gs9bW5Yhu7Xg1g5QGwGlj9+e7cGyWUCjAZ1lphxbOs6QGwerbD1VZA9bH38
M4uSWDntntoeh/Vvz2gAlPBIWT3VEFxWK9bBxtvH5yKx3FXS8ddZFhMLcrjHFhBi
Y6bYfDxwLnEJaP0qn336Epvq+YAy8x6T57/bfFKrWo6WfPUdZ5pphf7PvroVrDP8
nl3PWEOUZgGv0vNvH2IvmzWa4fc8TYsH6xKSbjcQwzJ46LCfPjYTuFxCXMxDM+nc
bkAEi3AIFWBWTzRFeGcPXmKneOpCkz+A6MnoV2vA1t8rCGf3RVbD/ZDwKK8lDT43
sANrglU4T9Eo1j2Ur2ekVKoch+Ul7iiyQhQd05BtGeQgfsdcpYiGxd2Lda49wFP/
oE3wKn+z8Rd09lzxQIRYDiLnhEt8joGkVvhTBsGd5Xq5C+QRYgjSiZTKSzCKvGg/
+JnhcJAfDh2Zq8PdQO7q+ckH+gRhg32Z5/LuAEJfGbXFONKsunoKYswAG602Ifsi
l4DziUgbwK97SEh9G5Fans2047L7r4wAxsPgX99ONUhVnbYWAzp2yQJScTliDlxm
vOuOkf6JgWoXC2PiRR8ix+35E9T+J/2f2PkRzzVHa03KVIMn6CIKYlDX5AdOWupw
QpwHVJZnmC5SbFs4GTTx9vqXzYQ3cFnKD7zT6gd8d9NhwmiBHGMmwaMLQimth5Mi
/STGWbWw00crrdUlh/rTZh+2QH6rDHklhRJJZJ23qTdTbMlFTBnAHtw35bCTWZyo
mGyfFvROXGtI91wr4puFyu6cM7ZpM8Upl4F/lY9KU/ILyLovJaqCkNDwwCjR2uAl
diJIwKuP3xnRTdqren2dIfgbfc+UUX1diES060wm+VaG59hdfsS3BD8MtROkYZIu
4Xgv9gd2cwa26DMBrTG0YrEDKCf8xBzTAHoo0wCuu8dCLKu4D1lBW6+5eyRKzMPF
KmcRWuBOUnY5tdyEAtHfXbO9uBOojXmNI63wN/dJITrIUoKjjrQ2h77Dlt3irxb5
zEwjgsB9Ais2ovtnMJ4t7SWFr67EViAryROiSZVV5LjdTgMcUi1EroScxkhGR0un
7pb1/ppskeYDsR5tZs3er8v9iryejdDil1YHimn9mCdsyrjZkCvjqLbdfEVED+Se
89pCG/KLHR2eg4Q50fW0EKq/uEGE93xPkvNOwHUwVeLulASzSJgvuJW2N+lklX4F
7T2v4/1M6jo18QO5RuBxxxpgcvGwhWpUndiuRwkHyJxwOw81Kn6cw5+sAB3Zl918
zNNNbru57K+JyOgljNMlwHmy+KcwmokX40a36s9YJ65o8sioFhqWwpQqNXlm0OO5
CSgTnkk8LNqEj51gvRZ3v9xfalqLDeMrW80bMXEN2g0eLJHg5JsDPxjDlSOnvv7K
SMDmcuBXF2fn3PWntwbsWzN1pWGHtigO2+yD/Aze/l5x7KUj0ipKZCPHp7Uutt/o
7pqHy37nvWngOVoBHoza3brvpkffSVE9XneTFWFdvCuluqoHGQVmN7GCbeyqzA7o
4K5T3sMPSpgGquHgZXIG5oGyJcX4AFY1hToiPwwAu+mCBAsVmY+HAr0XlN35ZS33
f7BIHDCwZM6Xo0Nz8B7KqaIsXNaJxYjnLAjGUZSB5HrSh/+cWAH4kDQwSJkP4hSO
208T5Rxl9i11PJqnabPIQEjK1wwI2iAwblqsR9fKcmPG8CckRUSRRV0gB6P48HR/
ihTgiYlI58q8CgOA+gqt/PTsh/PtmlY7Y4rSxvy4j3LoM16rYcKqHZD+ywrj+fzo
UEqpkCOsKUYpTmwfDxi4ifh8DFwpVnaSZxa4aKvRbDwk5y1jEUHrlLWh692IDwev
obd2dftk3jX5DKKCTqeNN2x/5DTDxytPWCZ1mRS8W/hLykJsMD/vdDAcQMqI5GCb
F6pcs9r23Al6iX1tQVCz8VLp497qNAgYNiYfIYXZ/D4isdzkHunOWl61bYc6pM9D
oQsDlhD+XxG4c5dUN80GtHFxXH5mgSgjhx6w8TLk6M+ItzrXm7Zdgb0NzvBSVDlD
Uj7FVLCNvjfZDvPRP1nGLD9RI1X8/A9ZAfbuKSNkGXlNKmGZA1+Z7Zvs5QBMS5wA
NBPEBuxkBY/ZD3f9a9p/rZ8mDcEINvrj/ucqUemERGmNDu74JVcyc+mgHMKtoUh/
EqC7loh1QblloJ/aGzgsTw619HNqLyaIrHU7GnN5KH1k45YBuo4e9G1ssS079IqD
fMCGNnJdW+t4SsrLtY8ue90lTGeEbln4Kk+dovnf26VaUu++AXE/M5l5/hQ2ql9T
7oE5S1aiTXYC/IkJzaV0KwzZFhQ9Nv6C19lLCM+8iR31nlxzyKaaQ7nfqYsRAGc6
DCrn/i84yllaWUcYZ72iselbaTFVd1CMwFH3a0Weg9iYxKqQmS6KzU5wJbbuMrYr
uMQHiTNLa45U+MON9HO77wm79Htt1J+JtAK4SWZzPinpz9o72c+5wkP53Otrqox0
F+bq5xX4V98p4tkqiJGU5zNJkaXPhK1xpMvZbdLp106nxgANlHmeoLZJt8CNfBmU
WFUYNXP5q7nz5bPmR0hgXVf2889RojHYRFf+JrrhOqj7r7eue+s0IPQGC9b5Tatm
NmkRrh7/9kTEs/DoqGMM9bhx8zs4FOm1Z0gCgaYj8kbzgYXmaqLI69f+jswDKK4J
sSu0B/htjERV5XlOYxxVBXZe0s/03JPqDUSKlScWiYfuEhbP3y1YzXjMCbmSiXw1
xOy6OKHHVC3HDAL9FENnOt/YWJSbvGS134j2YNfu/hH0Q4d9zvwMhRLPBZrk9Q74
K9he0wx5Rf1XXIK/n5X0AqU1plOrMy6KDHXWbyRFcwPdSAgk3T6YLVhp7/Iia1Ps
mEZf4l5caYYFjtQMnZuwVuqhjt4wMZerzBB62X/0dM/vFDcxhvsewKeoraDP8Tnv
8WnSYnjYdLiWYBTwIWzUIg6R7PXlj1aga9mjgnbUCcJDOQFv3HZuPco8y6KfuUge
690ANOEz54HCH+rixTtrtHO7obdrpZPMQyjFVox8caLfJvfinVkPdodwDN5WdgtR
i5PhFDYUywgyfED+Mxexnbdq2TUgPPAbgE8WxXiwJFVh7KruJ5VA7lcXa8Ohq0Hg
DItrewZ7cqi2Vk7M4xWEIrgZHP+7kOvhq41D/kGWkrXLEAzW0PXAZjqkNcrDBAxq
ijJvypYnENsw/VFyQ2UdCShYFRHDWZfoH2mDdWVlDt1c5pCnDQpjbT32lqTUuAAQ
5iEf9QcJREenjSKsUd9YupI3uEuxGnN6DdBVDWtaSuoE5OtthetzF3e/EE90EnSj
ylP0CyGifjupOdAN+fqkFMQapqG8ix+c12aXNkyZOO0lW1kaXieK9fr/2bFZ5Ppk
hRgInrEao5fIrOjsVAZihOuFbt8ObdZCqiXP2PCUcEA8rxl1Z78HKd2Jl2VGqjTH
XYob2qsQU3mMRAObcyFRkqj0hP6YkfZ8s+swf59eKTZN0Rpk6JY0fKn8Nx9ae/PI
MLYUBWhL8nSTHo1eq/qnVu1Wv34V8D4uIQHIcoeT7MeUv5PDqWeOhnC3GmmT+ZXo
AoVF+ENBmrD1yjnFufZ29a7RSYy8T6YWa1Ke3b1byEqEvDDEOMZRFc+4GYWJmyc8
bcJKW+nUQT+jzaRgipvruWsiUqIPN6RJs8IkhfFMf444RieTAeLoXKn28Ak992/m
sMrzb2o9nH/ex23ER/xpUyjjLGtz6xcxSIlJavnyr5Gw1kvKKA4Cni0Y5dNlRXfN
UWAidT7usK4ZClZydE6XQkcQoXcy0ibSDTvBRo6oWmJz/0coNY491JS1Xa+5dvrs
anPbR3LM5ZJJxm9IDngPNJQX7e0legzhnuByW2MLZPW3CqGYVnLWKTr3bMnx+MJY
4rfiiTV1IdKpqG3UFtXlMcNuVXOfYnE0hyV6r0Ao9PvCFqZ6J8jyfkSg4ddOXKia
m2+6qdSWpxet8rBv43h8c2DyHZFPDKL/FA9EdA+VV+vnNwgIYPsxsImSB1Le5ihp
JpsgNEh3rziggVaui6cfVm+APV89OxRXq5/KoA5QrKIOudSJJaw1Bm/0GUdiEGw1
ci4Qx0kuYvV6E2+5mmRttqaFnW1JFfXiIocHormktZoYpsZCRDK9L4TEXNBTvRRy
N931f9DozwkR5FzW1hSaX7KRnsePMwVbFC8v11wyojUQIb/72OVoDk5Rk8pwQT8a
LmQNJmiYlfn9gJPI4FzneMyyO1j6moF7xRwFGYB5wru01e4L6Utp3PoU08/eQLTI
d4MV+wO2v7tNvEB6ONogM5cBTIuIYpbivOppXNU2FT5RpZAbus/vpEWr2v1OrUfs
L3OjouzHKqySV7L5bpjNNsRhkujaISmEh8ApAqe+qpH8lDt8T4kj57EFJMnAd+QL
rNJlwwBgxz3ncf5ZINbUCjU1S/Msa3RHySNIlBi98zQXjl6abvT8YMp0TC3uFSeS
24Bh24JN2SVR4wvW3Sox6N+NLetf5ENA5OU8dsWLe3cZCRBrCLgoexgNOLfS1m6p
4uolttMFx89fcS9cjgYcFV1Su8cIJ3d0NO+KAta6RHFv09+x4ngUmVjBhu8B2mdm
95yLNENzVwqC0x/7uraZAXGpYhAZznNTZAPt/pCPrRPtenOqTcigitb+sjNZdV3t
Ai+o83o42CyVA8t8bbkS0SxQv3cXkvZ8Mwmzy3Ztbz10Ze9TNAJ1JMFHpWPEEC5z
PsT1k8tOWL3/o7FpB5FEljHQJoR2uKu+F1hkK9R50IQ9riB1HJqaMwJz+/frhX85
BnpOkJ5AFFqQrOoNKgXd4Y+y/Iu7eU3ArqICb6NrBlIcX5E4OniTnJ0jNgecs/kx
bCdvIwWCTvqQqaWt4tVdQ1i0SwDy1DYD1c0qq8U+RhBv7DcIC0PT//sBmbYjCnRZ
MWzYvortw8gxc6rGoS+TQ9pD5x9pMqSMrsBVY9BIJowL+tU3EGFOvAPuW48+OI7V
JNrIK1RhW1WG3a0/uz2tpovvc7r0iRaHRx1cAxUuxDmO0Yg7ZZO0LeU1ExNKoGlB
ZUqFTKSJwwg3naxUmwaszXKzkiYb/oJNSzBhGvs7zO7OOti30PfSN0K2+epN1tlF
GD9imuPSalqqD8g5dEu24b/5FWe7wHm3rh5RNZY1dZMNYUY4wEXQ0cllLE4ZhnVB
4XxrbaCbdwR2JAuJ7vPMVxEbpToSxK152CS7Jh7CzR8ILFy9PPEbKr1y7XopAzPA
E8mrb/ndmfqgkbZivBDp3Gba5LwRnqwo+8f37Y60cltvjV+dqDVkz7UbPlBXqdsl
DOeSKTGS0y653PWtrA6/DF3vAWZ3jDlk2Vypzie8EljXwevPPqK6/ap4Yt0O/n6f
LNf9BfmjogfvtjXF7dN2xb5ya/DBbZGgqqQXo0DaVHZjevKyYe+TndB9PZ4sZLSv
j99JZfEgis6pJCumonn8Py2rI3Gq1pBL6eUYyUH5uh/bkc+kv44ZCwx6K0OtvePF
zvTC8uoWbGIrux22tzGej03ninKHHV6dUVIZkWDuGFFN2a/ZKZOh++QMfxk7iAN+
xC0P4/BS46c1sRrNJr8LWZbJXremUchXSm23NBgwCyTVSxxB3ICcErimwKnMga41
zkirl+FvCMV/QvdRb9simb/IWgFk68G/kDKSGjQUHw71byCpUm3cUuuUIGDuzydF
G8culCsjahf6huZHagsDypFWyf/8S7wj9htDlfDt/lfOixaNMbHVWTDYit45ggsy
SMxfjT9gBmAlwjGgRhyfwzW4s8iOrLneTy08+cRcGY29dvdhkbPUI41Qqp9GEjGV
sW4wWGPXuzgHxMV0BZl3YXrLspBBh4QnIuBRjMd8hqoMt/OaTzbtWydJPaTLD3cI
dq9Slt+P01hf+iN9DyGCbthNUNnT1wDSnWhUmOG5ous3TdsZ/0cK3Pxd91QuxoLH
PpIw7lqXeECOzzjkOb+tJhLft4muY4+edfGz0wOx6RKhZjt4t6GPtJEDTP8Spren
tE68zsOp/X49dZaSMOQ8XgOoYbsPcwGtMKyx4W6H1DTGgsVR/aJd7NnOeOIoVfgs
MfNEQAAuYBALxvBQb+8Fz+7dtrFJxLx/4GYgv5fXebcXfiendpD8lL+fmgIzqUg7
SkXs4YBpFqaKHUIGT4m1kOtaWj1Ph24cSVDimrETUExFibGQagYWsxnsVKK+JmOP
KVcHNj5udmNOWje12qE34N32HLk7Ozb+y81VafQIM32Q3ehF5GJ5fnxXjM1ATST+
Ikow60Rsw+lF1Dma5JLEPVXKqMWENQmhwoRcJkdLqhJAZU3WSrj+kdzR14069wkk
UWL4RasEkCmPRWQUZYPnhXzHe6ovAl7QQ6EGFN9PZVOPHm8rt4CnH99CzsFkpwoJ
c8r4T8wux7iI5ioQ1hxNARAv2Ez34IQvrcWTRbtK5iC+rcb0u74wk4kO9BKZatXs
e94zpt6zXXgLgTRt8bM7ZLPPtquyqg4bMNHmm20PPB6Ap/byCVjQFp39I6qz7TiW
WHaTf0ziWNlVeJ6df9KnMzS256IOKx9ssiTpEDHMzNlaOnW9MEK+iAafQZT/H3ff
ompb32RX0v8U/cenomKegWj8izsQfZUpnpGI9m/JerqAzdMaiyDEFSUZbW6kGK+Q
/CHFAJqG6TtMWiO1aRV/BuyK8vh3WFejZ3EzB1P2ifuZMwiUDdYWPoT0UZjxpNgX
ckAhJLXCUNTk3cSoMQo1gFooCpqFCp9OJVG10fXzihszkPVjjLGoSc5se0hozwhQ
fyxHadQP53Xv3KcQsRk/1e1ff1POCew8EH2blRUTZhJULrGvUeODsr7rIZgSJ+zw
GSF0zA/Agljpe0Jr0AiWLlbJPRfY0ZSFBt4sq5fMb8F3bNAH+Kp5VGbFLD8eqmCp
C7NzPqzYg9dvC2ef1zlqAWexyTiMbwYE2lRKYgb3+F0tRc7ZUp+0gaXZAXZLHpjR
a6OzxctkgvtnmMolyPHo8+m7E4F2IENRr5761wHenZQvSKhhRFvj3pBg63N8CEKB
lc1VTMocWsnj9Y0eD3ISzQlU9CG1L0eTY3QS6+RH/+bntnh17D9xYoOJe+z+v4i1
hb2X6Hr1tATCBBO6MuZe6sGI8Ck1f4iS1yfUzKRUIZsifQ02WIrNO3pWBl+CrJnZ
9p4SJ01ebhFwwbtmneoaTnndonbvvNuQwg/mvhq6E8qrxQvjA4uM4kQ3Z1EMhsIl
o8FVdqxyb5+25Fu8dIBRsozelzfXHfY3VW54/BM24xRI7xMAsanZaAz557ZcTDtW
9CX/NVBNASuBMvgOrTJxS2c578F1/aqV46c9t1GLlFusfXmmsWEURmUuTfvBzeJw
6uoSXl/62v5YDUzAYQXMBQVjAl0ZGucM8+KcHuTm+kblGTW7ZG/YD1gQ+uvMavC5
OMYJGBNbSHo4jsTX/tssvzhmUWr/T86JbogpYnfVElZqRnp5gaU1dldb6W2jN5e2
oNb/582+X7n9xJKBWSSPLbXe2r+corU3LKBBoompoH0Y/KXMKakKBxCmOMCmKRdR
eX3Ls9lF0xuu5CAlsSqUTgisdC+Stk1+doSh1+j1cmMzYP126VODBLHeM27nIV6K
wCX4Zn/c5HZ4mev4LHrKVjE7dlHylNfGQczTrDL6gmYhkWhkJf2VtueZo7Ua6w3A
/GoEV0XLG+SsjJ6dnhAuSLiClRWKznK/wpNFY6hXKATjyveAnIKCINW53M+xKHYU
VvGq07cWX4ScTIpic8cNXlhJ2dHTG0i1sN9VRhcmgc060Vly1B0XkwpcELEOh+77
0Nsg6fVzNmfbWItSgaOTIzJzWAdt+WRwS9u6Qc8AeZNpLnfDrdMWx5iGsVQnnGqf
5RNCuaz7QU/oGs6s2E1OUcmT2elCWOmP337qgQo/PIwSmd4NIXvi63yqPIw3sAsA
JNdu4UONvx1GQECg9zi0dP1eZmoAps/8G8VpaXreaytDnpravyr/H199Oc69xGKl
GQ9FQLqylZiYh0ZOO4AmlXB3tIlEq+7SK+qkb5Nho/3u8reVgPQoy+7YqOS8W1Lc
LL4vINH6WsDY3QXra7lYuwhiJJ//vlxKqPr8AZ21Toe+ispZRySYW3L7av/bNbr1
WNq/4z7kZZFk4xt2usXbzhbnEagJ2aEGb/k5Cn4ZpS6UNNJmWdTvl9ksY10KVtBM
KaPYZKJkx9KqmIRFn+b+MWAdtNcyFqWEQI9hJ32FijHIIt3JFJBg58tQASCdicF7
WXRoZePnFk5llgAmRwXD14TNwnLAwkrq5GZVKJXo6ulGcVzM98inxTYe27Rz2aEn
m0tmgXYXQkg9V7IU6eWadqjvk23udJLENRmYpShwQoAFSoZu4HiqCCjTrh4zRiXn
ZPG6FslKckb62wv97pxW/2YmWW4naFNCHulvl5UsijGswIlxABUeXCzOvoTAKGC0
0pjg9ubmcAL4SIDhqLJKqSorI3y7eZvNJPeLUIbDWcJgbppZzqoPJ+sZxNzKJpDG
dRPms/s5lz2Eiokw9E0mn2Bv5yv7Oagcc/6lfuYpY5FDmhBzmKUZb5okN071T+Ct
BxqRKVK9+/bX7PG6yP3bz7GYrMrGwRuhT4Hi9X3QP0SdC6kJViOVSD8FyMweUZaf
TCQxefr7U3nDImuF3ykzBwJ2786bpl/JJs5GSGFzZ/oI6KEB+WlcgUVW4Zm0IpuR
D4WG7FVUFsV068qYVurux15/JXMr2TDTknR+6drb/EeqIJnvij1s//W3Mk7QLw2u
7j+88NTAHF6EMGG7WwHVvAkyqOM4iB87hT65q6wBVI5b7RVPVDdva9UeDHoXsmym
GRwghtdgIZKjLlNjq42aVdtCq+CtfIDjcsI/1UiJt+YYmAzAGPPMBcPvwMRbRzky
t0LrVl+BVv7YkSNGIt1MKLx4EwFBbxI+cNBxplKtfLO1BpGaFLHYr80CSZaMIH/D
PyCZBntydsPPZJ9RoIefHmaX/N3BaOxIDpo6nv9N+j/bhjr7Zim2N2lC08FsfZ0M
jfLUfMzjaNOyA++zlPkImv94mEN7RPEnJERsZJol1pIBurMx0ci1buo83lG04eIh
4J6d5AKOTyc3eE95zlanuOFg4Si9QnTCWNhG5U6rxedwZRebcivwxtF7RzM9cFK7
soNeI0TPqBH2Hl0zpW2WOpf1cxsRN7Zdadu7021DLSyWiTAi+shafxTpwt6VwxET
ARCzHM74H6p1cYmcGJQPd0sbx7WTpC6u0QZirIpEFqeksjTcsKG4+4kSHYBhDV+d
PVZmfz50ATVjVybyMssIJyG3g01+RSDycs1xxcxRzfl/4JmBQuJDCSsEU2N+CMG1
Nq3LyWj+QPUxhaplWXDfcrekAmk7RwwKguCK8TGmK43VCKXHgkTQwDlWqeTVwx/v
PQtK0gemQCHXfM65FrQ+MhBOkktaPE553M4O69yRpulpFxY+WJajxtP8luRvk2Qu
5rBeoUni9NV03cpWgyVnROluLyZtik7cZoB/Pm3H4ABABcaYoJzYAUpIEjzOMH7S
g0/MpwvWZFBzsQED1k+2Ap5mNGH8bwLV6qV3JVGmRvCplGadbkAp+JdiZX9Q9QFV
thRbZn9kBIpC6RYGHqfOV/0R6w3146N2UxTqKURQfxsLXzrtbjXvOkLTIbpLf12r
rft3hit2VGaWcTKbVB9Z40Yzn/i0fIf8v/WGbgK/oSAFPc13q1jp/C0x/Y+lqcKq
wTr85ofwkqJdNboyCs1W6WyCob+CydEI4Z6xYKRLZ6TI+6WeNB/qMP8n188xhNDg
JN+qYzHQVsGkgkaQV+rSoewirJALJ01XR327SN9OchbmsedPzp+FaikgnqGhWjVC
yoe2eU4ToCt5oBDrrcBm2pSg0cPTjOXiayYs7527s6+QK9qSac6eizw/qyFjjnFh
q9/zGLveaZ3/2lBkIPNEEBUkFmunnFTpuRuKEiSuY/Q/6hMcd4rGS5mkLWnftbe3
yHJp579+Sq9boMJDm6pULQScPUvUDmk8h6mt9OXjz2+jlUhKIr8wn2SSbHhwvoRF
vD9i0z10XM2Rh2F4wnowuZfn2yWdM21jZWpwOUwXCUawQvUawutSjheYsbarEUzq
lh8wXPlcEgiCqHAK51IEh6+AXVjZZdjPMAID+87r6WsrtlqrTE6H8pL0hTdXhtgI
dXk7VRGZORCOMi0I2TYCxmjk8bTOygwcgADgRH55BSsoF93YGBdU7sR4krxdqtrD
wNG9Mmv5liwdxUQI1s7lNjIiZe31GbHu08R2Zj1DMZSZZmdKXoGojZBEQVPQjZ+o
uAAQ9+AcI7Jc1gPLQcc68UciUOuIZ+qefIzaQWyJJL6/vHP/82+6WI8VN1ZeqyRT
ftxg+gbC/akOd2cXi4FZ0frPer4DjhxJDFMIEEh4OA+gHWMowtKw2aZUHLG6nH3C
LtLB1QQZXDCnotrHxKrc9aSmd/rHHFD+AKcpf/PE9/nNI4w0Nw4YPcD64Cn9eTq1
XChV5r8vCQh6RMFTyfPM3NfFwJ3AOsR9swc79FvL3il6rIg1XmZJw7UZIMInpSNR
oO+1mf0B1UEf3rtwYneGe1NfqFDgnR+WhLBwFXRWOTPGLIIfM0KSBZHbKFmNy7bm
aCkZcG67YJFcqlnakUmgSZ44ZEhnnq3H2CbpbkA3myUA+EtIKT/mQDgoplEQj/xI
iXIHagOiN9q0pTmn6f8o5rfVEauuIEcpJOeBwZl8KBnNcdlEcXVAeQDgkyYKdGoj
XFhkTIu3rYlpwI9jI0GxStlEAGzYqmDsMkiCZmlSFtMx7RtAWAOubqbaAW8TRjiq
+A9s8FIzkFWqlmWTP/2vpah9s/RzHSkFy+kuqBDpGgRQox3uazvhqjsB8NcscyZZ
Q/W6YGjQ0485RTkr/CZb0kHe5cL/nMaEg21KLckq6AkHTJ5FWruME9u/DmEVlhPn
YUhAHyCpLeS0NFPErMvZ76i06/6l40iTea3GbjvKIy9pWhK8ZuD514/gadzQw2Jw
53RSQ9h7VApdWNu1AAx5yOJH+uq5yBtCB+BSFwPLpX3KKnKFQRDzlrGGwpV7FEry
+WX+hdd+HL/K0bXmJzHDoDGew+ZaJ1LVft8+QU8YfRavGFhwIl+efyuAyqzQI/vZ
tw7TbqpzET6O1g2tmyU1qfuoXKKnxVkAMI90bZEILbGmwjpQRfBww5NDsTpu91tO
UZl9wx9+TyANe7CxDPMLt1eUaTW9L5tH7faNUdHdJAlkzhaLhgypE7z2v6r+nABZ
YyGpTl+O5OhCluKNSZTUlH79K8UHdYlxbxALtU4r403m8mDWlM1e86ruccuM9h9V
MYN5c+vih4kGfC7y9y7E1mHpx4TzCq7CcxxTeIgwqSqeSM9ohOxKlvXhhS151qH+
g4A7ZxMQFI/X9uyaV55r21q9T6CiaiEgX1SRQLQRF8fhLrRSMlaWdAGoHl9JdPHF
0KQVHE3ZoiPktjPxXEbiAp4fobVMhXag4Bpk1V1kNb+2FA2kG527edlCXzS+Rdnl
nZd+Cuo+wvh42y064wlGDsErJUV1N56qzvm7L8o8UOvz+rngEy3/71D5ttku/dhA
yJMIaw+p5y+vczd+SsMYvotY1uOp0PN9saAE2ERYuJHd//CPsJ1xPemnsARD5asC
/g+alwWSISxfC+zmudEHa52IZDGpFUx+3RwehLAr6BeCwaoXpvyb5E1ngdSujkOQ
PuLhwFoZPLIc17A+j8Wc1CDcW3ucVWcHqLPe1SGwZ2p2j+5jD1/7EDvjLVryKpOv
g87MAUHd+gska4NrxSPTPEd1ZaDqjso1Jz/2c7JTdT1SfGaP3bCO7SUv4uc9XmLc
dbdJ0cxWFvMQuB5fEFDQaUWP/MgZbZxgOhKA47ErOMF4Pcizmp3AR+UwqoutaZ7b
A1WOm9jYb40I6RUYMdR9Add8GarlVS0zOiFsbswIJ3GuUm245s4bFbIykdBF3ati
0uKLumrwuykqGZ+PYlMGSYaS6gCZeVNpvpA0rJOMVpUOQAAfv99GAhHeH30XK2+z
L4lqjkQI9o4fXZ1uHfLtLJPzJ+QV10Ft9ERIpY10zT46z8gloSFsmlYvU7rOEKVs
uh72zvm26Qym7gEWFdg2neR5ahb7yt3FObTLTSEDg/MOhqKa2RODa9/WwLdvya9x
3hUgTh4oRZl1K7EhXyTDFz0VNyrq8/FuhVMkrzfdlZlVTG1mMJ14FJMBAIoCyoQY
y339IyxY3C1PLK4p5ZkZtjj09T8FeVCN0BLEXkJZAEG+aM0lXmnUU3bOzWJOEtdR
P54+I1ho+ANQ5m9yY7FU/EW7X1UFSYXcpLlgiv6FRiZ5JsU3NJOqKEWqMKSu0Md1
5ietZOOFmsN6gXk0g9FLyRA42JQhYeZBvVJ7hh3TDIrngjvYl6yP4mwN9FrqyPT4
IuHxTG7Zd9xUD0YhEkq5oJeJgC2phJPAHXOKy78ZrNXIKteuIj3WsTjfzJnBOxbW
UyKIjsvXy+UC4W8BSbH4n9G/FzETS/UG4BvsSMda6msU3hRuJPtMaoTzCwiZ4DgW
t4YfdeBamMks5V6RKgG/Aki8OXjxpA8wdKvX+0Ca5kAICiv6CT8ZduNLhZUk3uj1
LWSblmccLPKD6W2JLDu22qSWKtt5brG4nsybL4AhdjrDCXqtrj+L0srXA7V9z42w
9BQ5V0NdVmW+mS0aMxfGfmEcufvSqa2KAlKipWcXoTOFqGu/rEK6XgUeknQ9Edd7
lvgAtoBEdzyqsgNdEveHbAS7LFRsWt/AZBZe9a9Y4ZXxUQd77awmnFa6+NOZRwte
eYmkHfz4+7sIYENkyfjf2owKe/OUSmtQ1RR9cI5aOq2D82bmIPYtE1dxk/F7eCEJ
De1CrvCNb39kDt2QFC3dQuDM2IUGKULcJb62H8bbr0bJbI9GQsWGKIUUUkILXkw8
fH1SlUWBcDqCM+58Qh5ssREQXBLIVjM5l/J+dkg3H0Y7nzI9Ag52F60eGke93u+6
g4hdKXiJQe1Bc0ISAPWuWYq0Vz2CKLEDEWg5vaPvsfk5X+sTuglQAsNsoXIQjSga
x+/p1gTOJ/wOJ3/Ys23sNIFXh0whhaqAUcbRyUR98vHCC8/KrBLHCHKVB7nd0NCu
+1XujXqreoTGjmpHu0a61A2n5XxRb63kmllyWCZwtxiao1C7Z82s+uMkDmYZy+8+
Ays2d2ShTZUr/Yxj0Ka0sx21RRtVL27Uuy6jSza7iLoEDGWqG2f3LhHVhc6i1vRF
yN+KJCdVgn4bGfG11H22DyvJqqlg2aF/7FeX7zfa6KIolM9eM2aneFW6YbiObSJT
ibN3/hiOjOUyfk8vHOZPsr+i3rMB+4pylU8Zaf/OEVaLzHbRijWseNviS5stN0VM
2BhjmBI9l9RbEVjTgyzUJx4XPHvnK3bgK3fQTae9tZ1S/cHyG0ZqRQLDIXuqDG4V
fa28srflEn0VGza8IRru6HZGgJ8ejxePwpF2x/wcuR18NCXvFKRyAcsINDN/pVCx
7ZYG14ByYu4H5X53sA4SjVJLi1rxD6gTjEgdITNM5BZjh+hTy8Cl1oK6jOoTD9l1
rKzKlTQOFrL7exKlOe7n+LU83nnthutpe/wF/VGDO5qdfG+XN2qSLzcMk4BEALUz
espoRMdjmnh4azYjJvapUrl9Mhfznh8cVPvBOeMJcWuFJFd/wQqvj9J2pSFgOfxX
km2p5CRG8170pRBSNHSCFyuntzxyb6V15VmZCxyPUPuTg9JvpRkrFrjh6FRHvfkO
D3jkERHW7UWs26hsOR156bOxPyAxsDxwjFYaXjHkv148D8ZIoAO6v0l4UYwhhmBP
UmtWNNYGMDV8ONOAkX3d6Qp07n3aIOpBzryQ7iI9n1rg7y3dlRwgTVeUNKB2cI/U
UTjak59G6aX/jD6t1/DXiXCDmQsb7hPsC1ScoPIJdEkz2mw8oxBSpIW0T0YHrGii
bL/kI1wxitz+q7HCM9SP+uCoe/oTXH/ovqFgwa3cCC6Du9zuIbwU/vMoI2iKpwZt
jjjSgric4XXgRKIe/D/H4H1aS9Kcco1GDla49R+2qa+ax8eAPzdgo1CzjbRG908I
FT8+MCac6eVAH54zlq2em/w0MoJzszdq4htIw4DMbIJEIlKfqsVPeCDmRHXaUHyp
q9OkgQZz+cc78ep9zz85V5DndAwByTnxRnhrz7JBLhiZO8LLM6K5Z4QimfT4YOCN
CnsUIAL3hh75eU3cbbctBiP0zwc+xVq50E4zG1NeD+4i52SyPlcr36j1T9xnj7Yc
eQ4BI9Bs79F1AE+vW9Gvzu2uHxGzJW9hHpbhRShqphYtaOolAx3o4lPPERalt0eL
nZ9lUndRVm7pMNfavZ/8W02TIvvKDw+jbzorJYWuWy9vjoH8z3fEk9nqlC7CSJI2
GU4Xh1pOqtSgMm63cSwIGdqZVgVDiq251/2cCrFTzlqep8RkBU2mVhIPjltJUIw3
QGJ46fStW8aukPbV/M9J9kzV5GE2+VpbTR2Yx7C/DlmqbjkiynNXxsfUJxJhssjh
aM3SMCNiLnZWoxJQXUqKmJWK1t8FtWBFXhW+6Kbet/v0Ko+cAE4bk2nhhgT1nxKa
93EJyUPcbaMl+gwK0T6Gl3JxuTlu54p7vWDxr9ruit9EhNE5LVN9+GFBSPFLx5tR
96cGl7quEwIqLr+6qvEbInPHSyv6qU0Z63mMda1jqirk3qlFNH4m8A1GRzLwt05Y
3EzviuAyYorfF56vMu+0n3SI/O5vgyJpZMXLqvk0bwspX5+LQc/9tHs0Xk+3pIzn
amTWbtWrqeTOMhfRozBC2tJzUR1HXBp7ocIMyi2uuGG8sf6MvDrDB0Nuo9jAeHvj
i6VnttlVt/zhKOxQqobsuEnkdQbAxkQtGYoxEHcnvGP0Q6KFrQO0V0aqN+ZVhx9S
Go6V1NESko6nlWzgW0RY++eHmPUwPuaeqVxMqQT3bqdRXnQJNgBq8rbKFwYdRGR0
RJNvEzyidBrfnA33jfjAlAaw1ENNHziNISwKjAWMVvhLrxYXRTbcWo811ITLGKlR
1aVEbplqTm7OCdd1ZcK7dXt9Tw4iGQRcFdYHKf6hHqjQOjCRPDeESvfEZk+k6Ghp
dvDC9ggVXBw4rOnqKONc+dKCHKU5uzvmfUXztzAfRMYjKZg11FBO4vvXe00C0RhE
bYDygXfPvTKmAGH7Su639s2pRZqlPUc/xFTf/yUU+7V+QsOuCQ3FcU5uPFhtzL36
a0/kr2Wo6m+GL++013ETWO1Y8l7JoRxSuXmGopR0375RjCPwOPpf5RciSeYcW3UH
Le1WmD0jo35YwzibL124M68h0vu0whaKfuqaEUPAYXN9Sqrlam2z+27GlG+wI1yd
MHNcBQHKwobKLqDOSr+w+XMZ32fdSRuvlA2lM1Zu0uwoVn1Qk/PceMiAQDjOysMG
qt38OX9Tjkk2hxcsWUNWcYLl1gVqaMZBw69la8+2/uiRlwAKqIOgTMTxG33iTuKI
yc0eyK9/XqrEkrjVGwbO45BH2W3vIlZ1yOeP1CuaodBgeeL/Wf9ZIjLAYE2t1rmS
TNICsnCHZiNaO79WEJ7l4lRSlpWHSUoKjyIML/yzhlzeidAs3ncVu0Ap758oFKSI
LG5kkT7ksoKDPB1MRogvMZ3zipuitPDWX1KNJsojhUEpMHwV8Sd3dPFYjibWx8gH
bYbgqcUkGfjLmrowbzeb3MUgS+wRxQ1Lb+NUa88774d7xYmdPeyDwKSHWAhhDBRC
R8PSurnGFUqnwf9OorsKhwQ3Kmr69XCICe0n+J5u5aTU5lyXA578TGYALLQZBCbr
QdFW8zIXD97IQWy8EQnA1AcuOZmIxcCnzGDSyrAMjScGkF5rU2F1VJUq1BplhQER
Hgcn2vuGJOg1p4RK9vHeLVp0wNleCFbRYTQP5keos37BZn05GPsXzTnJ2wv5tCOH
WHjjpsWvDa5oFbv33n43RPBLaMdtogIoa+Hky4NVazDFiEQcN9CM6fVxtm8/B5K3
CVvz+8tbuJV2gyrb51UABxvSXzUa66aHRk0FSuBuHsIfKIQFfZfZqz4oLIavHTpg
vpgytp8AUtLNRjhiXY1ASFfZaW+WcSm/dooOLjk6iRBk7+RLMadGT9P7LQ3VRjsm
8WnBr1O0bwy3sA2ctliqhOgrKvJihW1KfMbjnj9N/ly8nMkLXItD0zg4AMbSKQ6G
IGid3f0NRj6gIo5yWcfmvm1HDhQV91zSzieNRwauFNODVvL3visNkbobu/hAxLUA
+M8nwXmeIlA+dhbmYnlFTLwee0lvVlrqlUf4UG3tWKG5xjM3uCdIfwJF8spHeyJW
bG0fl/1rOezYLJLrJGMorbgtvXQ3fBlbaUItk5gONHIdIl8t0PJ3q5ikNKoLe3GQ
YOnfpTyThzDFdlQvpOXSbM6JL5SPhPgamweJBXoh0lF38F29DuwqL0E15rDyZ+y+
D9E7+IPfIFRHxtKgCJ6hy5eRVP5CiRh8Bax6eypDw3KdtNmGoom1+eHiux7KJG3I
wkMAEvmH5uP2MaJ4j9xRsGlGEB+cyFBL0A5VJpPJ2Kelxcmw+SqaAw40OgoPPmMw
T33hLM+CgaP7ueSYl6hnhdlB+OkIrOWRhMYCykIPOrK6Pt09de+b12xdEI+z/cun
zkRhw0T58IVljBr5Mu8lKERwqu3XDbcfiGKKrBM1CFwncl6rf16FAeVYLV42K72L
t3hTQSA26zdCnR+lDuB3VxKuhFMHUeNA3AeejmvYh6UFk48ToQgRrkoOynp4cnAb
cYvFJO/1vCEd4UJNfsgWPGvElv9K41hWAswuG+0X6QVlvg/W0usDClUUlkfo2IPo
dhxvP9Cfby+KXbGsDRChUlgbFgAGBD+B0MuOssY5HSEy/Fo3UdII904fCV1mypN3
UZGu0xRC/UHcRv5s2tPPmeRqBskSHOJe9CV2sd7J8iZL69mSVwoPPXZWcIzbdYMa
Ky4Lja5iVR93b+XbYzIIJ3qSRiFekwq+sCdDj4eIAGeT4lmtzm0WpIFrMd9qF6Ol
fnnrrmFwSRPliMKMEcV2hwXBncZKh7xA4elop+EK7NFLYj+xCvGJ/9VZbJ/UT1YE
1EE925gUWyz4Zq/9cWUKAYnvd8QUcuL5GTrKN5sTV8NeqQfTZA+kmIQ/BBJHn+QG
7qKj4aIRr4P4eATbKJPtRLgTLT8RI2o/fCTsV/ZMOhdh6wyJT6IthpjthPtGuB/0
Zya0ppm84IL0rBNxBC33i+yJP6fVjzk8VUx8wFyBwE+HzwtacRP9QodYTPlVfGEv
K3BgmedNfXsOgzxbuYAHyqsyW37cqUtVCqrfYah9rGIjmfUk8Uo53Kdyln9zKQNN
I1Zs5eqqefpbdkoceICEs4fY60PYqQf97jhTZkLQzNSxM+QtAVT3tjSFdB0R9hHd
GVUB2Pr3vwRSwJVlfsGTCdN2B8CW0pGG70hvwKthqNkxxFGgiEe9OUq75MHrbLpR
/tCIsJT+S+uuvgZn3RFn2fG9nsIJXh960nE8Hqj4BXffKzt3kKs6oaUaTaeVkpuE
AEkzCcggVY/GeKY+bFPm2PfY1p3ZKY3YXqyjhRM8ns99mcsYRO8XqDP+BLsOCTRt
nwjYKhEBEYOCIuhDnuCPOdjKaDxgO48j42IrUTL5FVjQP7qZq9tORaljGFLkrZm6
zPSTO3m0iWX2btXFaPyv5AkLFx+/glJnGU8LerGyqgw62xohJBJkyAU1FkQyQ9pJ
p0L1tYBHXa0E16Y2S99ZN0HSTwiKAu/M4TG4RSdFPdY7IzDKHIdWqXbZfOwy3VKI
/7y+TcbfFU5mKzS/qbvzSa5TYgWUo/YGqoiwb8rxCqIIKSRPnH/I2BsqL8B0A9QC
M8hgRugLoAD3iMURTV8RaqR+hTJUxLOA5J9L/2ZPKB8IX/CKLZl51sPF2mo0TBb+
sWj8vnhPTEQq9LiX6jys40Nv1XGedEZ/bq/e3EfXF7WR+pWaEDr3LIGO0JEM45de
tYbfhJKP8+4/LiDLQyaapSkRwpyupZJlSjS96gs/vO0UMgazJd0tY1qmXwcB8JWp
Hd/FLsBMn/2554G409GFDaThpQ4o+7HvaNkeAj3zsMCMo8IZ8zBWVG74+QeFietC
6urE7pa8VUfHzgNgikXb0qW3D6JL7hKfYbAD9nvZl35vxcZms+YQ2cMvZbyjMYra
hPIDKPdMENtBpBKZklzZD0Lv29K1WvrWoNe5VmS/OJUB1+i07XZfISmlPw0BTaEi
Xs0m1Yy8NRRW1/kOxA+QlAPlC4Onzm7i+jD0lNUk5SAVykkphuXns+ESO132CuBT
VgYh9CyN+hBzADCOVUTiAlHCg7XuIK5mvvSLAyNaiW68mIefQ8OMhsZU5V+V70gt
tagJn+0dmEw/R9NKpKjIgpWEHAg5xXyolljfakuf3KcQqU25jISvVyT79aNL0ZoE
DgvBA8ectywYWHnqUbowYOPUuFvhkwBbxfDrxB3prMhrRfrXZBsgpI3tWNerSmJG
6L/L8BYnXpR9lWb2ors4K11kbgHxovH5DYmqHWlnlMPpfoT0ljUIXUPv+cEfPN43
a3VU4onWvBMefRg7Y94c71EcIcVS80SQg6cnJgEWa2AErbXBceRi6HbYnCaKPB+N
8uXYEYmAefYVCGf4WbUoS1cBB6RB3es8tZq5U7ORnforZTkeawO9QFLQZ7kkh3xX
jP6U/0kX/IZ3MsJqSE7ORCxbcI6h6UiBtRR+reynt6JvbHab1dqNf1L5+LLyIjCH
J9wsbhb5rCoN19xWiRrYX9mvCY2AK88/qPVSRzbO+3fyJ8eHQ/GcfLGY9SDW6LEY
vLWa77ftlyfThpDjeFDIzGNNLTBYnUGyOdqCd9ZgDLbKbL+AWwpIztEJBD2m/BSG
W0Slok2Lxt3b4o85LJjWtOC+uiEx+KC+5a1dhe2W7Z8DxlXOWshzZxh1rEQClLzc
lkRsNorMhM29OUizch2ViKukjSmoUlTo5nYUfGlmvgbC/PQgk022hXT9CfFNDO/0
zhzToNN8GAhC29se5gRBv7HNqyKRXPI2XfHPd4YDKCvqnxusXMyoNj7PIT3R18EG
lLw9bwShAyXNgCmnuVf9GibtxNX0vYDgqhd2oLu/y4g/Qwsh73fkXEolhJ+2NTfJ
M8o5Qzf/yDrYDqVl8IBEdXOPgstxFsh7Yna+DjbnszK5MBgfqUdzNXn3F4wnd/aP
P3rB2cCLHzwtM7SySzUWUyu3oD0SBgemNMBoHtS1EujQFOjeWlWydiqCDUxXW2xw
M1EMD7HzPgYMnkqKA40DgQhqu1rWGOW3ljOTu3k1NT4Z3GAq20KT763s7Mj2IV0N
EJ9L48QvXIFli2skGBxNqxdH2zz10MYcqa4TpYcLI/M9tZvpYDP0vapXb9HbMrP7
VeiVvCbd8osHtXhv5BC1/wWdIs4pA7bATvVHxaQReTaC+AHXLxk/4ai0LCg5ML+a
EI68OyacYafaoZEPCTn8VuUZN/Wq1P6vqcprGCx92t8S5+mMNE7Fq5LvREYR7szf
F/Q3wGrmnUWm3H6y3/zux5ty0n3A/lsyGYcOxFkop6VoR2h21ydX0AqLMWveFTSx
ZPri3127Tl5M4SkDApe7QgMfDELe0vxsADXPhuVAtxSqseVsZJTByxoPBFO7Glb2
WdOorz77TBkQMi0jTsmIj6x35pfO6fFZ3+8d6Sp88erPOk9vh+q7oArT7Z6rgYtU
Cm8K0y0g9EE2+WvDNFdvWEGQW3g+Q0OZrD8GDNRyL1uCicUia1alXhQTDATh6TEj
SW79FN1wwOjgDeL/dcjnSWEwz0Eba+nNXERaadjNfow9tkIAz1ecwMQxKi15DFbu
bfCTstkvR/3JNUb8r5Dr/5IPWlcyGTYcaxi5ISViHKh8QZmZRYYP/LEQgSOh20gT
jrhQ/s0efIypnPYngg3WPbAbEZZb6xx5um4itZR9TqQeZwS+Fqiw/Z6DUf86H37x
dhh+pkC4rAMWoNaac3cqaRUe8hYkuR+wouyoVBcTJvd+VpYxBB4ml1m0dVlvnJ8E
91IE2wqYRx9gSWPVaV4Tbm0ROORZ8uDl+z2q3e9CALne/wfmWmbRYhwrNIJ7kQnt
LbiQ7TnR4LyYr23sp4EZlaWsW7cocUTY/mR3O7BHf15K+8qERi+2RzxEU5WHg5Bg
sxdMd1wwtSwy9i9g7h1Hi+MGwS+cY3RMwCRi6MEeBIjCaYHWWS8hSmO5/SD5q5AH
6Ns/HygswoI9caSlnfnghLWg9QXZZ+goo0zVKi81YFjX0GG6Gg2kqef33bX3MLGM
W9mfmQa2k9Sp5bEqd53zVyGh1fHA0HJZjeGhrQ9CPTfSCOIbFMj2fd69lxv9Giq+
N719W3zVdCWRjo1KD8nVJG2yOJ2m+SJ/7C6cnSIt3WtmttchfN7/CB4jHg4EwJ5n
tk+GdFcmHobxul0R5JwfuAc2OizDsKxmBsLpJng8UFYvCUeP/HPHLxUV4j+WLPZR
sSF5eDeurV4md2tb87kuMkINpAXlwm0Z03jAWcj7sopKpSdvxnKeshhuvwb7zjdh
6oBtuq0PNE2L2QEJKEdy6SzToN4CpnaIub6NHA39tCCpG0QM/i0P+m3f7eEjkquJ
4r1Jdlvmop7nJ4HyzP+kRbcIHztXnSMDPXUlHuenITki2sH+IoyQKjozB3lC/ywM
0CX/nuDf/nStColgQIbVUFJOyL7TFSVQSPGZdL8QoNBqVKsrdw+DblMRqz/7bkDH
yYP392huvdg2wvAOiWh4ALj/q77FzKCTZunxhijVaZ8moMqg6PcmIgIbN/P1rSs0
HWQVYd19lSyl+IA264r2nF8bXr0mp1RRAezShh8Ep6ZXGEDZF4pj71zJ0s7+5rbM
ppVMXvAcJBtevqH7lKubjIAEZXrcZIPzU8KuX0r5RMol1EWm7LOpIX21aF9d7LLr
VQI6RYyoOIxN8oBrmlMvkkZPTJDOPAZMKlAeujSPWh7LlJbA8wRj2Xvzhi+PYJGY
pBjnizU6msPXj3P4/Z0XDT9BIh8n5sQkZPpRdG2IckJUTjyPMekn6bfuwdBkVkJb
Q3vmkbtfbBNNArsXW4RSCtekqffv0Z5iLkc1wWJhq0v+6Tu4VAnKU3f1ijC9/iIB
/mLusOdh8+SJH/IwUkgPzh+o3J7MV7+tgeVIGwKH8Zekcwv9OBsaZCVYtWsIH/0A
tDVbhgNGOdl+O41DCN3WpLLG5VgyAOQ3wwFDpIvXKP69FwlVjPNUlyHRTx8DbJQs
brkhYhkBuh8xpC2iu/KnSPB7vCKH0C40Jg1CUZrSkIIx49iDNgdncUqb1M9b8MtV
mVsmPg9DJ0yWlEIpUu7v8SSzgAukTBkJX30XrcEG61Jx02uYtGibxgeHemvhGqiS
RGg/Bj95J6vvn64nvFeDneyaxlj4NmipGwIN5fagdZpjB8Wec/F3SRWSG6KB0R1F
gg2QXqjrINYK5/zy0wgvPIc7HtTzEjxh0YRwayheVfJdLZ9CN+s6k3i3baygRG0n
nqj7kd98rjJdtm9Ul8JxT6RCxsQT3fyp24y825CttAFDrYbvtmQS0dT6sTbKeRCC
Vh5MITfcwcdA4+Zqr0/lHEsvn9xRA9o0oChKIfL+ZhDEIfyWFFNHNB60YqB2DIA5
t49OUhxcvEDuUZSk/Biy/4WVXrVOO4YwiWYa2JsAzoZ9pynlq50PU76ih9Q4ycY6
iprgjhNQKtTv0hF3UoQwg0ogAuYhOzVNPtUXq9EoRkzkYtmh9iuU0VMeDgTMZEZ0
40W2sIrRnLqkUXbNdT37WBGaod29ONBV9IcHG8uEr9eqDSm9K5vT0YiefJL1FnEb
PpG1487LKLei/BGbnSadAIpHnTvgLiatAZINVfU3QV3D3h3rkR/+gDdaMXlidNFF
zvdWi+9/ggtTww/5eFirOqRkSASXNuAHMVAQiJesWhxUQs159C4WEZOYb/YFdayJ
VfsgC/laDNwJnq862dN7bAUU1aYINchWDN6HzJb4PgTuQYusStB5K1SyP5qUHk7t
yZyelr9qjFuNhF9GyHXU7YLgRVLK0a+/KZwPnJv6LUTpttwHyy/xtVD46FMj50r3
XdXXOSADPLWPA2z1QSvX2MK2IEOAt5IbFqDjaF/nO6bNX/6Wo9j9KHvNEFoVLJ9F
oxuJ+ZQcmjmycILq8R2Pryepz9peoldt2RZIz/S31BOR53lZS2SMGONPbkBZLnCW
b8BqsqFIW4LBYTRdYtEHDtlvTu10NAsR+WCRdYrXGxa43zWlatb4hlI+22bCo65t
iWZKdJn8tEIFOYBaaIh1Gp6lFt9bJT4AijeJ5/K7J5+dmBTt0AT2JR8nYG53QCCW
/EePOO3+zqb+JLwvcmmCDe8WxDw8orWCJ96JM9x5Fzu2HxY0RhHi+0B67jxy+U5u
NsSo3j8WW+dD77A7LiOPeyJFUhO5rASx3KuOYRUCKJjm/d9Ua1HXepKFpctNZvWV
GGsNEO+g9hrbovIXKTVQshRS8muC0PmZRGRWJBlbfMsmvkq8Z0QPi/JqzPIF68ov
PUAQ1UXEle8rIKJqdUoj8sMUy+luQK34Ay2z/v2QT1Iglv993Kx09uO1VkWUI6CF
eRa9va4CSSb4Wu/CrRSGLoZylgJjfHXq7dMIpt41f1d6SowiiupNI86FzzEjwJtq
S5ZOJ2G2amiUBUfwLzzx/WrCmt3+QQwf2PV2BKvY7tAjpgcQik/D1SNFxn/0uLzc
EV4Xu+heah4hkBGnuwv0F4EYgizovVg6F1Q8jZ97r8IJcAp5YPXyLPt2HYPynjAw
eQE7c0OJ4Gm4o+FsYOXKdzN3z4yCe7XkhXmXguEKReZ2SbYOwHFVMSFyew9JN7Tr
riU2QiTMlXimruP9Y4DEGU15bW1AKFEvfHDLsKUiV0O5KQkk79/CO6o09QfWeR91
1g95koGuXwkwXwwEBIggnttMIQpfimXRmjLIiVz162f9yDsNctAOZPwzp6GSH50D
0KDuHJGyy8nipEFFeibh0LR3C1qSlmOpZ32icbZ9PXAOGwYE9v/O8h7ErFydZGu3
S5h5DzoJpp9Ccn5J3aCe7JX2hKcP5uxyori2RZPU+B1CEX1CeGcgZ0wpmixbp2Q3
kXz8+8t5S7Evq/BbZBsAub0zhQOICgVHXLP+P8S2+kJfOyoE39pI47/lcSHCmJ6k
eRQ8lI3bvjeieq4HQ7Zac51hvIiorOy2vu28aoIo3MlphKEkNrxOYYxqnvNmJudQ
EifFoZUOcJQTeB5f3Ao4fgUodL7JjG7+ibdSBwT3w31Ttx9CVVLsvjFcyBSrOCkY
mUy50f/F4QbFY7hH0iJQnm4OwvffdpOmwAbAqn3mSRn8yE1LWv3LYXLTwu2mfx0Y
LlDxyJV5A9AYqEGGtohf6PVCyQDrW9robEe4hCEhUBMlPQMDV7041qRU8p29PnmD
3E+YADQwJpV8lmNJPjz7+gnf+3kBSKHvkauV9h4QNkmoAgtGh0gvBZrPls09nJpr
wbQ/3TDYQvfQhqrlrDgAHawov4cOg6CMNEJWtga68fKw0y3HSGxUaDOepvyRxzH3
jbX0DkGnJ53lTYAVZ6dsi7m75mMDvqmPCJoPbjvsaELZ6787vpeArK/5EnP5BXqY
YbmHkOsY94fW06SmiKcAErcTyUijPColr2MHGfOrPJCM36E4LXEpTxO+4gS28irM
3x9yvbLd2PCyAgh85TyTVyj7V90EmrwcUCcthBqqdtY12HjvZbB8a46d9VGsh0LD
KQMioalNhUPt7RsnR6YGbgaxk8Ueu3T/CcfqTvbm4r4PmM3YEY9fgaUt/kFRDN4k
keRVyAOgkUBZe1Zyv1iT3WaMFlaXA9b5VWPtMwlFw5iH26OMgC+VZAXCONxebknp
UMvCE9b2X7F7yLho1t4mAax3CETlcHpV2QHmJm3z5l9RqdaxmRK/NOCbam60MgH0
HlhfOubgygonZ3CFPYgjEejjRrJdHuDdXlYHHsj22sTKO/xh8+Sq60UXzKLOboLd
TTx7MAd/FBEKEZKqvh6Yg427JZNykdKxKwqJx3N0nIkCHMFt8Y0+dvYjgA7TXGW9
TsY1XkTVYzBVCEcHzrFKU9XVOAdQWcGu1gdoM8SRR3XxRiDBcZGu8xopJSCwKLxP
GdZFATfdGT6L4CNFaohguIKKdAf8/y+1Z1LuHECfxmziUbJFZpMJa9Hnx8B1AHvd
Pkmya/c4/d9H/fDJTy7FNNJ4Uvp+XgsV6SP6OSiJnX9+4zHl83ASG0XSD8NNt5KM
Zs7VcJ0z5VUOHev6qBc6ju3EyMY3F9Qs7R1oyrOmYer0PxUW0z3lNsfOpjJAqIJ1
H6YiSChAf0hk9wv9pwwfjFazZ5kWH6OkENHCIr+SrazxE9cFCPq+XLurFRaFGD0a
SCUN+bCs+QBhAjLpLC5qja/9KKzTzePu/zIo5t9fGbx3hnWxdqm6N+5w4KHB8ozJ
phLDNwiEpfm7qhlErJWmkx8sCXs+HhbC6EH8hdDK0cBM6E+FnW/WQfu/IfCL3Dk2
0y5OX/wV2Unnsgx3+oKjsmaVadg0wTFvhljU4iV+a0anhJzaelnDVcaG6xss4W0P
+pIM/HYETGMmzLyO3rz7lETKLvXkY1qUlSsJe4XoHFawOLJDBGi3pefUZ2niY0nc
saICh1aJRuD9+rWPc+7OXphkDDvOmqdgVexHTjjyEiPQ7EKbMqqwCSomQySbvn1H
WriXKBJd50nVHxNSHUQDjq8lwGbAjqK1hSWakAzn59vaqO1jcd3dwQioejzs80PH
44DMl4I1QGO964m8tleZ3IAlWeKdI7MGBrqKkvU3xFkjyFffIdfUg+udUNnIXl3d
Eyua/hyfAaRsC0fcknaSTJFpWWm44nI8kZlvFLrvv2y3XwfeD5RDpttKUAEgr7Iz
0ojwxZlEfq2Hk3/WCNFN2k543lc5RkEv0hd/5TUmqcKbDGSdQrk9IivqlbPMsjo9
EBSJH+V/XhFiZ/IfOagdYAenn68oTCk6msnVw/Or2q5b5yW35A632WWgG0WGo52j
oaEHFydQt/EyUkOzLP62ERhZR6wqUNR39AOWiA7tQz3tAaFnCenxS48dy1N18+rW
RqOUPtQ9L2AuAOVzri9jUY8S1/ZKDntN3GHImoHCqUutCoD6AnEjby/b/WVpUJk9
h9AyWBB4tVW1yTCvpWwh5B6NkpaxjjcJl4UZAtAb8VMe1NsqAXpuZiTFPzeImFaz
zJVUCiYEVOU4sw+xPyzcYumK9kZRrFubFrsL1YMZqSxy5HU1hKIuqVE1+m7pSfNq
RmwKljOMd/GVTe9Th1A9tgeSUcOWqiRnPGbrsLsT3x3dWXXAFDV8R4vsHhbdZ/B9
zjzOlZlSoZPl7XXE1POroIS5k9kufWdWh7Oz18gHzEkmPebVIQk9mkIIRKDSupem
5cHokyyFmQbXWPJC/gOBP9z/1qDmN5cOdhS3pD2t8KesLni08Ob6q6JmgCUvX69+
HRi2DhvXBNlfbt8/Q/JTR8quKLHZqnEKrty9prrF3fEYKU3dB7A5o0TzTGTnro/p
shqjJSc5TGR6bM8F1oxVWUWOlBCK4cVlrEsdXBLdfu9tWPDUAm121T7tq51fyivO
jlyR0pYzbbUFYEMdlab7i3R/e+K6C58v0FvDuYAxejaK7JY0zMAtv3XbJCmxxQRv
4ELf18Mk5mCw8Hv4xNqQijPWvBTe9PF5py7K7HRQgYBDz1yuY13ZGFfduT2CYasK
SDSvfdOKbQwo9jMukSa1RJQ701yrqmjbYS1dBZMlWP+RVgzOfYMAuhAtuIa/Iu2E
G8CVASDmhopuQzYBufszU0VHTVdVIa93PKppffYNq0cfFfFEQomy85vw3Zk6g+uf
pw0AO+18X9NPnq3yS7TtO5WxhRTY0HukefE6BNgj2/kw5TZojgHncM57+IZIyBf2
jeMEJy3rkh2YpmhKWYgpnoWK5p2w8BLzy80BgJKKKGhNt9SCQb/Piki5lFsWyk6E
yNgDd745awTryNRJw1CgyWBkJNU++iQaZ1lBGwmGzoAUt6L5OFAPWQVA6aVzzMqL
7bHSYebBQampn2EvRn+sqC1rONuya9QJIq51nLjswe5pHctbmfXFS3n19d6x0rJY
+hE2wtEdvU1og6PC5qz3JH6O4TvQDcmPX2F/GwpKwtbCJAethPR/6Jsjgjs50KM9
KORWCyZCQN4642wbOwu7Q69Il/ptd3R3D4DvGx+pXVRwy4gPwLS+icXPGftV+RUD
wxFdP+95k9+Cwtp4pdTJ6r5M+v3Q//YF90HLrbQhtK2C2hPJfplLahw8yXcipXic
l9KwsHF5kIz0tVQOcfxYp1kXBjQufPTQXsG0Sy3femYdsKq3ill4B6fBJSNbs3+q
HPL80eFgYPi5Z18RqdOQ3+AdWpIDbmKAw/nKIgx57VlQioA0dnr7r8np5Hvp5vRv
Fk0VsZ16Nb4vPdLb7cufA0+qamWwZuK/Iwim5u5ylzJ2ZRe/NRnaKLjUGRWS/DOu
9pyiKM/CoR2KCe4LBk9cVH/rLfvzPCrDxPmWJ776PFknLkNaEDXbRO/DlqiN08ea
3aIJ5xaYbirKarrgGI7NGkDk150eD+4GMHmObc4wtdOxkO/6fp5z3euyR2xqhHI0
SR9VCBhL5dm7sZmZgiKAMxAze4aUgigwsSoigeLBpyj2YMC4DUj4POjCWVMprUKo
KbW5kfm5uteGi6L8aZkpx0JPsJsThqZ+Tv2EwJp4XzYCuPzY33sXXiMRrMG7wrQR
jyppC4cm2zFTIjL7ns4poKqzuVRGM1zvnbWbJGlG/zjsNNU17cwrmyD8Kx4x8ptF
Utibm4PTwkizrMEl+rl0DIBc6mTJ0VDD8DUrUGgGhl9eRlSE7daUHcS8KH3sKrrU
M/w/TtnKzUedCU7vf9NrLWEITi9y88EEi2wsDQCw7tqtrtsauLGYqQ2ThThDUtNz
GYg3CYo4s8P+1mMybROVz07aqajudepBrUW8It4uJLgQS8fERatsD6ziX6MbneRx
P7ODj1hDC9r7Djfxhrgqze0nlMFA2yVm4P816IkTxQF8O/F9v8Mza+oeZ27Um4Cy
A7aTM4NYaBQKSlm2Bmtzw8rLf0UdeQ/pRDpd2uIBpnx3hGpXvGt/cvMk29iTjoLu
fnzCOu/12PEw7XVzJ4bBv+/cepX1aIykPBdM/z5U8QQns6EqLFmvbFatSuz5TO9r
PdVOar13ByEmaJ4shORXUw702JbjuZffA0v2CEKCPe4qC3Hai/dPTqFUMGZpu4Na
hDoTJZ6KLa/eiD4Tnc8cRjMM8Zz0qp+5ykYnr7/o6hz2wFBxDyt2Nj9pj/CkzgGT
uOt7IuJgXr2IgmbOAWiQGd5KyNQowUjyF2/mCBjgqDBlQYBWEtUaZaYYHRkjAZk5
25xLlknRruUZi54k/L3g7E3z7Bhw8byxNdcVyqXIzC1pHbVny8pLuLourkQF6XC5
bczxWBXx1EWAl2ig31Pxg1/XbHmC6KzGy21BPePiXz7r6z/sfdehzDyyImyurGdh
yXtzG81euMvbdO+nIHh5IIeTB7CvV35VzbOOouu5WbgTTu/wIJfXHgHEanNt7Yhs
y+RaZ2N70B1HDLq9Nb695fu2Cms042WRYt8EUSoZD+eFEn4Z+vggEt7+0mQDFZqX
pGcf3EwEjsZvDroikMvBuxfOjTz2nhDNsfvXppM+yavLDdxhoq5rg9XIGeMgzhfM
gVtEvIg+1SIe/cFOQcg/t8xZlV5f4k0UhKu+QTZiJXPQdNcJEFNqErzkvjgWsVDR
2LA2GABkgBjqfKkaxSrvJ40Bd2swA0h/hY81U796W6wyDGgPMLgF5tTCdN4u++EI
HEU/WXqF7OYdnEZ9dsQ87/ePgj8ooW/MKs8c5ZROArh2XsN3w6RDCgyCUNQntpoL
31E7jq4hWi4iCkGdpCuw0dASWtCZ/KUSHDDtg8l/+xSWOXWUvpMf/b+Tzk+go6Rk
LBd58ipHpFCkEuX9HR1jZXZNmBoy53Zv0dgy6cTkdceDFvkRBBJB/Xq/0FJhKu2K
wTLmglZ4DkkzsT9n3lWqjvWyZIMQK3B4zjdO8NiE+kFoFzSuU7PZqLjNzdc5G2wN
QutxJFF34qSbE1XQtYSyCfUrVXVtxMb4BXx023z/XSDdPZGMBdyNlptPpGOW91hH
kNmXjTxPdFDQVsWLCqbvvgFrpXQwK3R+oMLUxWVTyN7J6j25q7un79bU9Zql6q+H
u4t21qw3N0ZTYMTVx7q58mbbeCkoUvTZXBhycyGlFsMbiknlbmIJxxIJBtmXfVA/
pYh9rB4D7DZMLO5YGzHl8TuDHCI+ZzU54Yce7A8az9Rfpl//5+lGRrAWmNlH1XmA
2OXDJjUgIhgTxGGaxo7PyqNLf7EcRnnDY0ia7pYea4gMYYGjF3vVLzIhf11xr7M8
MrladdWV+jseBhJXbSXzYDzwxMCwyUU7quE8b/P5FlhBAVkT1kGPoqoS02DxCy2b
eo0K1Skm6QqUvE/RxFAj0fVdUaKL9V1w/uNPaT0PVMPPZVHXRxaMRtcsx+p6GmNU
9AAOqOAKq62pULsuBWek08Gf2jS0Y4f9Yjcg4x5DefvLG0SY4FcR7g/xytNpWpG3
grSlYqlC8uy3hb1nWRNJshVHZmfkW532NqdtL6bnz+4tAwoZU1OMt0kmAYJMA7jL
JSIa4p7l/9mRWhYp3iW/HkkXvYV2OBbbQkRplo7F4syIZDzHDW6j8UBcuGirl43q
t5P88Mt6FrFX8Vt2JGaY+JBFqgIqMmU5PtBwWCUZhvFP7ALljhZFU3XxiVKR45Va
fEx4Xv/Jo21jgUAkORLC3OWCbljtsW2Ua/f4dVC/Tynt3C0Iyv21Y3F9zJT31ecJ
BOa0+CQjd14FaA9km1rqjiClA7QVELO6w5oEzS41u4muLMMir2M9HjApQSgLtm19
khhL10GK457wmBk4uTK+8qsTIp54cakWJ/J5rYxpatBl+w1BAMiufp0J49NBJCeO
C1PFREuQUZKeEgp6/WRppZ2RMF0eVFaUNGeQLaHcorhj3u1xcF/hrbvbgRvsmgbp
mnsjlFljGv+7333HdXgtmjxZfneayfoG5wo1ZwOJSkvO9THugpgUdpnE6U0sJOt8
2A/qHbfDq/EFYVgGenWj7HCw4N0dVxui5oxjjHBPobOS0gGFxqWK528zTTiFGu81
9MPuvvDIoi/utbIdFX4u4MMi5Go2VkMMiuPxOm4hSbTXTi6wj3VNF66hU9e9536I
2YYT6dgaOH1PVYCAhYE+CZcAP4VzhJ2CC+uhA/Mi7sDsjJ1vO5jBhR7/KUOkCkjS
05PpXu9+9pD/XwWZ/e9yeLnA0m/VyLFaigRHa4l00B97KxH9pZfCf/kxmcTj5/Je
Xxeigb9zjpuRIlqggL0BD97H7xHidOsY/MHxdTENKHRP5yOS725++oK/DoNX50Tv
K8obV547QlDVlhWEFI/BNA5aZ36qtrPDDPRebTLBe38P9SoFwLIY/g3qowPkkBQH
DkshpP00xG0a93sovjn6Uo20GmvO8/tBltpojbi94ANaNYto6rl4cA2+jPrqxNlo
yaOrEE0Hthk6itJ+moBNN1VNeG1Klj+S+CnlhNJKmOv82Mm+K8hHddPr8m400Zqg
1jGsWQmYxQ2KAt/18z/2YEwC07WnQErTCWZtJIJtrChWTDuTZrg3eJnN2hGlmSdp
1800rm5xZjtQfIJ/xN3XQ8FP/ELR98kTA7jrIPIx5kSCzCT6yGl51Lyt/aXoR+P3
ayXIdxAyFIeWRDubwPiGRqPWd/wtwTZznjKSM1NxPkkd1WutLSnh/zQUb6Potyof
xoI8q1x/UzRgSRViPNCgYmYW2GBq1kD4ug2xkZA1wa2BOWc2mN9/fF0UzKz5Z1+1
67bYf56Y42HZ3AVDcJgkHkMCPs2cjY5f6mi2A12WDIKwl3YWO8vPGC3uS6gI492Q
w3YCjvZjI+E23AtkREWd3G5CzQ36128XzkVuXoKzWKQjAp6o4x9SI7s6T2z2wlyi
IYomkfrruaPIT8/gc08y4mjNYGXWrCY/8DrwX/lMar8nvHPPwmL1lQoUYNz+E9wv
lJunCSGI7fmG/XdH6Dd6oqsWj32tV3TJvaZxL1DecQYF3f9ZyjIV8r9U1RWM8Xw7
GSTKO+tp4h10BxpKyUFOT40A7aStdGideuWO5wubcco8UIjHatT/R7qnu1bmFhve
SJ79gzVuIJGw1pqyo0K9K21zYXdGiKrAgrWGLxLCbsy/S7qOObOLpM8PJV98ts0b
2D+pj0bo62uH/gZk5dakHX63QG/JR/BFsdc2ePN7iD+U26IFnWGCx6piq9XmFb3g
ObeKG8xt7nwA7IKSyan+O9BcJdQvFXkV/YwxLv2hVpNdT9q0RUlqCie2NZNFB7IX
FoNHuO2jhwHY0f8vSrLyN7iROkboFxB+TKM63aQKyfddjX1nK/7lAjqjYvdImpBZ
0SHwVVXi4hBkCHzMax29hyt24YoKyJ1RNwLqQg+6MEeMjnxnOcvtrI+6mfqzyg/w
ipd7erDrMAw0eXht/FijulZNxDk7B9cGiR8afm11grCFz2mXIC4zjEy0YWHfV8IA
bXW2KVY+ZTbTKKfVb7cZyvwM2S8LYxzoZlLJjv7HFWzLLX5GAFfB4EPFTh1VPyVE
tIFcdVa6QEUkG7WNb1ORVVIyvFE/kipBGWjXZV61uYQzVuOK0B4vQ8p6Sd5vXMn3
g1hJbARckEdL2GsA2F5KtekM9lbPJB7zhOoo92+U7UGhw/7h2bi5WXsDGvPkPMEy
nLak+uRr90IfhGw4UrCfvdhgK0oB7ItCRdryzJb9CkhKzHEYw64TG7SNZVPj8zl7
M8hOyMYI2aLC5QrsQP5/zkDpi5q9jt7CzbI3qelvf6SKpB5xE+M2vd/wt0xYNfYV
8LhRjNyTj8SRHSXrsq9vsgnk7xtadzMLcH3rkGXguK1FPJwloVSOab1a0vI1Rc1q
0QSUs0mxowUIEQBFjkAk+iEuAo5+hn4xa5saV1zr/2PY6HZ6X8/u8fnaB6ESqZmy
qe8XqoIEKekOAYkaIa1xV5QBKPs0hWba5e1iLlBvp5l2eCtBAw3safNUg+ZOCYZH
HjBSEVz1Vx6fNdb/4ig/+Ybfgd7ZccPquX4t4OfYgTTjzmOeoPv26hmSExs3VsLg
4m+AW7oEGp0f+rlwknNvAEt7XE7BoMTZgSoLUiYzN+ZO4ysddxJ3AB1j7m5/dQRC
1fOz6gTA2f/ygKn82PLsbWGim5Xzftm32SUjbuiDErQUnl7QqQraIMx5FcNXv05O
7/IvUG5pqKWlo6kSp2I+z3efmgddKfrAHuD1eyn1sKsRbwP/wgEBethGctcd68JZ
FW3TFxeJPfaD0ENmvYqocmH/SAHoisWPcK05bmjQpqFTXxmwxWrBDzpSpk3m55Iz
GPra7A48p+oGgT7LPNemfJtCnGnyiITmRGZyz+xpyfpkkEZ6hFMi/C7u9azPtC2o
O7Act1i8Phc6Z6xZGXvxiNM0/YRiAL9iDyX0YASCDqiYhTQFK9+SvIw/xEXg/U0y
Y5kWmBzrkpuHPDUDN5DT6CxzkT+7y8OBFvdG4JAl8Z2sjuAdTeq4mj0N8hpah4hj
ReVD4hjwSXokR6u4RXI7Vl4+TLhHSeaPbwraTmmPK8VPhd1B+wmCX4pfK8zYkXGx
uoK6U5SfRXvCK612UHvjVKoAs1U4OIBskkeExrEbe5tS+Ld2qdCE20QyyyPDm8Fn
Bs/5EHQZolYnXy6SXs+O9btJch/gSj0WaX5tbD7FxvQSYNtzj0qmRsrBeEEqTPCB
kCIOnvS1j/jTTQKjwSRgRujBbcUsyacwFUwUIpJ2YShE4ORbgPeE8bOttqoqt7Xb
6SNUEIxV+T7Ml49jL15h+eacJd/9FiuIEXEiaAgLiouQQ1CFWNOKjN1Ics780hd5
i2i8tYPg+68pukFnXI9PHj7+L5l2c/wFL7uHA/7u+QdWxT8dcGFx7ZjVNFEjwHJS
ziabXsxRE5Tn1IxZXHxWleMRvjUtRoGweDZAePb2NMGnqXt5A8H0K7al9LTIBlGJ
9GTD71SyZ64pj55gWrPQcSsFji6zlOW2TUl22zcBKOjv0SYsTnQCrXuC5s2UgLmG
O6x9jCZYlcipUQy3DY3myDZP8OAc1CI8QBn1zWG26nOW+ept9XGcKJ0iR7D3lwPk
yAxyX28km1N/WGMaERcO9ShpRj3DF8fEC3l1ixBmR17gkQunNeAUjEcl/iZlFFe7
/zxJY0yTmLlQviLU7cyeh9yG2k/CLMLbp4ScNjV2IF8KgolxFdWWgT8nanIln7V0
hc6+zBWHS9LaoZwxVIx3Gvk9hRJgIWsjHiSv2DU1+4zOA4MzT6oqryyWb7+R2Tnq
kl9W91bK2/Z3fTPFhTLJYFuyu8nVoLAfREd2T5Joyz7eVCIkELGDW9PDVMoK0kCK
dSCFBzpau+ljvizzRetX3nM2AVIjCCd2qBeYEXjwKdI/I9kiE43tCtkOlpFxuciy
dHANwcjReVvO2OYZ4nIJUEjD/MYwOylaLf/x87QDQQWaUHvswOx63eKgwzlzyZlE
edQI7kwUKDN0YBRJFZwhaYgaljpJnjDQ/u01ylr9JHBQjqI3jaJsY315RQCjrQWX
B7qfdDzgmWvXAXMtlK14/GpbSQllU4wDrY+bj1yrMqfzzgIh0X6CnjWnQGHfzvOO
xmAupzHrBoPIEuJ4kbJRki2J8w26I5KXT3k5eUrOs84tXikRdWhDYIhEX0EJnO3N
8L9FRvOQHc39cSSGs67gO7iFTZzn0epY8+bzk2WMzXQv78GJ6l3E0ZS+tlTCyaA/
bNVWbPVfh0WvFpqkbmOZgt70pf37ib+uSgMGybXUFkdk0SuzBcGVpgnE1NA/4BCP
l/a6vfHNri4wZtqvtKsUFP1XkKQEZjSEIIYI0JCV/VrnFefKlaenyh9qW6Uakx8P
1nFNOukJgXGvfPEEmrhLrwVnrlKHMZ4PZDK7dKx8/4E5ZmDKdWHEaPNwT4qgV+DA
tyItrKsdqMWef8EhWw4zdit/fOYMNz1KpcDre4/yoCBf6rPLqDal05v4jeZY48Ls
B/vSX/2PJOYL84G+1yAjb2ZHQOkzEDp5UMOQaC0UrId+rSEvyMWym72wi0W/ntyQ
XSStGQg09AqPq6njmjKPcdAF80M1Z+pLuGihLIA24SgnAeihA27va8lxUwF0BWu7
Yhmy6KTOj/WR9vn3KqtzSCblbsHxq2Ftxyx2j5+wB2sSW7t/0oKEojaLmgqu5OOl
VKtrc6KMEMWek5dwFIBfZ1KdlNbitLsujoiCwhavLlV6IMXLB0Z8Md+QXDcd5RZr
ft7/fXWz8qnGJJx+xJ7u3pEgdgJYg7RwloRQjn4DSh9isEpGsU3r5NLy1bwmHDAZ
vb+M0r/Kuy6QO1fK/jMSK73hJ220S8k3mzbLn5zxSaNnvvnzTPl+TeEBZTaJUhW/
Xxt/dGPeL3UHwmkNlW03KaTcWYXEaYMJwfGp7ewjnMLDB5kPedb7f+GV2b5yAMxn
ncA6r7i+iG/dU+UwIHfJR/oJ4SFgYXGN7k/+zFrfgCfIoBhWEOowtuaojqRhSC+S
Q8UsfD75+rJAMFQp7DsHRRSHc8YHLBdsDu+XH1/xL8RvbpGjUG9jWaJf2lYOSa7G
b4Wb4KPeGCBt9Bn0T9oTuLbb09/SPeNR+I+1N9bUvMOnX811rT9EjfCkrIDQwgmu
W2CyfdiNTbwXE/hOEyF90VHvqYEpAXp6MDpBslUDdsNF8SZzzse/DTjmEC8R5F9Y
I8piuPyMcZCPYSAJix9z+59bMmi7sUkGy3oli6hUaVxo0d5tLHxqIbkioKWNQkRW
X1V6/DRdbOhRPP5hvo88FcrbxEeTRxrmvQvb/GjKzodsoM6QqbY+1MfqqnvjR9X8
ESLS8HFMMvLXMK35buYdx8xilWJdQv8e9oZwpg8iPBQJz7Ypgo8NLxy6LFkyacwt
wdNUJnnaUGgPC+NqUoR0KLkTowV0lKXsTrgoN3+NyCKXuwQbyx4DZRakXU9RV31M
NODpxxdbpxE6i/bhBTpHPlxqEVFFQaNhRvwH//CdlCsaXczu9gqDXuZDMNKnK807
5MKrRlWw2XlPztefm205U/cmkA12LLgikFWtFFjLXsxfJ/zJKJSjy7kbXl5f/23l
yJ9DAA13btEjuXyLiCq9xVOiXVJ7VSYIdCZqlDhlcYQzDHtX77dq4JDUjdoQWk71
jZe1tVMDbYgmf7Seg/Zq6xR3AvKTMOO2ifdg7ttjVsvL01p3L3d1eJi7PIt3dA8k
PJC0kSFF1jRRjygJ8/mIPsbHtNcqHoEPY+AYXnfNJffvL+4M63fD3qQqHUvOg0OO
HYfUAuqWDnKb4B/fVkGvikUll6fSn64vlBRSUfClOGMIRxQLnvzyq3igy6q7MhvE
fjekS8KcWAUrplGmJ1g/vVMXmdi5CvFBA9RROeLsjtNqcung7j98aNFxCuiqrjch
SRGKN+WzllGNACmNvXUGhSwY1RcPXhiv4of+bDegvzwfsIV8o/84qY+xo24NI8Xt
XP3jWP/J43DZ1QlpSvWeSp8IME+5c03bsTq0PtsJq7QJ7Z/8jtlaGEuPiMWm7hNb
HjcuVP+R8vGOu+6OZrEuQLhWPhS8uz+4IK2olQjo6g+p/TIGVWHpbLeus/WcCrjD
LgrFq703fTx7PNLASlXpVVqMOUuMfcwNdGYV+ExTYcIM6SKYSACgujsogydrXLBj
Ya20Rb/071s3L/VIUKKimCuRSidYcyDUQowwQ2t3Qoe5AyAnp5z4njoDVeG8aMY0
R10NryHJ5Kgg1NDOnmj57KPtCWp9pjgDj7cT+t9NmcX3dj+WjSFm+s+ewSRn3+jG
sgRLQpUiBGqXEJ5u4gU/Z4fi+Ja7oSz3ekytdPaq+/LKZOOe/Gmuj/I+EaiwArEj
f4mQ+e6SSq77KCLjDgeuPpR8yqLbrUEdV/sCRrcGDymATZg4+VldwxjCRu9jnrhp
3RWkA0LkaLGDX2BoHBuehW5NhcPFD3u07QD5xqGX7H7xC4l2+rPaFl5aGdF45aov
EhZJONvxa1+/zI2/1ByOY29qT634hVh+RSx77Uk6DNpin85Tdpjnal6B6LQwjVMw
XqwYeG8YGtBj+qkzJ30afPpdYuJmyk/V3mJzua+gbZR9+8kuE3+8aVNjaPPEKuED
MmX9shxW3xHI2MpxhlaHEqsXmEWvrszXRIQPZ3IrYmVXNsp0YrsyDmE8sSfCT6e9
FS9QQ+L1I3FFaJhGGEi4p6fL5TlNF5oP9WFmyDulqmWzCvJywk9j5J0RHtRMuHXb
xvnRvVUcdoWhtNmS/mAuMjHSzzUcWVGVukLMBWk4N95eKKOg8Q5q3R4EpD4lhckQ
J2M5DkBY6FKcIswfKLBIQ6DWVL0C4kk0h2tBppn3yH4KfPm21mP47gzSd/8+lrz0
EDphiGVSw348M8XPP2UROV2wi6XSC5GkXaxP19rLvnDFgzEu1V+DH9hYbqlkEOM4
nvQhwby9wirZtn0bnJbjFijqwMsxRPsXdTeD0DyabMINE0k3rDghFXJXaizIezoA
HZ3QasqfHOWcIjgLW6j+zERxEPWBQhuOhS8nS4EtTfjXOnAu/1D7CxutnxbHPvWu
B3Nt6CU79n8abiTPN68dFzlEOXpByPdptcyrYDoJRGBzeg7WpHrRvrW+N33y8kpt
gULODYgurQmWYQn6cGnVAEHBg0pLWFYvaCxOhoUNYOdTjeYoGEx5DoW94X3M7FZX
6sjqxCj7s+ersc/c5HDaP6VAcau72j11XLyc1mZs56HgnbO9iyZowm7ew9m2sciW
xRNC7/i4LUe1rXMrMQV8bixUsYTngKk9embXXhwZT8dd3egGgWPFY8MsCfyZWiBF
CKBwq0Yq67VDrDkLsSFng2fokIInkIYttR/gi8bW8MKr62et/U8CBn398YC52hLE
KKyDHCAfUzOEmqRoMi6APZp1FO9BLNEBD8ExbuH5XXnLR9EMKVs+r94wZ1fLFvCk
nB+5BGE58ZqbWYUeFPHZwnPrqCc+0q7Xs7Bvp4b68YC2HhQ/xpZmE4cXXgM8dKMt
18Q6hGMcNz7lHmnfFZjK1umzoTKKSG2EMmmluvAtBB9xFCM662CLltXVSpAfnBxl
c8ulAOCm/UzTj18uNxeDMhYj+oDg3SHqAFLWOpKToqAhTRS/iJtTgaxL3BlSOLdN
p0N/iCDShHFt+SGEe2rpPe0Q26vTbnXHGDSypOmJOHXYQn0vIskP5SLemkVvhuNk
pzDaXxNkYDB8Hi6/7P1aozlm/SBZHaeXsdzaZ+0tbQ/xOWcGD9J9SCWfeCjgBTP+
8DQs3gwKfeqVw1W4/dYhmx1KAKA4m3jXYI6cx0NDE/2Wi9RQESGmSuaVopOq137Z
/l/vEjhtTWnIpxpDuyXLPz5pQiuJ3D1+vCgaunmU3TgmdfRSUscEFGyUzqb5kBIF
c1Oiql+BMOtqwbl54FPDDkSSnBg5y+nIIlndoUxWO/FxPP+UFVHFnYmkFf0zSTtr
3ZXnbrf0ijNX/Fc6O6XiOE+Rq//D/sOik3YOsQu4fklETQQSHC63/T+gvlKYcYn0
gmGaEv1h791oCAfIJ5XlOU7iQVKnxBVT0qiVk8au/kUERxv63/AEEvN3paVW2NUX
1QwUVa4vstfnp1DtS+g/Pe8Ze78eltThItIlWMVJ3bgFNKq3qUn7/WeYyyBHrnvb
jvWQGgVkOwUM9ZxOQ6MFrB8U0euiB+Se/GTX0ousVjHtbM36ZLZTx+fr94syb0I0
htsjADg+cOS1u92UNHkbaUuP1RJbJ3N71/BSKKjIESVD88EavugdlT51CjFxunRp
oDJBCEIFipvrBuHmplMqRDQk5JQt7FjLCtayPhE+T2/vYGhhc1YaUAUwEM0Sb1Q7
cRIujlr4WRd6HdgePa8VsA5aAgXF3B/Lu2ye/MXoHXsNCLo+WPiTexIyugPUGYha
6J3Ht8OzPrszft/IX+3Y7LADT2xqchXLlU4di3CxPTF79sgkndC3mUF/wQnonI5i
tdG6vI8320GX92RhNqrXuY/qbssLzByR3Zqwif0vunpPajEgEkoDaulVLKEt3fbJ
mFQdP+gtnXLNd9+NHluJy29n/SlnB7JgRWVs+CpHvenzL1hYPDz3K0y4C1NlxZ6u
A9cqTenczMYwQ+v2Ff41T28MCIHVm2gd7rU8C0M1Z+kqyFf0jsfzwMC1oWiEXKzz
xAnP/XaeA/+swN/t64qBmpTorg2AWldY9SPa+O1FvumPPCQEgxXK6zNMW/ArEGNI
0C68m8CyYSHT8p+9xEuSoOIpR7RGefoNSfaWEgSLxXDGVg0ijJmwdB5540yX3CYU
Of+z+DZGZ5nDyZ5vek7tBttftgOZc0uSblNnmEavPUYkk5M4LNuBR5SXIErtBoO+
Fwbn0P06+OSEUq5ylG2KcdWOz2MMNks9lKn00lxemHQPqKyfy23XX/DnbUo2TWb/
JDaNYHD1SxC2ow9FwJjlu5oF141S+vV/kW+3+5hLjWivki02i1O5UypsvlEP5fV8
BLP++ZOrcpkYm/Q5N1a5/T83KatMx22WMSD9Uounq6vkT34yk38TcamufXemTDGJ
zRZg/ZD9vJCtcvscKoZCZ0QaeGr87Z+7msQ2rzQeVNZAFEuGB5DdfW72BYc1+MDx
pJhAgzMQFLAY74z8zPITaI5D6cF+LQbBxnkoOe8GQ0nY27lDcefhYMipCo4TWhTb
vtUiFM5rmrLo23qiRScr9TojQHm1m9xF3Twq9EAO7kn06+jxRRuK8CwyVDXKqjPG
PD61SMxuX4vduxNifmPqPKxWoeYhG6NGX1ci87TlQRhflaP8G9NSPWz3UZJ677RK
i8+lIHtaFmt+PGjOixuIfJKJApaKszbWqyIgN2Osn80appKkfLvpobXDLK36een9
Z1Rn4i/py6+b6KBdtoxhMbFFJm5nWT9WXvdnXrG2aBygXpM9kSDG1+KfoQ2fyKXZ
n8kuJCtovIhWOKdcSnCFsyq+YJoBNkh9VUOE7+T5TBb5vm+sM/s5+GxyxpZWLc5D
nDOES4hLe5jssdKME9dVtPLnGDx96N3RNgjHgm1yw4rP32Bj3A5CFfZa3t38nrcg
JFstKZSQMzj8+ek71U2aX2a0AKFvbUbE0+g9nOpZT/FksHKSAHRhA4tqManuTuzq
kfHeoFofwe44dkS5QaJWDWgqjSCDTWTGWsyE7HVurG2OjvYgC4wIUP+kIZlFSZRC
iY4rY9XXQEU1hhBWV5eYxiSPprRsrkuP1pWXt4GCHYbJC7WvaXfOYGwf9Nw0TUdR
S3pnQJ/1RCENPOZ6FkmOW6q3GuEECh9GV+1anyrxBrRnbgNqSM+n+Sb6aIUF+c8v
7tRfPoF6woH3p3C+jZBBP+Z2/189wIP9LZWeJv8VLqXyTn1/QGZVgDBgFVncPC/P
r4JRRRXy42WQ1SLn9OVTCHRKc0w4m3OUI6EBAux555G0Rs/jNm100fDxLXz8BddD
W6Rsw2m9GkGVuOWMMC2AUGcz1giF57mXkAQPh0fwPcxMTDrRaLInbuBK9/EApMOq
UVyfqyOR7ZRem9o66k1eIATvF8xnSEPG3Z8hR9dkgWvQQOYC/QwA9Qj9Hqe7xH8O
c1ZDKfPbtbRgo/ALnXKhPoYXMQlI+oQ2q4co/1h6GJCsj0SkWcX50iR4HJOg71Gu
MU/HZwl0YFJNfVCjkJ06nW/7PEtU+zS68C9BVFceUINrFQaGoByND/0vS0FqjFPA
ex6r/zyNzu+WEA3E+kENx2xMZUfa01GyM+WUfVtjdwaVMOxSKXrGzLe/d2d7FDNr
eY4rwX7c9FGX4V8smjGlQEzTepb3V6LYzbIBnSeWaiCJC6xnG8RQVYCuVsaZTCx0
M5sqzq3NyRxofIFh+XGqR/2gf1A7G89alvfSBDoCNKzlHrt/y/N5Ju5BRHjFf9V9
XUd6wGJItKWGwY1qsJ6M6lpnasjMbNGlR9r/XL1xOauivo42fIzu3z/PvjXUTxIW
N3a3mwJnMvnnr6ypXMEHLcWJrKJYPwAkwZRWNx1mNHLwDjqNNTdlJh461lzsNe4X
lPm05Eokwqy2kKiYJJcDDhDFdrt0vAmm5kLjc1F6OD6mIS/tZK/dCOP64uQvII/d
S8t1oxBfpWVIIJfuIs7Mx6Bligwg5pQ8RvVQJWotyEIj/Pvoa2Z2bc7pE9vKGIK6
+arbl61UpCQHiDKc4aEQkvRVibxGszJz+vBu6lV98ILBZHFJDip9bb4eLUd9SC/E
ADqCXBV2/dnBa8KDObZ2uOEMslB1nHT+VBozrByFR1sisiAqfiqI/jVjkBQ8uTvz
037yLi5wVsteGr9ndCxjVnmCWpv0tY0OOy6g2sFWKSgSnT55LSU0zbuEu5ZCVv7C
II74SlSD12tIXrWcGZ9DOuQ7jUwoqq9sR3IHB70aX7oeCIDxA7+oB7QPnRinMXPq
gSU/aFLb0fWLvvnjc/E7cwBc1kbPKLngAIY3KNpcv+VW8ZT5gSCwRLtTQMY3fNhy
Wvr4KNJai25F9AKrxW0QHHoxLcepCo+0SC1UVGy8cuG4LRdFk3ypyf2wHHBn3LC/
YjNIA7YqxmMRapbA1f8wY7bImvkbV/ShzuHU33z5Rv5Y+L8tCB+soJFBzMB24WFl
RuyOEcMNTjzF5ORtFR54SNuLskOcIcVSbLwMP7MnYJsBuEtxwxhigLFyZepPWcT+
MW/hJYzRseKtmr9y8MEYEGmqljyDlXiKC05hCEtJsheJcjN9ucPSphXHdtzccvtV
Dx0qU+ANxhcpa8YI1RCulZky+Jo3ZbNr+ES1nA53C8Fre6cjxdY/84Ljim9o9xNJ
AubF7KQqe9YYaPI9Lcq6JusTHMzcS9p15kWJJEHGvMFH7tAxdTQxUtJNYnEgDpdj
adGpZ26TvoVFC8BS3F4Hldt1KUWU3PBVoQbi41F5WXwZ7tmNNOPInytxxlf3E9Q3
rOAO7RpGtGN26gLFQhMG7aDzrsDjLQ/oAGkYv7vm/AVTYvBFMV6gpkLfdw77eIPk
XgqfKBTIEULtqCjTnD0VQxhwrlvNpF6pykTpTbuvx1DzKe81Dm/LAsGe5BGeC7qn
YcbdxxxRn25tWEf3GBDvqRNxTOTkWk1R60eBiI7ekVrVsLvW44zzw2q6ah0Brn2/
IFCcbFSDMaPmme233vge36SDgY9a4vKXC5wj0OPeEQ5zw16DeK5xGAhdY7rz8rLF
ZEM/HWATRlGZsYD7MiSKl8g9kCoKrA2GERv7r9WE/Kuu1HDYG0BXmgGR1Et9Ss1z
4eYwm/2VUhIs+Esbm9+CrH1Q4JUDhem+2ozXgvbzUomjxLir6hgvU+WpE4kLEdwW
E38zl6/M+dmoW4hCJB44zw8gWMjYHe88te1lf0NjaJCNORTzhUse58eOBRgRniNF
94TcSBgQ6C7zCu8CsEMTZvLIcBent4C9XfSVV2hZmgpnexRJ++v10g0KZ6F3uvls
U54mN+bXycNyxFqscmiRoiH5fKmVo9EVUYDa2yeGWdvn6lFDIEit0mw5dKtYqlpe
MFuMPEWz8dHWVfpl/DjtuAlIQhjvhrFQ5jWvNGKcoIcK9SHLqpxmXFq/p3bFlGZQ
7iRxTw7iEED+mcJvXJtEGFkQUhqgV9TXTWwE/1kz8LO2g9tRg+tU49VF+3I8tzZ/
uuPDmWftLEZcBSiwHoCFf6CZ3P+VGxgdzs4JZZPabjfUcCOmVE90nkfgQ6MXkw0D
c+FRvNIKCcSv0Bjk1TajjygGpac7k4deBEK8v2kd1KcDCZPEi1jXVhH5jbPlvX3m
zelB5QZMxNuWIFBB043rNSdSDZg1LZ1N5fPvFY/+rQWl3dpCQgwOir9Bf6SJqnu9
QHBTTLm2Zhjo5AdEJnWUSLh+vAn8KCbPOQhxvSUZYiEnC9wvBk8RxIsALlHlgS1f
ENtykB2TnmPC7eNSeghO/0BDHaAFkQ3ByqRGACkvppC6EwkO2VK2OD0tXo9o+smL
XFdq02L+rw4qxKckmhNcS9czxIjiOyFUCb/7XDmMGttt5+Pd0mEkiNoRL6y3D7nw
tDFXD1hvlVmQ8UgGP6D/f7M9nghuTx5k8QgLI2j13PpMu1hwKNhPlBv60Ws8LPT5
mAhYFhGnmVm/oM31IgYN6wph5qabCwaE80Sy1ma1OyHTsxWwlzGM7v/RiqMQg42q
X1TxtN5O+gjGSUdurEbH2jj03Hng/9FmYsdY8VPRyhusYTxewDejFjnnrl83cxsu
M7NHNrURVhqZfST1AM6zH80WDZWqqksgPe5o+0Ya243yk6V97zRUx/RVaasoWXvp
IMHerNZvcIWizVLgZjCG8+cMKPJahFcJvokXXmW3pZt++J5a8tS3FxSCP1zMIC3Q
xaa6GAoKrfTz0PBQL/Cy/G+kbVw+5FZVaoqlwidn3xro1I9tVeXkKlIRjxBE0jIA
DWs+5gtLwhw2fn4fBhxsNfUFNW4b85Y7KKB2wMUNM/VGTkTVPAfqL+bi14bC5cy3
3K1v8d7v3Rk+MIyCMmcekqYI/AhHdoIgwAlopnm5R07+zyEbun1O9mzRKZ1rBzhl
sKfdnxc3GOzxyjPodj7mZnQABqYoqI0pzSqef2sPmpbHwMYn6zACzIahK9ykjAf5
WITJ77eV6D+3XsR2BzPbG5eyK1fwrEru6OWN6EHOESW21QxiJ0nDfT4v4W0K5Dcg
JBn53wtJk62h1Q+y0KZwruOnMU0xYJXEcWGoMm2HeUU4rfaFxx4qm8tqJrb+AfZM
1xJ7kOQlV/aBTUSnrHd7tzg9FcO+19MkOzXYQQ4uzr8N4wJ/qp0R5eeDMQBKZlsa
zFsLKMDyQGxXMW9N+2BJ+uGLngzB4HohVpe9KTjnnWvCyZ18oyo62jligpIRCERj
Pzq29vlQ7ulvm+cufAaCnkV4z8f2LeTT/eOziWB+jdJlJINZLn15HLaUlHRQ3duO
4OSx3ZoEft/oBrT341xWYNvDOcfwcnpH0nYX+36uYpTGSK7bsIZVKLLIQy3RSOM6
Xy4+ai8acl6zl3TwYZ9jRmgscBXVWJye1O7aGm/4A/Om4Hgg6ZuK5v5HMBdwx08H
pOZllVNuv6SXOSZiX+A5ALb09dny7/H/+HJVkYLskT9QHmCEAumiMIyf9zvcOREz
fA/gWejTvIqwH9C9X72aKLF1v1Of9A3E6ovMQWoEeKRy61ZlHitnOMAwFNKyYuNN
zx91PE+Lzi7j6hz0Yag04yHgP9vn/IJwi2PBsFyMLnPBR3kh87JfpPRzn10zfyXg
aCHZCmYlsGngA7ZQUe9U58gA9T3K3xUs/PyfgwfN5DV/kA7oiFW+V/9sDmjYRFDO
k3SWemd6/14rW/LximV4OeYJiazgB2T7ah4uiOie0CNmfsuvr6LFRAI6n7v/x2G8
Yfg4DYut2NLPlwC2b06cNX3WSaHBMBKdjUiFkgetuw03awW7lkKxMK1Iald/CWGU
EwWXo/ElW+xATcfCf+xXBZimRlaSF2p/iiA5F8pOXQfYVs5ZeOV9nUSbs6VYo35V
uZEM6k/S0tJ/OcoEpBFyHTq76OF5W40X3RGHlvfW/TVHpYTA+bs+YundlbMDmR9i
gtWACkTITgIfvvifS1JA6E2zalMgcirLwwuRYuzkash2+IoVi6Ni0eQVu2LrZYQG
ewcUjUsJVthkojgk9zeUMm+gzCxXdQSUvgM/20tvNzgerfN466JQEGqoAYbBULOr
jtgnCnx5vOOlNoEPuvBFm+l+XvZPFogIP9rukGMjha/eeKVqmXuVorzeAu13OkIt
jwrOVS9m8+AraioLI4TxWNfca/P0A4z2oriEaPNrTZZqF5cyrDY+HbAqfZBExPvY
a3v3q1SAihE/5/QoNW1RkYmdSpgfdjmRqMs6D19PY96BpefrMp2pAVGH9wLxDxb9
Sm26pvof0JwICSydyYg58rcc2mynKKArqmxe5lF+di5Vw9TlH6wW5M7+jwOUO0Tl
WK1xF9uwgNFAR37ydLX4cKtLRBn2DJ4Alea9SWL1PsOC27g+tfWH2qPO17BdEqf6
H07Hxa3ioLxW40fni+wGaUJW2uPYcBpzHffc3uwXC/umCk9/+YotsmT2eZnasy1f
2VN7BboT+Za+4Vh1neOz5Y5fSfjoM6PxrHZ+k3XYXEZrv66VUcbek0gUZWM3Zmdr
jviIIsiX+BKtWgIqQGGCOQ==
`pragma protect end_protected
