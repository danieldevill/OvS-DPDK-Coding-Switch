-- megafunction wizard: %Cyclone V Hard IP for PCI Express Intel FPGA IP v18.1%
-- GENERATION: XML
-- pcie.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pcie is
	port (
		npor               : in  std_logic                      := '0';             --               npor.npor
		pin_perst          : in  std_logic                      := '0';             --                   .pin_perst
		test_in            : in  std_logic_vector(31 downto 0)  := (others => '0'); --           hip_ctrl.test_in
		simu_mode_pipe     : in  std_logic                      := '0';             --                   .simu_mode_pipe
		pld_clk            : in  std_logic                      := '0';             --            pld_clk.clk
		coreclkout         : out std_logic;                                         --     coreclkout_hip.clk
		refclk             : in  std_logic                      := '0';             --             refclk.clk
		rx_in0             : in  std_logic                      := '0';             --         hip_serial.rx_in0
		rx_in1             : in  std_logic                      := '0';             --                   .rx_in1
		rx_in2             : in  std_logic                      := '0';             --                   .rx_in2
		rx_in3             : in  std_logic                      := '0';             --                   .rx_in3
		tx_out0            : out std_logic;                                         --                   .tx_out0
		tx_out1            : out std_logic;                                         --                   .tx_out1
		tx_out2            : out std_logic;                                         --                   .tx_out2
		tx_out3            : out std_logic;                                         --                   .tx_out3
		rx_st_valid        : out std_logic;                                         --              rx_st.valid
		rx_st_sop          : out std_logic;                                         --                   .startofpacket
		rx_st_eop          : out std_logic;                                         --                   .endofpacket
		rx_st_ready        : in  std_logic                      := '0';             --                   .ready
		rx_st_err          : out std_logic;                                         --                   .error
		rx_st_data         : out std_logic_vector(63 downto 0);                     --                   .data
		rx_st_bar          : out std_logic_vector(7 downto 0);                      --          rx_bar_be.rx_st_bar
		rx_st_mask         : in  std_logic                      := '0';             --                   .rx_st_mask
		tx_st_valid        : in  std_logic                      := '0';             --              tx_st.valid
		tx_st_sop          : in  std_logic                      := '0';             --                   .startofpacket
		tx_st_eop          : in  std_logic                      := '0';             --                   .endofpacket
		tx_st_ready        : out std_logic;                                         --                   .ready
		tx_st_err          : in  std_logic                      := '0';             --                   .error
		tx_st_data         : in  std_logic_vector(63 downto 0)  := (others => '0'); --                   .data
		tx_fifo_empty      : out std_logic;                                         --            tx_fifo.fifo_empty
		tx_cred_datafccp   : out std_logic_vector(11 downto 0);                     --            tx_cred.tx_cred_datafccp
		tx_cred_datafcnp   : out std_logic_vector(11 downto 0);                     --                   .tx_cred_datafcnp
		tx_cred_datafcp    : out std_logic_vector(11 downto 0);                     --                   .tx_cred_datafcp
		tx_cred_fchipcons  : out std_logic_vector(5 downto 0);                      --                   .tx_cred_fchipcons
		tx_cred_fcinfinite : out std_logic_vector(5 downto 0);                      --                   .tx_cred_fcinfinite
		tx_cred_hdrfccp    : out std_logic_vector(7 downto 0);                      --                   .tx_cred_hdrfccp
		tx_cred_hdrfcnp    : out std_logic_vector(7 downto 0);                      --                   .tx_cred_hdrfcnp
		tx_cred_hdrfcp     : out std_logic_vector(7 downto 0);                      --                   .tx_cred_hdrfcp
		sim_pipe_pclk_in   : in  std_logic                      := '0';             --           hip_pipe.sim_pipe_pclk_in
		sim_pipe_rate      : out std_logic_vector(1 downto 0);                      --                   .sim_pipe_rate
		sim_ltssmstate     : out std_logic_vector(4 downto 0);                      --                   .sim_ltssmstate
		eidleinfersel0     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel0
		eidleinfersel1     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel1
		eidleinfersel2     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel2
		eidleinfersel3     : out std_logic_vector(2 downto 0);                      --                   .eidleinfersel3
		powerdown0         : out std_logic_vector(1 downto 0);                      --                   .powerdown0
		powerdown1         : out std_logic_vector(1 downto 0);                      --                   .powerdown1
		powerdown2         : out std_logic_vector(1 downto 0);                      --                   .powerdown2
		powerdown3         : out std_logic_vector(1 downto 0);                      --                   .powerdown3
		rxpolarity0        : out std_logic;                                         --                   .rxpolarity0
		rxpolarity1        : out std_logic;                                         --                   .rxpolarity1
		rxpolarity2        : out std_logic;                                         --                   .rxpolarity2
		rxpolarity3        : out std_logic;                                         --                   .rxpolarity3
		txcompl0           : out std_logic;                                         --                   .txcompl0
		txcompl1           : out std_logic;                                         --                   .txcompl1
		txcompl2           : out std_logic;                                         --                   .txcompl2
		txcompl3           : out std_logic;                                         --                   .txcompl3
		txdata0            : out std_logic_vector(7 downto 0);                      --                   .txdata0
		txdata1            : out std_logic_vector(7 downto 0);                      --                   .txdata1
		txdata2            : out std_logic_vector(7 downto 0);                      --                   .txdata2
		txdata3            : out std_logic_vector(7 downto 0);                      --                   .txdata3
		txdatak0           : out std_logic;                                         --                   .txdatak0
		txdatak1           : out std_logic;                                         --                   .txdatak1
		txdatak2           : out std_logic;                                         --                   .txdatak2
		txdatak3           : out std_logic;                                         --                   .txdatak3
		txdetectrx0        : out std_logic;                                         --                   .txdetectrx0
		txdetectrx1        : out std_logic;                                         --                   .txdetectrx1
		txdetectrx2        : out std_logic;                                         --                   .txdetectrx2
		txdetectrx3        : out std_logic;                                         --                   .txdetectrx3
		txelecidle0        : out std_logic;                                         --                   .txelecidle0
		txelecidle1        : out std_logic;                                         --                   .txelecidle1
		txelecidle2        : out std_logic;                                         --                   .txelecidle2
		txelecidle3        : out std_logic;                                         --                   .txelecidle3
		txswing0           : out std_logic;                                         --                   .txswing0
		txswing1           : out std_logic;                                         --                   .txswing1
		txswing2           : out std_logic;                                         --                   .txswing2
		txswing3           : out std_logic;                                         --                   .txswing3
		txmargin0          : out std_logic_vector(2 downto 0);                      --                   .txmargin0
		txmargin1          : out std_logic_vector(2 downto 0);                      --                   .txmargin1
		txmargin2          : out std_logic_vector(2 downto 0);                      --                   .txmargin2
		txmargin3          : out std_logic_vector(2 downto 0);                      --                   .txmargin3
		txdeemph0          : out std_logic;                                         --                   .txdeemph0
		txdeemph1          : out std_logic;                                         --                   .txdeemph1
		txdeemph2          : out std_logic;                                         --                   .txdeemph2
		txdeemph3          : out std_logic;                                         --                   .txdeemph3
		phystatus0         : in  std_logic                      := '0';             --                   .phystatus0
		phystatus1         : in  std_logic                      := '0';             --                   .phystatus1
		phystatus2         : in  std_logic                      := '0';             --                   .phystatus2
		phystatus3         : in  std_logic                      := '0';             --                   .phystatus3
		rxdata0            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata0
		rxdata1            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata1
		rxdata2            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata2
		rxdata3            : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .rxdata3
		rxdatak0           : in  std_logic                      := '0';             --                   .rxdatak0
		rxdatak1           : in  std_logic                      := '0';             --                   .rxdatak1
		rxdatak2           : in  std_logic                      := '0';             --                   .rxdatak2
		rxdatak3           : in  std_logic                      := '0';             --                   .rxdatak3
		rxelecidle0        : in  std_logic                      := '0';             --                   .rxelecidle0
		rxelecidle1        : in  std_logic                      := '0';             --                   .rxelecidle1
		rxelecidle2        : in  std_logic                      := '0';             --                   .rxelecidle2
		rxelecidle3        : in  std_logic                      := '0';             --                   .rxelecidle3
		rxstatus0          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus0
		rxstatus1          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus1
		rxstatus2          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus2
		rxstatus3          : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .rxstatus3
		rxvalid0           : in  std_logic                      := '0';             --                   .rxvalid0
		rxvalid1           : in  std_logic                      := '0';             --                   .rxvalid1
		rxvalid2           : in  std_logic                      := '0';             --                   .rxvalid2
		rxvalid3           : in  std_logic                      := '0';             --                   .rxvalid3
		reset_status       : out std_logic;                                         --            hip_rst.reset_status
		serdes_pll_locked  : out std_logic;                                         --                   .serdes_pll_locked
		pld_clk_inuse      : out std_logic;                                         --                   .pld_clk_inuse
		pld_core_ready     : in  std_logic                      := '0';             --                   .pld_core_ready
		testin_zero        : out std_logic;                                         --                   .testin_zero
		lmi_addr           : in  std_logic_vector(11 downto 0)  := (others => '0'); --                lmi.lmi_addr
		lmi_din            : in  std_logic_vector(31 downto 0)  := (others => '0'); --                   .lmi_din
		lmi_rden           : in  std_logic                      := '0';             --                   .lmi_rden
		lmi_wren           : in  std_logic                      := '0';             --                   .lmi_wren
		lmi_ack            : out std_logic;                                         --                   .lmi_ack
		lmi_dout           : out std_logic_vector(31 downto 0);                     --                   .lmi_dout
		pm_auxpwr          : in  std_logic                      := '0';             --         power_mngt.pm_auxpwr
		pm_data            : in  std_logic_vector(9 downto 0)   := (others => '0'); --                   .pm_data
		pme_to_cr          : in  std_logic                      := '0';             --                   .pme_to_cr
		pm_event           : in  std_logic                      := '0';             --                   .pm_event
		pme_to_sr          : out std_logic;                                         --                   .pme_to_sr
		reconfig_to_xcvr   : in  std_logic_vector(349 downto 0) := (others => '0'); --   reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr : out std_logic_vector(229 downto 0);                    -- reconfig_from_xcvr.reconfig_from_xcvr
		app_msi_num        : in  std_logic_vector(4 downto 0)   := (others => '0'); --            int_msi.app_msi_num
		app_msi_req        : in  std_logic                      := '0';             --                   .app_msi_req
		app_msi_tc         : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .app_msi_tc
		app_msi_ack        : out std_logic;                                         --                   .app_msi_ack
		app_int_sts_vec    : in  std_logic                      := '0';             --                   .app_int_sts
		tl_hpg_ctrl_er     : in  std_logic_vector(4 downto 0)   := (others => '0'); --          config_tl.hpg_ctrler
		tl_cfg_ctl         : out std_logic_vector(31 downto 0);                     --                   .tl_cfg_ctl
		cpl_err            : in  std_logic_vector(6 downto 0)   := (others => '0'); --                   .cpl_err
		tl_cfg_add         : out std_logic_vector(3 downto 0);                      --                   .tl_cfg_add
		tl_cfg_ctl_wr      : out std_logic;                                         --                   .tl_cfg_ctl_wr
		tl_cfg_sts_wr      : out std_logic;                                         --                   .tl_cfg_sts_wr
		tl_cfg_sts         : out std_logic_vector(52 downto 0);                     --                   .tl_cfg_sts
		cpl_pending        : in  std_logic_vector(0 downto 0)   := (others => '0'); --                   .cpl_pending
		derr_cor_ext_rcv0  : out std_logic;                                         --         hip_status.derr_cor_ext_rcv
		derr_cor_ext_rpl   : out std_logic;                                         --                   .derr_cor_ext_rpl
		derr_rpl           : out std_logic;                                         --                   .derr_rpl
		dlup_exit          : out std_logic;                                         --                   .dlup_exit
		dl_ltssm           : out std_logic_vector(4 downto 0);                      --                   .ltssmstate
		ev128ns            : out std_logic;                                         --                   .ev128ns
		ev1us              : out std_logic;                                         --                   .ev1us
		hotrst_exit        : out std_logic;                                         --                   .hotrst_exit
		int_status         : out std_logic_vector(3 downto 0);                      --                   .int_status
		l2_exit            : out std_logic;                                         --                   .l2_exit
		lane_act           : out std_logic_vector(3 downto 0);                      --                   .lane_act
		ko_cpl_spc_header  : out std_logic_vector(7 downto 0);                      --                   .ko_cpl_spc_header
		ko_cpl_spc_data    : out std_logic_vector(11 downto 0);                     --                   .ko_cpl_spc_data
		dl_current_speed   : out std_logic_vector(1 downto 0)                       --   hip_currentspeed.currentspeed
	);
end entity pcie;

architecture rtl of pcie is
	component altpcie_cv_hip_ast_hwtcl is
		generic (
			ACDS_VERSION_HWTCL                        : string  := "18.1";
			lane_mask_hwtcl                           : string  := "x4";
			gen12_lane_rate_mode_hwtcl                : string  := "Gen1 (2.5 Gbps)";
			pcie_spec_version_hwtcl                   : string  := "2.1";
			ast_width_hwtcl                           : string  := "Avalon-ST 64-bit";
			pll_refclk_freq_hwtcl                     : string  := "100 MHz";
			set_pld_clk_x1_625MHz_hwtcl               : integer := 0;
			in_cvp_mode_hwtcl                         : integer := 0;
			hip_reconfig_hwtcl                        : integer := 0;
			num_of_func_hwtcl                         : integer := 1;
			use_crc_forwarding_hwtcl                  : integer := 0;
			port_link_number_hwtcl                    : integer := 1;
			slotclkcfg_hwtcl                          : integer := 1;
			enable_slot_register_hwtcl                : integer := 0;
			vsec_id_hwtcl                             : integer := 4466;
			vsec_rev_hwtcl                            : integer := 0;
			user_id_hwtcl                             : integer := 0;
			porttype_func0_hwtcl                      : string  := "Native endpoint";
			bar0_size_mask_0_hwtcl                    : integer := 28;
			bar0_io_space_0_hwtcl                     : string  := "Disabled";
			bar0_64bit_mem_space_0_hwtcl              : string  := "Enabled";
			bar0_prefetchable_0_hwtcl                 : string  := "Enabled";
			bar1_size_mask_0_hwtcl                    : integer := 0;
			bar1_io_space_0_hwtcl                     : string  := "Disabled";
			bar1_prefetchable_0_hwtcl                 : string  := "Disabled";
			bar2_size_mask_0_hwtcl                    : integer := 0;
			bar2_io_space_0_hwtcl                     : string  := "Disabled";
			bar2_64bit_mem_space_0_hwtcl              : string  := "Disabled";
			bar2_prefetchable_0_hwtcl                 : string  := "Disabled";
			bar3_size_mask_0_hwtcl                    : integer := 0;
			bar3_io_space_0_hwtcl                     : string  := "Disabled";
			bar3_prefetchable_0_hwtcl                 : string  := "Disabled";
			bar4_size_mask_0_hwtcl                    : integer := 0;
			bar4_io_space_0_hwtcl                     : string  := "Disabled";
			bar4_64bit_mem_space_0_hwtcl              : string  := "Disabled";
			bar4_prefetchable_0_hwtcl                 : string  := "Disabled";
			bar5_size_mask_0_hwtcl                    : integer := 0;
			bar5_io_space_0_hwtcl                     : string  := "Disabled";
			bar5_prefetchable_0_hwtcl                 : string  := "Disabled";
			expansion_base_address_register_0_hwtcl   : integer := 0;
			io_window_addr_width_hwtcl                : integer := 0;
			prefetchable_mem_window_addr_width_hwtcl  : integer := 0;
			vendor_id_0_hwtcl                         : integer := 0;
			device_id_0_hwtcl                         : integer := 1;
			revision_id_0_hwtcl                       : integer := 1;
			class_code_0_hwtcl                        : integer := 0;
			subsystem_vendor_id_0_hwtcl               : integer := 0;
			subsystem_device_id_0_hwtcl               : integer := 0;
			max_payload_size_0_hwtcl                  : integer := 128;
			extend_tag_field_0_hwtcl                  : string  := "32";
			completion_timeout_0_hwtcl                : string  := "ABCD";
			enable_completion_timeout_disable_0_hwtcl : integer := 1;
			flr_capability_0_hwtcl                    : integer := 0;
			use_aer_0_hwtcl                           : integer := 0;
			ecrc_check_capable_0_hwtcl                : integer := 0;
			ecrc_gen_capable_0_hwtcl                  : integer := 0;
			dll_active_report_support_0_hwtcl         : integer := 0;
			surprise_down_error_support_0_hwtcl       : integer := 0;
			msi_multi_message_capable_0_hwtcl         : string  := "4";
			msi_64bit_addressing_capable_0_hwtcl      : string  := "true";
			msi_masking_capable_0_hwtcl               : string  := "false";
			msi_support_0_hwtcl                       : string  := "true";
			enable_function_msix_support_0_hwtcl      : integer := 0;
			msix_table_size_0_hwtcl                   : integer := 0;
			msix_table_offset_0_hwtcl                 : string  := "0";
			msix_table_bir_0_hwtcl                    : integer := 0;
			msix_pba_offset_0_hwtcl                   : string  := "0";
			msix_pba_bir_0_hwtcl                      : integer := 0;
			interrupt_pin_0_hwtcl                     : string  := "inta";
			slot_power_scale_0_hwtcl                  : integer := 0;
			slot_power_limit_0_hwtcl                  : integer := 0;
			slot_number_0_hwtcl                       : integer := 0;
			rx_ei_l0s_0_hwtcl                         : integer := 0;
			endpoint_l0_latency_0_hwtcl               : integer := 0;
			endpoint_l1_latency_0_hwtcl               : integer := 0;
			reconfig_to_xcvr_width                    : integer := 10;
			hip_hard_reset_hwtcl                      : integer := 0;
			reconfig_from_xcvr_width                  : integer := 10;
			single_rx_detect_hwtcl                    : integer := 0;
			enable_l0s_aspm_hwtcl                     : string  := "false";
			aspm_optionality_hwtcl                    : string  := "false";
			enable_adapter_half_rate_mode_hwtcl       : string  := "false";
			millisecond_cycle_count_hwtcl             : integer := 248500;
			credit_buffer_allocation_aux_hwtcl        : string  := "balanced";
			vc0_rx_flow_ctrl_posted_header_hwtcl      : integer := 50;
			vc0_rx_flow_ctrl_posted_data_hwtcl        : integer := 360;
			vc0_rx_flow_ctrl_nonposted_header_hwtcl   : integer := 54;
			vc0_rx_flow_ctrl_nonposted_data_hwtcl     : integer := 0;
			vc0_rx_flow_ctrl_compl_header_hwtcl       : integer := 112;
			vc0_rx_flow_ctrl_compl_data_hwtcl         : integer := 448;
			cpl_spc_header_hwtcl                      : integer := 112;
			cpl_spc_data_hwtcl                        : integer := 448;
			port_width_data_hwtcl                     : integer := 64;
			bypass_clk_switch_hwtcl                   : string  := "disable";
			cvp_rate_sel_hwtcl                        : string  := "full_rate";
			cvp_data_compressed_hwtcl                 : string  := "false";
			cvp_data_encrypted_hwtcl                  : string  := "false";
			cvp_mode_reset_hwtcl                      : string  := "false";
			cvp_clk_reset_hwtcl                       : string  := "false";
			core_clk_sel_hwtcl                        : string  := "pld_clk";
			enable_rx_buffer_checking_hwtcl           : string  := "false";
			disable_link_x2_support_hwtcl             : string  := "false";
			device_number_hwtcl                       : integer := 0;
			pipex1_debug_sel_hwtcl                    : string  := "disable";
			pclk_out_sel_hwtcl                        : string  := "pclk";
			no_soft_reset_hwtcl                       : string  := "false";
			d1_support_hwtcl                          : string  := "false";
			d2_support_hwtcl                          : string  := "false";
			d0_pme_hwtcl                              : string  := "false";
			d1_pme_hwtcl                              : string  := "false";
			d2_pme_hwtcl                              : string  := "false";
			d3_hot_pme_hwtcl                          : string  := "false";
			d3_cold_pme_hwtcl                         : string  := "false";
			low_priority_vc_hwtcl                     : string  := "single_vc";
			enable_l1_aspm_hwtcl                      : string  := "false";
			l1_exit_latency_sameclock_hwtcl           : integer := 0;
			l1_exit_latency_diffclock_hwtcl           : integer := 0;
			hot_plug_support_hwtcl                    : integer := 0;
			no_command_completed_hwtcl                : string  := "false";
			eie_before_nfts_count_hwtcl               : integer := 4;
			gen2_diffclock_nfts_count_hwtcl           : integer := 255;
			gen2_sameclock_nfts_count_hwtcl           : integer := 255;
			deemphasis_enable_hwtcl                   : string  := "false";
			l0_exit_latency_sameclock_hwtcl           : integer := 6;
			l0_exit_latency_diffclock_hwtcl           : integer := 6;
			vc0_clk_enable_hwtcl                      : string  := "true";
			register_pipe_signals_hwtcl               : string  := "true";
			tx_cdc_almost_empty_hwtcl                 : integer := 5;
			rx_l0s_count_idl_hwtcl                    : integer := 0;
			cdc_dummy_insert_limit_hwtcl              : integer := 11;
			ei_delay_powerdown_count_hwtcl            : integer := 10;
			skp_os_schedule_count_hwtcl               : integer := 0;
			fc_init_timer_hwtcl                       : integer := 1024;
			l01_entry_latency_hwtcl                   : integer := 31;
			flow_control_update_count_hwtcl           : integer := 30;
			flow_control_timeout_count_hwtcl          : integer := 200;
			retry_buffer_last_active_address_hwtcl    : integer := 255;
			reserved_debug_hwtcl                      : integer := 0;
			use_tl_cfg_sync_hwtcl                     : integer := 1;
			diffclock_nfts_count_hwtcl                : integer := 255;
			sameclock_nfts_count_hwtcl                : integer := 255;
			l2_async_logic_hwtcl                      : string  := "disable";
			rx_cdc_almost_full_hwtcl                  : integer := 12;
			tx_cdc_almost_full_hwtcl                  : integer := 11;
			indicator_hwtcl                           : integer := 0;
			maximum_current_0_hwtcl                   : integer := 0;
			disable_snoop_packet_0_hwtcl              : string  := "false";
			bridge_port_vga_enable_0_hwtcl            : string  := "false";
			bridge_port_ssid_support_0_hwtcl          : string  := "false";
			ssvid_0_hwtcl                             : integer := 0;
			ssid_0_hwtcl                              : integer := 0;
			porttype_func1_hwtcl                      : string  := "Native endpoint";
			bar0_size_mask_1_hwtcl                    : integer := 28;
			bar0_io_space_1_hwtcl                     : string  := "Disabled";
			bar0_64bit_mem_space_1_hwtcl              : string  := "Enabled";
			bar0_prefetchable_1_hwtcl                 : string  := "Enabled";
			bar1_size_mask_1_hwtcl                    : integer := 0;
			bar1_io_space_1_hwtcl                     : string  := "Disabled";
			bar1_prefetchable_1_hwtcl                 : string  := "Disabled";
			bar2_size_mask_1_hwtcl                    : integer := 0;
			bar2_io_space_1_hwtcl                     : string  := "Disabled";
			bar2_64bit_mem_space_1_hwtcl              : string  := "Disabled";
			bar2_prefetchable_1_hwtcl                 : string  := "Disabled";
			bar3_size_mask_1_hwtcl                    : integer := 0;
			bar3_io_space_1_hwtcl                     : string  := "Disabled";
			bar3_prefetchable_1_hwtcl                 : string  := "Disabled";
			bar4_size_mask_1_hwtcl                    : integer := 0;
			bar4_io_space_1_hwtcl                     : string  := "Disabled";
			bar4_64bit_mem_space_1_hwtcl              : string  := "Disabled";
			bar4_prefetchable_1_hwtcl                 : string  := "Disabled";
			bar5_size_mask_1_hwtcl                    : integer := 0;
			bar5_io_space_1_hwtcl                     : string  := "Disabled";
			bar5_prefetchable_1_hwtcl                 : string  := "Disabled";
			expansion_base_address_register_1_hwtcl   : integer := 0;
			vendor_id_1_hwtcl                         : integer := 0;
			device_id_1_hwtcl                         : integer := 1;
			revision_id_1_hwtcl                       : integer := 1;
			class_code_1_hwtcl                        : integer := 0;
			subsystem_vendor_id_1_hwtcl               : integer := 0;
			subsystem_device_id_1_hwtcl               : integer := 0;
			max_payload_size_1_hwtcl                  : integer := 128;
			extend_tag_field_1_hwtcl                  : string  := "32";
			completion_timeout_1_hwtcl                : string  := "ABCD";
			enable_completion_timeout_disable_1_hwtcl : integer := 1;
			flr_capability_1_hwtcl                    : integer := 0;
			use_aer_1_hwtcl                           : integer := 0;
			ecrc_check_capable_1_hwtcl                : integer := 0;
			ecrc_gen_capable_1_hwtcl                  : integer := 0;
			dll_active_report_support_1_hwtcl         : integer := 0;
			surprise_down_error_support_1_hwtcl       : integer := 0;
			msi_multi_message_capable_1_hwtcl         : string  := "4";
			msi_64bit_addressing_capable_1_hwtcl      : string  := "true";
			msi_masking_capable_1_hwtcl               : string  := "false";
			msi_support_1_hwtcl                       : string  := "true";
			enable_function_msix_support_1_hwtcl      : integer := 0;
			msix_table_size_1_hwtcl                   : integer := 0;
			msix_table_offset_1_hwtcl                 : string  := "0";
			msix_table_bir_1_hwtcl                    : integer := 0;
			msix_pba_offset_1_hwtcl                   : string  := "0";
			msix_pba_bir_1_hwtcl                      : integer := 0;
			interrupt_pin_1_hwtcl                     : string  := "inta";
			slot_power_scale_1_hwtcl                  : integer := 0;
			slot_power_limit_1_hwtcl                  : integer := 0;
			slot_number_1_hwtcl                       : integer := 0;
			rx_ei_l0s_1_hwtcl                         : integer := 0;
			endpoint_l0_latency_1_hwtcl               : integer := 0;
			endpoint_l1_latency_1_hwtcl               : integer := 0;
			maximum_current_1_hwtcl                   : integer := 0;
			disable_snoop_packet_1_hwtcl              : string  := "false";
			bridge_port_vga_enable_1_hwtcl            : string  := "false";
			bridge_port_ssid_support_1_hwtcl          : string  := "false";
			ssvid_1_hwtcl                             : integer := 0;
			ssid_1_hwtcl                              : integer := 0;
			porttype_func2_hwtcl                      : string  := "Native endpoint";
			bar0_size_mask_2_hwtcl                    : integer := 28;
			bar0_io_space_2_hwtcl                     : string  := "Disabled";
			bar0_64bit_mem_space_2_hwtcl              : string  := "Enabled";
			bar0_prefetchable_2_hwtcl                 : string  := "Enabled";
			bar1_size_mask_2_hwtcl                    : integer := 0;
			bar1_io_space_2_hwtcl                     : string  := "Disabled";
			bar1_prefetchable_2_hwtcl                 : string  := "Disabled";
			bar2_size_mask_2_hwtcl                    : integer := 0;
			bar2_io_space_2_hwtcl                     : string  := "Disabled";
			bar2_64bit_mem_space_2_hwtcl              : string  := "Disabled";
			bar2_prefetchable_2_hwtcl                 : string  := "Disabled";
			bar3_size_mask_2_hwtcl                    : integer := 0;
			bar3_io_space_2_hwtcl                     : string  := "Disabled";
			bar3_prefetchable_2_hwtcl                 : string  := "Disabled";
			bar4_size_mask_2_hwtcl                    : integer := 0;
			bar4_io_space_2_hwtcl                     : string  := "Disabled";
			bar4_64bit_mem_space_2_hwtcl              : string  := "Disabled";
			bar4_prefetchable_2_hwtcl                 : string  := "Disabled";
			bar5_size_mask_2_hwtcl                    : integer := 0;
			bar5_io_space_2_hwtcl                     : string  := "Disabled";
			bar5_prefetchable_2_hwtcl                 : string  := "Disabled";
			expansion_base_address_register_2_hwtcl   : integer := 0;
			vendor_id_2_hwtcl                         : integer := 0;
			device_id_2_hwtcl                         : integer := 1;
			revision_id_2_hwtcl                       : integer := 1;
			class_code_2_hwtcl                        : integer := 0;
			subsystem_vendor_id_2_hwtcl               : integer := 0;
			subsystem_device_id_2_hwtcl               : integer := 0;
			max_payload_size_2_hwtcl                  : integer := 128;
			extend_tag_field_2_hwtcl                  : string  := "32";
			completion_timeout_2_hwtcl                : string  := "ABCD";
			enable_completion_timeout_disable_2_hwtcl : integer := 1;
			flr_capability_2_hwtcl                    : integer := 0;
			use_aer_2_hwtcl                           : integer := 0;
			ecrc_check_capable_2_hwtcl                : integer := 0;
			ecrc_gen_capable_2_hwtcl                  : integer := 0;
			dll_active_report_support_2_hwtcl         : integer := 0;
			surprise_down_error_support_2_hwtcl       : integer := 0;
			msi_multi_message_capable_2_hwtcl         : string  := "4";
			msi_64bit_addressing_capable_2_hwtcl      : string  := "true";
			msi_masking_capable_2_hwtcl               : string  := "false";
			msi_support_2_hwtcl                       : string  := "true";
			enable_function_msix_support_2_hwtcl      : integer := 0;
			msix_table_size_2_hwtcl                   : integer := 0;
			msix_table_offset_2_hwtcl                 : string  := "0";
			msix_table_bir_2_hwtcl                    : integer := 0;
			msix_pba_offset_2_hwtcl                   : string  := "0";
			msix_pba_bir_2_hwtcl                      : integer := 0;
			interrupt_pin_2_hwtcl                     : string  := "inta";
			slot_power_scale_2_hwtcl                  : integer := 0;
			slot_power_limit_2_hwtcl                  : integer := 0;
			slot_number_2_hwtcl                       : integer := 0;
			rx_ei_l0s_2_hwtcl                         : integer := 0;
			endpoint_l0_latency_2_hwtcl               : integer := 0;
			endpoint_l1_latency_2_hwtcl               : integer := 0;
			maximum_current_2_hwtcl                   : integer := 0;
			disable_snoop_packet_2_hwtcl              : string  := "false";
			bridge_port_vga_enable_2_hwtcl            : string  := "false";
			bridge_port_ssid_support_2_hwtcl          : string  := "false";
			ssvid_2_hwtcl                             : integer := 0;
			ssid_2_hwtcl                              : integer := 0;
			porttype_func3_hwtcl                      : string  := "Native endpoint";
			bar0_size_mask_3_hwtcl                    : integer := 28;
			bar0_io_space_3_hwtcl                     : string  := "Disabled";
			bar0_64bit_mem_space_3_hwtcl              : string  := "Enabled";
			bar0_prefetchable_3_hwtcl                 : string  := "Enabled";
			bar1_size_mask_3_hwtcl                    : integer := 0;
			bar1_io_space_3_hwtcl                     : string  := "Disabled";
			bar1_prefetchable_3_hwtcl                 : string  := "Disabled";
			bar2_size_mask_3_hwtcl                    : integer := 0;
			bar2_io_space_3_hwtcl                     : string  := "Disabled";
			bar2_64bit_mem_space_3_hwtcl              : string  := "Disabled";
			bar2_prefetchable_3_hwtcl                 : string  := "Disabled";
			bar3_size_mask_3_hwtcl                    : integer := 0;
			bar3_io_space_3_hwtcl                     : string  := "Disabled";
			bar3_prefetchable_3_hwtcl                 : string  := "Disabled";
			bar4_size_mask_3_hwtcl                    : integer := 0;
			bar4_io_space_3_hwtcl                     : string  := "Disabled";
			bar4_64bit_mem_space_3_hwtcl              : string  := "Disabled";
			bar4_prefetchable_3_hwtcl                 : string  := "Disabled";
			bar5_size_mask_3_hwtcl                    : integer := 0;
			bar5_io_space_3_hwtcl                     : string  := "Disabled";
			bar5_prefetchable_3_hwtcl                 : string  := "Disabled";
			expansion_base_address_register_3_hwtcl   : integer := 0;
			vendor_id_3_hwtcl                         : integer := 0;
			device_id_3_hwtcl                         : integer := 1;
			revision_id_3_hwtcl                       : integer := 1;
			class_code_3_hwtcl                        : integer := 0;
			subsystem_vendor_id_3_hwtcl               : integer := 0;
			subsystem_device_id_3_hwtcl               : integer := 0;
			max_payload_size_3_hwtcl                  : integer := 128;
			extend_tag_field_3_hwtcl                  : string  := "32";
			completion_timeout_3_hwtcl                : string  := "ABCD";
			enable_completion_timeout_disable_3_hwtcl : integer := 1;
			flr_capability_3_hwtcl                    : integer := 0;
			use_aer_3_hwtcl                           : integer := 0;
			ecrc_check_capable_3_hwtcl                : integer := 0;
			ecrc_gen_capable_3_hwtcl                  : integer := 0;
			dll_active_report_support_3_hwtcl         : integer := 0;
			surprise_down_error_support_3_hwtcl       : integer := 0;
			msi_multi_message_capable_3_hwtcl         : string  := "4";
			msi_64bit_addressing_capable_3_hwtcl      : string  := "true";
			msi_masking_capable_3_hwtcl               : string  := "false";
			msi_support_3_hwtcl                       : string  := "true";
			enable_function_msix_support_3_hwtcl      : integer := 0;
			msix_table_size_3_hwtcl                   : integer := 0;
			msix_table_offset_3_hwtcl                 : string  := "0";
			msix_table_bir_3_hwtcl                    : integer := 0;
			msix_pba_offset_3_hwtcl                   : string  := "0";
			msix_pba_bir_3_hwtcl                      : integer := 0;
			interrupt_pin_3_hwtcl                     : string  := "inta";
			slot_power_scale_3_hwtcl                  : integer := 0;
			slot_power_limit_3_hwtcl                  : integer := 0;
			slot_number_3_hwtcl                       : integer := 0;
			rx_ei_l0s_3_hwtcl                         : integer := 0;
			endpoint_l0_latency_3_hwtcl               : integer := 0;
			endpoint_l1_latency_3_hwtcl               : integer := 0;
			maximum_current_3_hwtcl                   : integer := 0;
			disable_snoop_packet_3_hwtcl              : string  := "false";
			bridge_port_vga_enable_3_hwtcl            : string  := "false";
			bridge_port_ssid_support_3_hwtcl          : string  := "false";
			ssvid_3_hwtcl                             : integer := 0;
			ssid_3_hwtcl                              : integer := 0;
			porttype_func4_hwtcl                      : string  := "Native endpoint";
			bar0_size_mask_4_hwtcl                    : integer := 28;
			bar0_io_space_4_hwtcl                     : string  := "Disabled";
			bar0_64bit_mem_space_4_hwtcl              : string  := "Enabled";
			bar0_prefetchable_4_hwtcl                 : string  := "Enabled";
			bar1_size_mask_4_hwtcl                    : integer := 0;
			bar1_io_space_4_hwtcl                     : string  := "Disabled";
			bar1_prefetchable_4_hwtcl                 : string  := "Disabled";
			bar2_size_mask_4_hwtcl                    : integer := 0;
			bar2_io_space_4_hwtcl                     : string  := "Disabled";
			bar2_64bit_mem_space_4_hwtcl              : string  := "Disabled";
			bar2_prefetchable_4_hwtcl                 : string  := "Disabled";
			bar3_size_mask_4_hwtcl                    : integer := 0;
			bar3_io_space_4_hwtcl                     : string  := "Disabled";
			bar3_prefetchable_4_hwtcl                 : string  := "Disabled";
			bar4_size_mask_4_hwtcl                    : integer := 0;
			bar4_io_space_4_hwtcl                     : string  := "Disabled";
			bar4_64bit_mem_space_4_hwtcl              : string  := "Disabled";
			bar4_prefetchable_4_hwtcl                 : string  := "Disabled";
			bar5_size_mask_4_hwtcl                    : integer := 0;
			bar5_io_space_4_hwtcl                     : string  := "Disabled";
			bar5_prefetchable_4_hwtcl                 : string  := "Disabled";
			expansion_base_address_register_4_hwtcl   : integer := 0;
			vendor_id_4_hwtcl                         : integer := 0;
			device_id_4_hwtcl                         : integer := 1;
			revision_id_4_hwtcl                       : integer := 1;
			class_code_4_hwtcl                        : integer := 0;
			subsystem_vendor_id_4_hwtcl               : integer := 0;
			subsystem_device_id_4_hwtcl               : integer := 0;
			max_payload_size_4_hwtcl                  : integer := 128;
			extend_tag_field_4_hwtcl                  : string  := "32";
			completion_timeout_4_hwtcl                : string  := "ABCD";
			enable_completion_timeout_disable_4_hwtcl : integer := 1;
			flr_capability_4_hwtcl                    : integer := 0;
			use_aer_4_hwtcl                           : integer := 0;
			ecrc_check_capable_4_hwtcl                : integer := 0;
			ecrc_gen_capable_4_hwtcl                  : integer := 0;
			dll_active_report_support_4_hwtcl         : integer := 0;
			surprise_down_error_support_4_hwtcl       : integer := 0;
			msi_multi_message_capable_4_hwtcl         : string  := "4";
			msi_64bit_addressing_capable_4_hwtcl      : string  := "true";
			msi_masking_capable_4_hwtcl               : string  := "false";
			msi_support_4_hwtcl                       : string  := "true";
			enable_function_msix_support_4_hwtcl      : integer := 0;
			msix_table_size_4_hwtcl                   : integer := 0;
			msix_table_offset_4_hwtcl                 : string  := "0";
			msix_table_bir_4_hwtcl                    : integer := 0;
			msix_pba_offset_4_hwtcl                   : string  := "0";
			msix_pba_bir_4_hwtcl                      : integer := 0;
			interrupt_pin_4_hwtcl                     : string  := "inta";
			slot_power_scale_4_hwtcl                  : integer := 0;
			slot_power_limit_4_hwtcl                  : integer := 0;
			slot_number_4_hwtcl                       : integer := 0;
			rx_ei_l0s_4_hwtcl                         : integer := 0;
			endpoint_l0_latency_4_hwtcl               : integer := 0;
			endpoint_l1_latency_4_hwtcl               : integer := 0;
			maximum_current_4_hwtcl                   : integer := 0;
			disable_snoop_packet_4_hwtcl              : string  := "false";
			bridge_port_vga_enable_4_hwtcl            : string  := "false";
			bridge_port_ssid_support_4_hwtcl          : string  := "false";
			ssvid_4_hwtcl                             : integer := 0;
			ssid_4_hwtcl                              : integer := 0;
			porttype_func5_hwtcl                      : string  := "Native endpoint";
			bar0_size_mask_5_hwtcl                    : integer := 28;
			bar0_io_space_5_hwtcl                     : string  := "Disabled";
			bar0_64bit_mem_space_5_hwtcl              : string  := "Enabled";
			bar0_prefetchable_5_hwtcl                 : string  := "Enabled";
			bar1_size_mask_5_hwtcl                    : integer := 0;
			bar1_io_space_5_hwtcl                     : string  := "Disabled";
			bar1_prefetchable_5_hwtcl                 : string  := "Disabled";
			bar2_size_mask_5_hwtcl                    : integer := 0;
			bar2_io_space_5_hwtcl                     : string  := "Disabled";
			bar2_64bit_mem_space_5_hwtcl              : string  := "Disabled";
			bar2_prefetchable_5_hwtcl                 : string  := "Disabled";
			bar3_size_mask_5_hwtcl                    : integer := 0;
			bar3_io_space_5_hwtcl                     : string  := "Disabled";
			bar3_prefetchable_5_hwtcl                 : string  := "Disabled";
			bar4_size_mask_5_hwtcl                    : integer := 0;
			bar4_io_space_5_hwtcl                     : string  := "Disabled";
			bar4_64bit_mem_space_5_hwtcl              : string  := "Disabled";
			bar4_prefetchable_5_hwtcl                 : string  := "Disabled";
			bar5_size_mask_5_hwtcl                    : integer := 0;
			bar5_io_space_5_hwtcl                     : string  := "Disabled";
			bar5_prefetchable_5_hwtcl                 : string  := "Disabled";
			expansion_base_address_register_5_hwtcl   : integer := 0;
			vendor_id_5_hwtcl                         : integer := 0;
			device_id_5_hwtcl                         : integer := 1;
			revision_id_5_hwtcl                       : integer := 1;
			class_code_5_hwtcl                        : integer := 0;
			subsystem_vendor_id_5_hwtcl               : integer := 0;
			subsystem_device_id_5_hwtcl               : integer := 0;
			max_payload_size_5_hwtcl                  : integer := 128;
			extend_tag_field_5_hwtcl                  : string  := "32";
			completion_timeout_5_hwtcl                : string  := "ABCD";
			enable_completion_timeout_disable_5_hwtcl : integer := 1;
			flr_capability_5_hwtcl                    : integer := 0;
			use_aer_5_hwtcl                           : integer := 0;
			ecrc_check_capable_5_hwtcl                : integer := 0;
			ecrc_gen_capable_5_hwtcl                  : integer := 0;
			dll_active_report_support_5_hwtcl         : integer := 0;
			surprise_down_error_support_5_hwtcl       : integer := 0;
			msi_multi_message_capable_5_hwtcl         : string  := "4";
			msi_64bit_addressing_capable_5_hwtcl      : string  := "true";
			msi_masking_capable_5_hwtcl               : string  := "false";
			msi_support_5_hwtcl                       : string  := "true";
			enable_function_msix_support_5_hwtcl      : integer := 0;
			msix_table_size_5_hwtcl                   : integer := 0;
			msix_table_offset_5_hwtcl                 : string  := "0";
			msix_table_bir_5_hwtcl                    : integer := 0;
			msix_pba_offset_5_hwtcl                   : string  := "0";
			msix_pba_bir_5_hwtcl                      : integer := 0;
			interrupt_pin_5_hwtcl                     : string  := "inta";
			slot_power_scale_5_hwtcl                  : integer := 0;
			slot_power_limit_5_hwtcl                  : integer := 0;
			slot_number_5_hwtcl                       : integer := 0;
			rx_ei_l0s_5_hwtcl                         : integer := 0;
			endpoint_l0_latency_5_hwtcl               : integer := 0;
			endpoint_l1_latency_5_hwtcl               : integer := 0;
			maximum_current_5_hwtcl                   : integer := 0;
			disable_snoop_packet_5_hwtcl              : string  := "false";
			bridge_port_vga_enable_5_hwtcl            : string  := "false";
			bridge_port_ssid_support_5_hwtcl          : string  := "false";
			ssvid_5_hwtcl                             : integer := 0;
			ssid_5_hwtcl                              : integer := 0;
			porttype_func6_hwtcl                      : string  := "Native endpoint";
			bar0_size_mask_6_hwtcl                    : integer := 28;
			bar0_io_space_6_hwtcl                     : string  := "Disabled";
			bar0_64bit_mem_space_6_hwtcl              : string  := "Enabled";
			bar0_prefetchable_6_hwtcl                 : string  := "Enabled";
			bar1_size_mask_6_hwtcl                    : integer := 0;
			bar1_io_space_6_hwtcl                     : string  := "Disabled";
			bar1_prefetchable_6_hwtcl                 : string  := "Disabled";
			bar2_size_mask_6_hwtcl                    : integer := 0;
			bar2_io_space_6_hwtcl                     : string  := "Disabled";
			bar2_64bit_mem_space_6_hwtcl              : string  := "Disabled";
			bar2_prefetchable_6_hwtcl                 : string  := "Disabled";
			bar3_size_mask_6_hwtcl                    : integer := 0;
			bar3_io_space_6_hwtcl                     : string  := "Disabled";
			bar3_prefetchable_6_hwtcl                 : string  := "Disabled";
			bar4_size_mask_6_hwtcl                    : integer := 0;
			bar4_io_space_6_hwtcl                     : string  := "Disabled";
			bar4_64bit_mem_space_6_hwtcl              : string  := "Disabled";
			bar4_prefetchable_6_hwtcl                 : string  := "Disabled";
			bar5_size_mask_6_hwtcl                    : integer := 0;
			bar5_io_space_6_hwtcl                     : string  := "Disabled";
			bar5_prefetchable_6_hwtcl                 : string  := "Disabled";
			expansion_base_address_register_6_hwtcl   : integer := 0;
			vendor_id_6_hwtcl                         : integer := 0;
			device_id_6_hwtcl                         : integer := 1;
			revision_id_6_hwtcl                       : integer := 1;
			class_code_6_hwtcl                        : integer := 0;
			subsystem_vendor_id_6_hwtcl               : integer := 0;
			subsystem_device_id_6_hwtcl               : integer := 0;
			max_payload_size_6_hwtcl                  : integer := 128;
			extend_tag_field_6_hwtcl                  : string  := "32";
			completion_timeout_6_hwtcl                : string  := "ABCD";
			enable_completion_timeout_disable_6_hwtcl : integer := 1;
			flr_capability_6_hwtcl                    : integer := 0;
			use_aer_6_hwtcl                           : integer := 0;
			ecrc_check_capable_6_hwtcl                : integer := 0;
			ecrc_gen_capable_6_hwtcl                  : integer := 0;
			dll_active_report_support_6_hwtcl         : integer := 0;
			surprise_down_error_support_6_hwtcl       : integer := 0;
			msi_multi_message_capable_6_hwtcl         : string  := "4";
			msi_64bit_addressing_capable_6_hwtcl      : string  := "true";
			msi_masking_capable_6_hwtcl               : string  := "false";
			msi_support_6_hwtcl                       : string  := "true";
			enable_function_msix_support_6_hwtcl      : integer := 0;
			msix_table_size_6_hwtcl                   : integer := 0;
			msix_table_offset_6_hwtcl                 : string  := "0";
			msix_table_bir_6_hwtcl                    : integer := 0;
			msix_pba_offset_6_hwtcl                   : string  := "0";
			msix_pba_bir_6_hwtcl                      : integer := 0;
			interrupt_pin_6_hwtcl                     : string  := "inta";
			slot_power_scale_6_hwtcl                  : integer := 0;
			slot_power_limit_6_hwtcl                  : integer := 0;
			slot_number_6_hwtcl                       : integer := 0;
			rx_ei_l0s_6_hwtcl                         : integer := 0;
			endpoint_l0_latency_6_hwtcl               : integer := 0;
			endpoint_l1_latency_6_hwtcl               : integer := 0;
			maximum_current_6_hwtcl                   : integer := 0;
			disable_snoop_packet_6_hwtcl              : string  := "false";
			bridge_port_vga_enable_6_hwtcl            : string  := "false";
			bridge_port_ssid_support_6_hwtcl          : string  := "false";
			ssvid_6_hwtcl                             : integer := 0;
			ssid_6_hwtcl                              : integer := 0;
			porttype_func7_hwtcl                      : string  := "Native endpoint";
			bar0_size_mask_7_hwtcl                    : integer := 28;
			bar0_io_space_7_hwtcl                     : string  := "Disabled";
			bar0_64bit_mem_space_7_hwtcl              : string  := "Enabled";
			bar0_prefetchable_7_hwtcl                 : string  := "Enabled";
			bar1_size_mask_7_hwtcl                    : integer := 0;
			bar1_io_space_7_hwtcl                     : string  := "Disabled";
			bar1_prefetchable_7_hwtcl                 : string  := "Disabled";
			bar2_size_mask_7_hwtcl                    : integer := 0;
			bar2_io_space_7_hwtcl                     : string  := "Disabled";
			bar2_64bit_mem_space_7_hwtcl              : string  := "Disabled";
			bar2_prefetchable_7_hwtcl                 : string  := "Disabled";
			bar3_size_mask_7_hwtcl                    : integer := 0;
			bar3_io_space_7_hwtcl                     : string  := "Disabled";
			bar3_prefetchable_7_hwtcl                 : string  := "Disabled";
			bar4_size_mask_7_hwtcl                    : integer := 0;
			bar4_io_space_7_hwtcl                     : string  := "Disabled";
			bar4_64bit_mem_space_7_hwtcl              : string  := "Disabled";
			bar4_prefetchable_7_hwtcl                 : string  := "Disabled";
			bar5_size_mask_7_hwtcl                    : integer := 0;
			bar5_io_space_7_hwtcl                     : string  := "Disabled";
			bar5_prefetchable_7_hwtcl                 : string  := "Disabled";
			expansion_base_address_register_7_hwtcl   : integer := 0;
			vendor_id_7_hwtcl                         : integer := 0;
			device_id_7_hwtcl                         : integer := 1;
			revision_id_7_hwtcl                       : integer := 1;
			class_code_7_hwtcl                        : integer := 0;
			subsystem_vendor_id_7_hwtcl               : integer := 0;
			subsystem_device_id_7_hwtcl               : integer := 0;
			max_payload_size_7_hwtcl                  : integer := 128;
			extend_tag_field_7_hwtcl                  : string  := "32";
			completion_timeout_7_hwtcl                : string  := "ABCD";
			enable_completion_timeout_disable_7_hwtcl : integer := 1;
			flr_capability_7_hwtcl                    : integer := 0;
			use_aer_7_hwtcl                           : integer := 0;
			ecrc_check_capable_7_hwtcl                : integer := 0;
			ecrc_gen_capable_7_hwtcl                  : integer := 0;
			dll_active_report_support_7_hwtcl         : integer := 0;
			surprise_down_error_support_7_hwtcl       : integer := 0;
			msi_multi_message_capable_7_hwtcl         : string  := "4";
			msi_64bit_addressing_capable_7_hwtcl      : string  := "true";
			msi_masking_capable_7_hwtcl               : string  := "false";
			msi_support_7_hwtcl                       : string  := "true";
			enable_function_msix_support_7_hwtcl      : integer := 0;
			msix_table_size_7_hwtcl                   : integer := 0;
			msix_table_offset_7_hwtcl                 : string  := "0";
			msix_table_bir_7_hwtcl                    : integer := 0;
			msix_pba_offset_7_hwtcl                   : string  := "0";
			msix_pba_bir_7_hwtcl                      : integer := 0;
			interrupt_pin_7_hwtcl                     : string  := "inta";
			slot_power_scale_7_hwtcl                  : integer := 0;
			slot_power_limit_7_hwtcl                  : integer := 0;
			slot_number_7_hwtcl                       : integer := 0;
			rx_ei_l0s_7_hwtcl                         : integer := 0;
			endpoint_l0_latency_7_hwtcl               : integer := 0;
			endpoint_l1_latency_7_hwtcl               : integer := 0;
			maximum_current_7_hwtcl                   : integer := 0;
			disable_snoop_packet_7_hwtcl              : string  := "false";
			bridge_port_vga_enable_7_hwtcl            : string  := "false";
			bridge_port_ssid_support_7_hwtcl          : string  := "false";
			ssvid_7_hwtcl                             : integer := 0;
			ssid_7_hwtcl                              : integer := 0;
			rpre_emph_a_val_hwtcl                     : integer := 11;
			rpre_emph_b_val_hwtcl                     : integer := 0;
			rpre_emph_c_val_hwtcl                     : integer := 22;
			rpre_emph_d_val_hwtcl                     : integer := 12;
			rpre_emph_e_val_hwtcl                     : integer := 21;
			rvod_sel_a_val_hwtcl                      : integer := 50;
			rvod_sel_b_val_hwtcl                      : integer := 34;
			rvod_sel_c_val_hwtcl                      : integer := 50;
			rvod_sel_d_val_hwtcl                      : integer := 50;
			rvod_sel_e_val_hwtcl                      : integer := 9
		);
		port (
			npor                   : in  std_logic                      := 'X';             -- npor
			pin_perst              : in  std_logic                      := 'X';             -- pin_perst
			test_in                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- test_in
			simu_mode_pipe         : in  std_logic                      := 'X';             -- simu_mode_pipe
			pld_clk                : in  std_logic                      := 'X';             -- clk
			coreclkout             : out std_logic;                                         -- clk
			refclk                 : in  std_logic                      := 'X';             -- clk
			rx_in0                 : in  std_logic                      := 'X';             -- rx_in0
			rx_in1                 : in  std_logic                      := 'X';             -- rx_in1
			rx_in2                 : in  std_logic                      := 'X';             -- rx_in2
			rx_in3                 : in  std_logic                      := 'X';             -- rx_in3
			tx_out0                : out std_logic;                                         -- tx_out0
			tx_out1                : out std_logic;                                         -- tx_out1
			tx_out2                : out std_logic;                                         -- tx_out2
			tx_out3                : out std_logic;                                         -- tx_out3
			rx_st_valid            : out std_logic;                                         -- valid
			rx_st_sop              : out std_logic;                                         -- startofpacket
			rx_st_eop              : out std_logic;                                         -- endofpacket
			rx_st_ready            : in  std_logic                      := 'X';             -- ready
			rx_st_err              : out std_logic;                                         -- error
			rx_st_data             : out std_logic_vector(63 downto 0);                     -- data
			rx_st_bar              : out std_logic_vector(7 downto 0);                      -- rx_st_bar
			rx_st_mask             : in  std_logic                      := 'X';             -- rx_st_mask
			tx_st_valid            : in  std_logic                      := 'X';             -- valid
			tx_st_sop              : in  std_logic                      := 'X';             -- startofpacket
			tx_st_eop              : in  std_logic                      := 'X';             -- endofpacket
			tx_st_ready            : out std_logic;                                         -- ready
			tx_st_err              : in  std_logic                      := 'X';             -- error
			tx_st_data             : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- data
			tx_fifo_empty          : out std_logic;                                         -- fifo_empty
			tx_cred_datafccp       : out std_logic_vector(11 downto 0);                     -- tx_cred_datafccp
			tx_cred_datafcnp       : out std_logic_vector(11 downto 0);                     -- tx_cred_datafcnp
			tx_cred_datafcp        : out std_logic_vector(11 downto 0);                     -- tx_cred_datafcp
			tx_cred_fchipcons      : out std_logic_vector(5 downto 0);                      -- tx_cred_fchipcons
			tx_cred_fcinfinite     : out std_logic_vector(5 downto 0);                      -- tx_cred_fcinfinite
			tx_cred_hdrfccp        : out std_logic_vector(7 downto 0);                      -- tx_cred_hdrfccp
			tx_cred_hdrfcnp        : out std_logic_vector(7 downto 0);                      -- tx_cred_hdrfcnp
			tx_cred_hdrfcp         : out std_logic_vector(7 downto 0);                      -- tx_cred_hdrfcp
			sim_pipe_pclk_in       : in  std_logic                      := 'X';             -- sim_pipe_pclk_in
			sim_pipe_rate          : out std_logic_vector(1 downto 0);                      -- sim_pipe_rate
			sim_ltssmstate         : out std_logic_vector(4 downto 0);                      -- sim_ltssmstate
			eidleinfersel0         : out std_logic_vector(2 downto 0);                      -- eidleinfersel0
			eidleinfersel1         : out std_logic_vector(2 downto 0);                      -- eidleinfersel1
			eidleinfersel2         : out std_logic_vector(2 downto 0);                      -- eidleinfersel2
			eidleinfersel3         : out std_logic_vector(2 downto 0);                      -- eidleinfersel3
			powerdown0             : out std_logic_vector(1 downto 0);                      -- powerdown0
			powerdown1             : out std_logic_vector(1 downto 0);                      -- powerdown1
			powerdown2             : out std_logic_vector(1 downto 0);                      -- powerdown2
			powerdown3             : out std_logic_vector(1 downto 0);                      -- powerdown3
			rxpolarity0            : out std_logic;                                         -- rxpolarity0
			rxpolarity1            : out std_logic;                                         -- rxpolarity1
			rxpolarity2            : out std_logic;                                         -- rxpolarity2
			rxpolarity3            : out std_logic;                                         -- rxpolarity3
			txcompl0               : out std_logic;                                         -- txcompl0
			txcompl1               : out std_logic;                                         -- txcompl1
			txcompl2               : out std_logic;                                         -- txcompl2
			txcompl3               : out std_logic;                                         -- txcompl3
			txdata0                : out std_logic_vector(7 downto 0);                      -- txdata0
			txdata1                : out std_logic_vector(7 downto 0);                      -- txdata1
			txdata2                : out std_logic_vector(7 downto 0);                      -- txdata2
			txdata3                : out std_logic_vector(7 downto 0);                      -- txdata3
			txdatak0               : out std_logic;                                         -- txdatak0
			txdatak1               : out std_logic;                                         -- txdatak1
			txdatak2               : out std_logic;                                         -- txdatak2
			txdatak3               : out std_logic;                                         -- txdatak3
			txdetectrx0            : out std_logic;                                         -- txdetectrx0
			txdetectrx1            : out std_logic;                                         -- txdetectrx1
			txdetectrx2            : out std_logic;                                         -- txdetectrx2
			txdetectrx3            : out std_logic;                                         -- txdetectrx3
			txelecidle0            : out std_logic;                                         -- txelecidle0
			txelecidle1            : out std_logic;                                         -- txelecidle1
			txelecidle2            : out std_logic;                                         -- txelecidle2
			txelecidle3            : out std_logic;                                         -- txelecidle3
			txswing0               : out std_logic;                                         -- txswing0
			txswing1               : out std_logic;                                         -- txswing1
			txswing2               : out std_logic;                                         -- txswing2
			txswing3               : out std_logic;                                         -- txswing3
			txmargin0              : out std_logic_vector(2 downto 0);                      -- txmargin0
			txmargin1              : out std_logic_vector(2 downto 0);                      -- txmargin1
			txmargin2              : out std_logic_vector(2 downto 0);                      -- txmargin2
			txmargin3              : out std_logic_vector(2 downto 0);                      -- txmargin3
			txdeemph0              : out std_logic;                                         -- txdeemph0
			txdeemph1              : out std_logic;                                         -- txdeemph1
			txdeemph2              : out std_logic;                                         -- txdeemph2
			txdeemph3              : out std_logic;                                         -- txdeemph3
			phystatus0             : in  std_logic                      := 'X';             -- phystatus0
			phystatus1             : in  std_logic                      := 'X';             -- phystatus1
			phystatus2             : in  std_logic                      := 'X';             -- phystatus2
			phystatus3             : in  std_logic                      := 'X';             -- phystatus3
			rxdata0                : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rxdata0
			rxdata1                : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rxdata1
			rxdata2                : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rxdata2
			rxdata3                : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rxdata3
			rxdatak0               : in  std_logic                      := 'X';             -- rxdatak0
			rxdatak1               : in  std_logic                      := 'X';             -- rxdatak1
			rxdatak2               : in  std_logic                      := 'X';             -- rxdatak2
			rxdatak3               : in  std_logic                      := 'X';             -- rxdatak3
			rxelecidle0            : in  std_logic                      := 'X';             -- rxelecidle0
			rxelecidle1            : in  std_logic                      := 'X';             -- rxelecidle1
			rxelecidle2            : in  std_logic                      := 'X';             -- rxelecidle2
			rxelecidle3            : in  std_logic                      := 'X';             -- rxelecidle3
			rxstatus0              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rxstatus0
			rxstatus1              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rxstatus1
			rxstatus2              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rxstatus2
			rxstatus3              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rxstatus3
			rxvalid0               : in  std_logic                      := 'X';             -- rxvalid0
			rxvalid1               : in  std_logic                      := 'X';             -- rxvalid1
			rxvalid2               : in  std_logic                      := 'X';             -- rxvalid2
			rxvalid3               : in  std_logic                      := 'X';             -- rxvalid3
			reset_status           : out std_logic;                                         -- reset_status
			serdes_pll_locked      : out std_logic;                                         -- serdes_pll_locked
			pld_clk_inuse          : out std_logic;                                         -- pld_clk_inuse
			pld_core_ready         : in  std_logic                      := 'X';             -- pld_core_ready
			testin_zero            : out std_logic;                                         -- testin_zero
			lmi_addr               : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- lmi_addr
			lmi_din                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- lmi_din
			lmi_rden               : in  std_logic                      := 'X';             -- lmi_rden
			lmi_wren               : in  std_logic                      := 'X';             -- lmi_wren
			lmi_ack                : out std_logic;                                         -- lmi_ack
			lmi_dout               : out std_logic_vector(31 downto 0);                     -- lmi_dout
			pm_auxpwr              : in  std_logic                      := 'X';             -- pm_auxpwr
			pm_data                : in  std_logic_vector(9 downto 0)   := (others => 'X'); -- pm_data
			pme_to_cr              : in  std_logic                      := 'X';             -- pme_to_cr
			pm_event               : in  std_logic                      := 'X';             -- pm_event
			pme_to_sr              : out std_logic;                                         -- pme_to_sr
			reconfig_to_xcvr       : in  std_logic_vector(349 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr     : out std_logic_vector(229 downto 0);                    -- reconfig_from_xcvr
			app_msi_num            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- app_msi_num
			app_msi_req            : in  std_logic                      := 'X';             -- app_msi_req
			app_msi_tc             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- app_msi_tc
			app_msi_ack            : out std_logic;                                         -- app_msi_ack
			app_int_sts_vec        : in  std_logic                      := 'X';             -- app_int_sts
			tl_hpg_ctrl_er         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- hpg_ctrler
			tl_cfg_ctl             : out std_logic_vector(31 downto 0);                     -- tl_cfg_ctl
			cpl_err                : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- cpl_err
			tl_cfg_add             : out std_logic_vector(3 downto 0);                      -- tl_cfg_add
			tl_cfg_ctl_wr          : out std_logic;                                         -- tl_cfg_ctl_wr
			tl_cfg_sts_wr          : out std_logic;                                         -- tl_cfg_sts_wr
			tl_cfg_sts             : out std_logic_vector(52 downto 0);                     -- tl_cfg_sts
			cpl_pending            : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- cpl_pending
			derr_cor_ext_rcv0      : out std_logic;                                         -- derr_cor_ext_rcv
			derr_cor_ext_rpl       : out std_logic;                                         -- derr_cor_ext_rpl
			derr_rpl               : out std_logic;                                         -- derr_rpl
			dlup_exit              : out std_logic;                                         -- dlup_exit
			dl_ltssm               : out std_logic_vector(4 downto 0);                      -- ltssmstate
			ev128ns                : out std_logic;                                         -- ev128ns
			ev1us                  : out std_logic;                                         -- ev1us
			hotrst_exit            : out std_logic;                                         -- hotrst_exit
			int_status             : out std_logic_vector(3 downto 0);                      -- int_status
			l2_exit                : out std_logic;                                         -- l2_exit
			lane_act               : out std_logic_vector(3 downto 0);                      -- lane_act
			ko_cpl_spc_header      : out std_logic_vector(7 downto 0);                      -- ko_cpl_spc_header
			ko_cpl_spc_data        : out std_logic_vector(11 downto 0);                     -- ko_cpl_spc_data
			dl_current_speed       : out std_logic_vector(1 downto 0);                      -- currentspeed
			rx_in4                 : in  std_logic                      := 'X';             -- rx_in4
			rx_in5                 : in  std_logic                      := 'X';             -- rx_in5
			rx_in6                 : in  std_logic                      := 'X';             -- rx_in6
			rx_in7                 : in  std_logic                      := 'X';             -- rx_in7
			tx_out4                : out std_logic;                                         -- tx_out4
			tx_out5                : out std_logic;                                         -- tx_out5
			tx_out6                : out std_logic;                                         -- tx_out6
			tx_out7                : out std_logic;                                         -- tx_out7
			rx_st_empty            : out std_logic;                                         -- rx_st_empty
			rx_fifo_empty          : out std_logic;                                         -- rx_fifo_empty
			rx_fifo_full           : out std_logic;                                         -- rx_fifo_full
			rx_bar_dec_func_num    : out std_logic_vector(2 downto 0);                      -- rx_bar_dec_func_num
			rx_st_be               : out std_logic_vector(7 downto 0);                      -- rx_st_be
			tx_st_empty            : in  std_logic                      := 'X';             -- tx_st_empty
			tx_fifo_full           : out std_logic;                                         -- tx_fifo_full
			tx_fifo_rdp            : out std_logic_vector(3 downto 0);                      -- tx_fifo_rdp
			tx_fifo_wrp            : out std_logic_vector(3 downto 0);                      -- tx_fifo_wrp
			eidleinfersel4         : out std_logic_vector(2 downto 0);                      -- eidleinfersel4
			eidleinfersel5         : out std_logic_vector(2 downto 0);                      -- eidleinfersel5
			eidleinfersel6         : out std_logic_vector(2 downto 0);                      -- eidleinfersel6
			eidleinfersel7         : out std_logic_vector(2 downto 0);                      -- eidleinfersel7
			powerdown4             : out std_logic_vector(1 downto 0);                      -- powerdown4
			powerdown5             : out std_logic_vector(1 downto 0);                      -- powerdown5
			powerdown6             : out std_logic_vector(1 downto 0);                      -- powerdown6
			powerdown7             : out std_logic_vector(1 downto 0);                      -- powerdown7
			rxpolarity4            : out std_logic;                                         -- rxpolarity4
			rxpolarity5            : out std_logic;                                         -- rxpolarity5
			rxpolarity6            : out std_logic;                                         -- rxpolarity6
			rxpolarity7            : out std_logic;                                         -- rxpolarity7
			txcompl4               : out std_logic;                                         -- txcompl4
			txcompl5               : out std_logic;                                         -- txcompl5
			txcompl6               : out std_logic;                                         -- txcompl6
			txcompl7               : out std_logic;                                         -- txcompl7
			txdata4                : out std_logic_vector(7 downto 0);                      -- txdata4
			txdata5                : out std_logic_vector(7 downto 0);                      -- txdata5
			txdata6                : out std_logic_vector(7 downto 0);                      -- txdata6
			txdata7                : out std_logic_vector(7 downto 0);                      -- txdata7
			txdatak4               : out std_logic;                                         -- txdatak4
			txdatak5               : out std_logic;                                         -- txdatak5
			txdatak6               : out std_logic;                                         -- txdatak6
			txdatak7               : out std_logic;                                         -- txdatak7
			txdetectrx4            : out std_logic;                                         -- txdetectrx4
			txdetectrx5            : out std_logic;                                         -- txdetectrx5
			txdetectrx6            : out std_logic;                                         -- txdetectrx6
			txdetectrx7            : out std_logic;                                         -- txdetectrx7
			txelecidle4            : out std_logic;                                         -- txelecidle4
			txelecidle5            : out std_logic;                                         -- txelecidle5
			txelecidle6            : out std_logic;                                         -- txelecidle6
			txelecidle7            : out std_logic;                                         -- txelecidle7
			txswing4               : out std_logic;                                         -- txswing4
			txswing5               : out std_logic;                                         -- txswing5
			txswing6               : out std_logic;                                         -- txswing6
			txswing7               : out std_logic;                                         -- txswing7
			txmargin4              : out std_logic_vector(2 downto 0);                      -- txmargin4
			txmargin5              : out std_logic_vector(2 downto 0);                      -- txmargin5
			txmargin6              : out std_logic_vector(2 downto 0);                      -- txmargin6
			txmargin7              : out std_logic_vector(2 downto 0);                      -- txmargin7
			txdeemph4              : out std_logic;                                         -- txdeemph4
			txdeemph5              : out std_logic;                                         -- txdeemph5
			txdeemph6              : out std_logic;                                         -- txdeemph6
			txdeemph7              : out std_logic;                                         -- txdeemph7
			phystatus4             : in  std_logic                      := 'X';             -- phystatus4
			phystatus5             : in  std_logic                      := 'X';             -- phystatus5
			phystatus6             : in  std_logic                      := 'X';             -- phystatus6
			phystatus7             : in  std_logic                      := 'X';             -- phystatus7
			rxdata4                : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rxdata4
			rxdata5                : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rxdata5
			rxdata6                : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rxdata6
			rxdata7                : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rxdata7
			rxdatak4               : in  std_logic                      := 'X';             -- rxdatak4
			rxdatak5               : in  std_logic                      := 'X';             -- rxdatak5
			rxdatak6               : in  std_logic                      := 'X';             -- rxdatak6
			rxdatak7               : in  std_logic                      := 'X';             -- rxdatak7
			rxelecidle4            : in  std_logic                      := 'X';             -- rxelecidle4
			rxelecidle5            : in  std_logic                      := 'X';             -- rxelecidle5
			rxelecidle6            : in  std_logic                      := 'X';             -- rxelecidle6
			rxelecidle7            : in  std_logic                      := 'X';             -- rxelecidle7
			rxstatus4              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rxstatus4
			rxstatus5              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rxstatus5
			rxstatus6              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rxstatus6
			rxstatus7              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rxstatus7
			rxvalid4               : in  std_logic                      := 'X';             -- rxvalid4
			rxvalid5               : in  std_logic                      := 'X';             -- rxvalid5
			rxvalid6               : in  std_logic                      := 'X';             -- rxvalid6
			rxvalid7               : in  std_logic                      := 'X';             -- rxvalid7
			sim_pipe_pclk_out      : out std_logic;                                         -- sim_pipe_pclk_out
			pm_event_func          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- pm_event_func
			hip_reconfig_clk       : in  std_logic                      := 'X';             -- hip_reconfig_clk
			hip_reconfig_rst_n     : in  std_logic                      := 'X';             -- hip_reconfig_rst_n
			hip_reconfig_address   : in  std_logic_vector(9 downto 0)   := (others => 'X'); -- hip_reconfig_address
			hip_reconfig_byte_en   : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- hip_reconfig_byte_en
			hip_reconfig_read      : in  std_logic                      := 'X';             -- hip_reconfig_read
			hip_reconfig_readdata  : out std_logic_vector(15 downto 0);                     -- hip_reconfig_readdata
			hip_reconfig_write     : in  std_logic                      := 'X';             -- hip_reconfig_write
			hip_reconfig_writedata : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- hip_reconfig_writedata
			ser_shift_load         : in  std_logic                      := 'X';             -- ser_shift_load
			interface_sel          : in  std_logic                      := 'X';             -- interface_sel
			app_msi_func           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- app_msi_func
			serr_out               : out std_logic;                                         -- serr_out
			aer_msi_num            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- aer_msi_num
			pex_msi_num            : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- pex_msi_num
			cpl_err_func           : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- cpl_err_func
		);
	end component altpcie_cv_hip_ast_hwtcl;

begin

	pcie_inst : component altpcie_cv_hip_ast_hwtcl
		generic map (
			ACDS_VERSION_HWTCL                        => "18.1",
			lane_mask_hwtcl                           => "x4",
			gen12_lane_rate_mode_hwtcl                => "Gen1 (2.5 Gbps)",
			pcie_spec_version_hwtcl                   => "2.1",
			ast_width_hwtcl                           => "Avalon-ST 64-bit",
			pll_refclk_freq_hwtcl                     => "100 MHz",
			set_pld_clk_x1_625MHz_hwtcl               => 0,
			in_cvp_mode_hwtcl                         => 0,
			hip_reconfig_hwtcl                        => 0,
			num_of_func_hwtcl                         => 1,
			use_crc_forwarding_hwtcl                  => 0,
			port_link_number_hwtcl                    => 1,
			slotclkcfg_hwtcl                          => 1,
			enable_slot_register_hwtcl                => 0,
			vsec_id_hwtcl                             => 4466,
			vsec_rev_hwtcl                            => 0,
			user_id_hwtcl                             => 0,
			porttype_func0_hwtcl                      => "Native endpoint",
			bar0_size_mask_0_hwtcl                    => 16,
			bar0_io_space_0_hwtcl                     => "Disabled",
			bar0_64bit_mem_space_0_hwtcl              => "Enabled",
			bar0_prefetchable_0_hwtcl                 => "Enabled",
			bar1_size_mask_0_hwtcl                    => 0,
			bar1_io_space_0_hwtcl                     => "Disabled",
			bar1_prefetchable_0_hwtcl                 => "Disabled",
			bar2_size_mask_0_hwtcl                    => 0,
			bar2_io_space_0_hwtcl                     => "Disabled",
			bar2_64bit_mem_space_0_hwtcl              => "Disabled",
			bar2_prefetchable_0_hwtcl                 => "Disabled",
			bar3_size_mask_0_hwtcl                    => 0,
			bar3_io_space_0_hwtcl                     => "Disabled",
			bar3_prefetchable_0_hwtcl                 => "Disabled",
			bar4_size_mask_0_hwtcl                    => 16,
			bar4_io_space_0_hwtcl                     => "Disabled",
			bar4_64bit_mem_space_0_hwtcl              => "Enabled",
			bar4_prefetchable_0_hwtcl                 => "Enabled",
			bar5_size_mask_0_hwtcl                    => 0,
			bar5_io_space_0_hwtcl                     => "Disabled",
			bar5_prefetchable_0_hwtcl                 => "Disabled",
			expansion_base_address_register_0_hwtcl   => 0,
			io_window_addr_width_hwtcl                => 0,
			prefetchable_mem_window_addr_width_hwtcl  => 0,
			vendor_id_0_hwtcl                         => 4466,
			device_id_0_hwtcl                         => 57347,
			revision_id_0_hwtcl                       => 1,
			class_code_0_hwtcl                        => 0,
			subsystem_vendor_id_0_hwtcl               => 0,
			subsystem_device_id_0_hwtcl               => 10337,
			max_payload_size_0_hwtcl                  => 256,
			extend_tag_field_0_hwtcl                  => "32",
			completion_timeout_0_hwtcl                => "ABCD",
			enable_completion_timeout_disable_0_hwtcl => 1,
			flr_capability_0_hwtcl                    => 0,
			use_aer_0_hwtcl                           => 0,
			ecrc_check_capable_0_hwtcl                => 0,
			ecrc_gen_capable_0_hwtcl                  => 0,
			dll_active_report_support_0_hwtcl         => 0,
			surprise_down_error_support_0_hwtcl       => 0,
			msi_multi_message_capable_0_hwtcl         => "1",
			msi_64bit_addressing_capable_0_hwtcl      => "true",
			msi_masking_capable_0_hwtcl               => "false",
			msi_support_0_hwtcl                       => "true",
			enable_function_msix_support_0_hwtcl      => 0,
			msix_table_size_0_hwtcl                   => 0,
			msix_table_offset_0_hwtcl                 => "0",
			msix_table_bir_0_hwtcl                    => 0,
			msix_pba_offset_0_hwtcl                   => "0",
			msix_pba_bir_0_hwtcl                      => 0,
			interrupt_pin_0_hwtcl                     => "inta",
			slot_power_scale_0_hwtcl                  => 0,
			slot_power_limit_0_hwtcl                  => 0,
			slot_number_0_hwtcl                       => 0,
			rx_ei_l0s_0_hwtcl                         => 0,
			endpoint_l0_latency_0_hwtcl               => 0,
			endpoint_l1_latency_0_hwtcl               => 0,
			reconfig_to_xcvr_width                    => 350,
			hip_hard_reset_hwtcl                      => 1,
			reconfig_from_xcvr_width                  => 230,
			single_rx_detect_hwtcl                    => 4,
			enable_l0s_aspm_hwtcl                     => "false",
			aspm_optionality_hwtcl                    => "true",
			enable_adapter_half_rate_mode_hwtcl       => "false",
			millisecond_cycle_count_hwtcl             => 124250,
			credit_buffer_allocation_aux_hwtcl        => "absolute",
			vc0_rx_flow_ctrl_posted_header_hwtcl      => 16,
			vc0_rx_flow_ctrl_posted_data_hwtcl        => 16,
			vc0_rx_flow_ctrl_nonposted_header_hwtcl   => 16,
			vc0_rx_flow_ctrl_nonposted_data_hwtcl     => 0,
			vc0_rx_flow_ctrl_compl_header_hwtcl       => 0,
			vc0_rx_flow_ctrl_compl_data_hwtcl         => 0,
			cpl_spc_header_hwtcl                      => 67,
			cpl_spc_data_hwtcl                        => 269,
			port_width_data_hwtcl                     => 64,
			bypass_clk_switch_hwtcl                   => "disable",
			cvp_rate_sel_hwtcl                        => "full_rate",
			cvp_data_compressed_hwtcl                 => "false",
			cvp_data_encrypted_hwtcl                  => "false",
			cvp_mode_reset_hwtcl                      => "false",
			cvp_clk_reset_hwtcl                       => "false",
			core_clk_sel_hwtcl                        => "pld_clk",
			enable_rx_buffer_checking_hwtcl           => "false",
			disable_link_x2_support_hwtcl             => "false",
			device_number_hwtcl                       => 0,
			pipex1_debug_sel_hwtcl                    => "disable",
			pclk_out_sel_hwtcl                        => "pclk",
			no_soft_reset_hwtcl                       => "false",
			d1_support_hwtcl                          => "false",
			d2_support_hwtcl                          => "false",
			d0_pme_hwtcl                              => "false",
			d1_pme_hwtcl                              => "false",
			d2_pme_hwtcl                              => "false",
			d3_hot_pme_hwtcl                          => "false",
			d3_cold_pme_hwtcl                         => "false",
			low_priority_vc_hwtcl                     => "single_vc",
			enable_l1_aspm_hwtcl                      => "false",
			l1_exit_latency_sameclock_hwtcl           => 0,
			l1_exit_latency_diffclock_hwtcl           => 0,
			hot_plug_support_hwtcl                    => 0,
			no_command_completed_hwtcl                => "false",
			eie_before_nfts_count_hwtcl               => 4,
			gen2_diffclock_nfts_count_hwtcl           => 255,
			gen2_sameclock_nfts_count_hwtcl           => 255,
			deemphasis_enable_hwtcl                   => "false",
			l0_exit_latency_sameclock_hwtcl           => 6,
			l0_exit_latency_diffclock_hwtcl           => 6,
			vc0_clk_enable_hwtcl                      => "true",
			register_pipe_signals_hwtcl               => "true",
			tx_cdc_almost_empty_hwtcl                 => 5,
			rx_l0s_count_idl_hwtcl                    => 0,
			cdc_dummy_insert_limit_hwtcl              => 11,
			ei_delay_powerdown_count_hwtcl            => 10,
			skp_os_schedule_count_hwtcl               => 0,
			fc_init_timer_hwtcl                       => 1024,
			l01_entry_latency_hwtcl                   => 31,
			flow_control_update_count_hwtcl           => 30,
			flow_control_timeout_count_hwtcl          => 200,
			retry_buffer_last_active_address_hwtcl    => 255,
			reserved_debug_hwtcl                      => 0,
			use_tl_cfg_sync_hwtcl                     => 1,
			diffclock_nfts_count_hwtcl                => 255,
			sameclock_nfts_count_hwtcl                => 255,
			l2_async_logic_hwtcl                      => "disable",
			rx_cdc_almost_full_hwtcl                  => 12,
			tx_cdc_almost_full_hwtcl                  => 11,
			indicator_hwtcl                           => 0,
			maximum_current_0_hwtcl                   => 0,
			disable_snoop_packet_0_hwtcl              => "false",
			bridge_port_vga_enable_0_hwtcl            => "false",
			bridge_port_ssid_support_0_hwtcl          => "false",
			ssvid_0_hwtcl                             => 0,
			ssid_0_hwtcl                              => 0,
			porttype_func1_hwtcl                      => "Native endpoint",
			bar0_size_mask_1_hwtcl                    => 28,
			bar0_io_space_1_hwtcl                     => "Disabled",
			bar0_64bit_mem_space_1_hwtcl              => "Enabled",
			bar0_prefetchable_1_hwtcl                 => "Enabled",
			bar1_size_mask_1_hwtcl                    => 0,
			bar1_io_space_1_hwtcl                     => "Disabled",
			bar1_prefetchable_1_hwtcl                 => "Disabled",
			bar2_size_mask_1_hwtcl                    => 0,
			bar2_io_space_1_hwtcl                     => "Disabled",
			bar2_64bit_mem_space_1_hwtcl              => "Disabled",
			bar2_prefetchable_1_hwtcl                 => "Disabled",
			bar3_size_mask_1_hwtcl                    => 0,
			bar3_io_space_1_hwtcl                     => "Disabled",
			bar3_prefetchable_1_hwtcl                 => "Disabled",
			bar4_size_mask_1_hwtcl                    => 0,
			bar4_io_space_1_hwtcl                     => "Disabled",
			bar4_64bit_mem_space_1_hwtcl              => "Disabled",
			bar4_prefetchable_1_hwtcl                 => "Disabled",
			bar5_size_mask_1_hwtcl                    => 0,
			bar5_io_space_1_hwtcl                     => "Disabled",
			bar5_prefetchable_1_hwtcl                 => "Disabled",
			expansion_base_address_register_1_hwtcl   => 0,
			vendor_id_1_hwtcl                         => 0,
			device_id_1_hwtcl                         => 1,
			revision_id_1_hwtcl                       => 1,
			class_code_1_hwtcl                        => 0,
			subsystem_vendor_id_1_hwtcl               => 0,
			subsystem_device_id_1_hwtcl               => 0,
			max_payload_size_1_hwtcl                  => 256,
			extend_tag_field_1_hwtcl                  => "32",
			completion_timeout_1_hwtcl                => "ABCD",
			enable_completion_timeout_disable_1_hwtcl => 1,
			flr_capability_1_hwtcl                    => 0,
			use_aer_1_hwtcl                           => 0,
			ecrc_check_capable_1_hwtcl                => 0,
			ecrc_gen_capable_1_hwtcl                  => 0,
			dll_active_report_support_1_hwtcl         => 0,
			surprise_down_error_support_1_hwtcl       => 0,
			msi_multi_message_capable_1_hwtcl         => "4",
			msi_64bit_addressing_capable_1_hwtcl      => "true",
			msi_masking_capable_1_hwtcl               => "false",
			msi_support_1_hwtcl                       => "true",
			enable_function_msix_support_1_hwtcl      => 0,
			msix_table_size_1_hwtcl                   => 0,
			msix_table_offset_1_hwtcl                 => "0",
			msix_table_bir_1_hwtcl                    => 0,
			msix_pba_offset_1_hwtcl                   => "0",
			msix_pba_bir_1_hwtcl                      => 0,
			interrupt_pin_1_hwtcl                     => "inta",
			slot_power_scale_1_hwtcl                  => 0,
			slot_power_limit_1_hwtcl                  => 0,
			slot_number_1_hwtcl                       => 0,
			rx_ei_l0s_1_hwtcl                         => 0,
			endpoint_l0_latency_1_hwtcl               => 0,
			endpoint_l1_latency_1_hwtcl               => 0,
			maximum_current_1_hwtcl                   => 0,
			disable_snoop_packet_1_hwtcl              => "false",
			bridge_port_vga_enable_1_hwtcl            => "false",
			bridge_port_ssid_support_1_hwtcl          => "false",
			ssvid_1_hwtcl                             => 0,
			ssid_1_hwtcl                              => 0,
			porttype_func2_hwtcl                      => "Native endpoint",
			bar0_size_mask_2_hwtcl                    => 28,
			bar0_io_space_2_hwtcl                     => "Disabled",
			bar0_64bit_mem_space_2_hwtcl              => "Enabled",
			bar0_prefetchable_2_hwtcl                 => "Enabled",
			bar1_size_mask_2_hwtcl                    => 0,
			bar1_io_space_2_hwtcl                     => "Disabled",
			bar1_prefetchable_2_hwtcl                 => "Disabled",
			bar2_size_mask_2_hwtcl                    => 0,
			bar2_io_space_2_hwtcl                     => "Disabled",
			bar2_64bit_mem_space_2_hwtcl              => "Disabled",
			bar2_prefetchable_2_hwtcl                 => "Disabled",
			bar3_size_mask_2_hwtcl                    => 0,
			bar3_io_space_2_hwtcl                     => "Disabled",
			bar3_prefetchable_2_hwtcl                 => "Disabled",
			bar4_size_mask_2_hwtcl                    => 0,
			bar4_io_space_2_hwtcl                     => "Disabled",
			bar4_64bit_mem_space_2_hwtcl              => "Disabled",
			bar4_prefetchable_2_hwtcl                 => "Disabled",
			bar5_size_mask_2_hwtcl                    => 0,
			bar5_io_space_2_hwtcl                     => "Disabled",
			bar5_prefetchable_2_hwtcl                 => "Disabled",
			expansion_base_address_register_2_hwtcl   => 0,
			vendor_id_2_hwtcl                         => 0,
			device_id_2_hwtcl                         => 1,
			revision_id_2_hwtcl                       => 1,
			class_code_2_hwtcl                        => 0,
			subsystem_vendor_id_2_hwtcl               => 0,
			subsystem_device_id_2_hwtcl               => 0,
			max_payload_size_2_hwtcl                  => 256,
			extend_tag_field_2_hwtcl                  => "32",
			completion_timeout_2_hwtcl                => "ABCD",
			enable_completion_timeout_disable_2_hwtcl => 1,
			flr_capability_2_hwtcl                    => 0,
			use_aer_2_hwtcl                           => 0,
			ecrc_check_capable_2_hwtcl                => 0,
			ecrc_gen_capable_2_hwtcl                  => 0,
			dll_active_report_support_2_hwtcl         => 0,
			surprise_down_error_support_2_hwtcl       => 0,
			msi_multi_message_capable_2_hwtcl         => "4",
			msi_64bit_addressing_capable_2_hwtcl      => "true",
			msi_masking_capable_2_hwtcl               => "false",
			msi_support_2_hwtcl                       => "true",
			enable_function_msix_support_2_hwtcl      => 0,
			msix_table_size_2_hwtcl                   => 0,
			msix_table_offset_2_hwtcl                 => "0",
			msix_table_bir_2_hwtcl                    => 0,
			msix_pba_offset_2_hwtcl                   => "0",
			msix_pba_bir_2_hwtcl                      => 0,
			interrupt_pin_2_hwtcl                     => "inta",
			slot_power_scale_2_hwtcl                  => 0,
			slot_power_limit_2_hwtcl                  => 0,
			slot_number_2_hwtcl                       => 0,
			rx_ei_l0s_2_hwtcl                         => 0,
			endpoint_l0_latency_2_hwtcl               => 0,
			endpoint_l1_latency_2_hwtcl               => 0,
			maximum_current_2_hwtcl                   => 0,
			disable_snoop_packet_2_hwtcl              => "false",
			bridge_port_vga_enable_2_hwtcl            => "false",
			bridge_port_ssid_support_2_hwtcl          => "false",
			ssvid_2_hwtcl                             => 0,
			ssid_2_hwtcl                              => 0,
			porttype_func3_hwtcl                      => "Native endpoint",
			bar0_size_mask_3_hwtcl                    => 28,
			bar0_io_space_3_hwtcl                     => "Disabled",
			bar0_64bit_mem_space_3_hwtcl              => "Enabled",
			bar0_prefetchable_3_hwtcl                 => "Enabled",
			bar1_size_mask_3_hwtcl                    => 0,
			bar1_io_space_3_hwtcl                     => "Disabled",
			bar1_prefetchable_3_hwtcl                 => "Disabled",
			bar2_size_mask_3_hwtcl                    => 0,
			bar2_io_space_3_hwtcl                     => "Disabled",
			bar2_64bit_mem_space_3_hwtcl              => "Disabled",
			bar2_prefetchable_3_hwtcl                 => "Disabled",
			bar3_size_mask_3_hwtcl                    => 0,
			bar3_io_space_3_hwtcl                     => "Disabled",
			bar3_prefetchable_3_hwtcl                 => "Disabled",
			bar4_size_mask_3_hwtcl                    => 0,
			bar4_io_space_3_hwtcl                     => "Disabled",
			bar4_64bit_mem_space_3_hwtcl              => "Disabled",
			bar4_prefetchable_3_hwtcl                 => "Disabled",
			bar5_size_mask_3_hwtcl                    => 0,
			bar5_io_space_3_hwtcl                     => "Disabled",
			bar5_prefetchable_3_hwtcl                 => "Disabled",
			expansion_base_address_register_3_hwtcl   => 0,
			vendor_id_3_hwtcl                         => 0,
			device_id_3_hwtcl                         => 1,
			revision_id_3_hwtcl                       => 1,
			class_code_3_hwtcl                        => 0,
			subsystem_vendor_id_3_hwtcl               => 0,
			subsystem_device_id_3_hwtcl               => 0,
			max_payload_size_3_hwtcl                  => 256,
			extend_tag_field_3_hwtcl                  => "32",
			completion_timeout_3_hwtcl                => "ABCD",
			enable_completion_timeout_disable_3_hwtcl => 1,
			flr_capability_3_hwtcl                    => 0,
			use_aer_3_hwtcl                           => 0,
			ecrc_check_capable_3_hwtcl                => 0,
			ecrc_gen_capable_3_hwtcl                  => 0,
			dll_active_report_support_3_hwtcl         => 0,
			surprise_down_error_support_3_hwtcl       => 0,
			msi_multi_message_capable_3_hwtcl         => "4",
			msi_64bit_addressing_capable_3_hwtcl      => "true",
			msi_masking_capable_3_hwtcl               => "false",
			msi_support_3_hwtcl                       => "true",
			enable_function_msix_support_3_hwtcl      => 0,
			msix_table_size_3_hwtcl                   => 0,
			msix_table_offset_3_hwtcl                 => "0",
			msix_table_bir_3_hwtcl                    => 0,
			msix_pba_offset_3_hwtcl                   => "0",
			msix_pba_bir_3_hwtcl                      => 0,
			interrupt_pin_3_hwtcl                     => "inta",
			slot_power_scale_3_hwtcl                  => 0,
			slot_power_limit_3_hwtcl                  => 0,
			slot_number_3_hwtcl                       => 0,
			rx_ei_l0s_3_hwtcl                         => 0,
			endpoint_l0_latency_3_hwtcl               => 0,
			endpoint_l1_latency_3_hwtcl               => 0,
			maximum_current_3_hwtcl                   => 0,
			disable_snoop_packet_3_hwtcl              => "false",
			bridge_port_vga_enable_3_hwtcl            => "false",
			bridge_port_ssid_support_3_hwtcl          => "false",
			ssvid_3_hwtcl                             => 0,
			ssid_3_hwtcl                              => 0,
			porttype_func4_hwtcl                      => "Native endpoint",
			bar0_size_mask_4_hwtcl                    => 28,
			bar0_io_space_4_hwtcl                     => "Disabled",
			bar0_64bit_mem_space_4_hwtcl              => "Enabled",
			bar0_prefetchable_4_hwtcl                 => "Enabled",
			bar1_size_mask_4_hwtcl                    => 0,
			bar1_io_space_4_hwtcl                     => "Disabled",
			bar1_prefetchable_4_hwtcl                 => "Disabled",
			bar2_size_mask_4_hwtcl                    => 0,
			bar2_io_space_4_hwtcl                     => "Disabled",
			bar2_64bit_mem_space_4_hwtcl              => "Disabled",
			bar2_prefetchable_4_hwtcl                 => "Disabled",
			bar3_size_mask_4_hwtcl                    => 0,
			bar3_io_space_4_hwtcl                     => "Disabled",
			bar3_prefetchable_4_hwtcl                 => "Disabled",
			bar4_size_mask_4_hwtcl                    => 0,
			bar4_io_space_4_hwtcl                     => "Disabled",
			bar4_64bit_mem_space_4_hwtcl              => "Disabled",
			bar4_prefetchable_4_hwtcl                 => "Disabled",
			bar5_size_mask_4_hwtcl                    => 0,
			bar5_io_space_4_hwtcl                     => "Disabled",
			bar5_prefetchable_4_hwtcl                 => "Disabled",
			expansion_base_address_register_4_hwtcl   => 0,
			vendor_id_4_hwtcl                         => 0,
			device_id_4_hwtcl                         => 1,
			revision_id_4_hwtcl                       => 1,
			class_code_4_hwtcl                        => 0,
			subsystem_vendor_id_4_hwtcl               => 0,
			subsystem_device_id_4_hwtcl               => 0,
			max_payload_size_4_hwtcl                  => 256,
			extend_tag_field_4_hwtcl                  => "32",
			completion_timeout_4_hwtcl                => "ABCD",
			enable_completion_timeout_disable_4_hwtcl => 1,
			flr_capability_4_hwtcl                    => 0,
			use_aer_4_hwtcl                           => 0,
			ecrc_check_capable_4_hwtcl                => 0,
			ecrc_gen_capable_4_hwtcl                  => 0,
			dll_active_report_support_4_hwtcl         => 0,
			surprise_down_error_support_4_hwtcl       => 0,
			msi_multi_message_capable_4_hwtcl         => "4",
			msi_64bit_addressing_capable_4_hwtcl      => "true",
			msi_masking_capable_4_hwtcl               => "false",
			msi_support_4_hwtcl                       => "true",
			enable_function_msix_support_4_hwtcl      => 0,
			msix_table_size_4_hwtcl                   => 0,
			msix_table_offset_4_hwtcl                 => "0",
			msix_table_bir_4_hwtcl                    => 0,
			msix_pba_offset_4_hwtcl                   => "0",
			msix_pba_bir_4_hwtcl                      => 0,
			interrupt_pin_4_hwtcl                     => "inta",
			slot_power_scale_4_hwtcl                  => 0,
			slot_power_limit_4_hwtcl                  => 0,
			slot_number_4_hwtcl                       => 0,
			rx_ei_l0s_4_hwtcl                         => 0,
			endpoint_l0_latency_4_hwtcl               => 0,
			endpoint_l1_latency_4_hwtcl               => 0,
			maximum_current_4_hwtcl                   => 0,
			disable_snoop_packet_4_hwtcl              => "false",
			bridge_port_vga_enable_4_hwtcl            => "false",
			bridge_port_ssid_support_4_hwtcl          => "false",
			ssvid_4_hwtcl                             => 0,
			ssid_4_hwtcl                              => 0,
			porttype_func5_hwtcl                      => "Native endpoint",
			bar0_size_mask_5_hwtcl                    => 28,
			bar0_io_space_5_hwtcl                     => "Disabled",
			bar0_64bit_mem_space_5_hwtcl              => "Enabled",
			bar0_prefetchable_5_hwtcl                 => "Enabled",
			bar1_size_mask_5_hwtcl                    => 0,
			bar1_io_space_5_hwtcl                     => "Disabled",
			bar1_prefetchable_5_hwtcl                 => "Disabled",
			bar2_size_mask_5_hwtcl                    => 0,
			bar2_io_space_5_hwtcl                     => "Disabled",
			bar2_64bit_mem_space_5_hwtcl              => "Disabled",
			bar2_prefetchable_5_hwtcl                 => "Disabled",
			bar3_size_mask_5_hwtcl                    => 0,
			bar3_io_space_5_hwtcl                     => "Disabled",
			bar3_prefetchable_5_hwtcl                 => "Disabled",
			bar4_size_mask_5_hwtcl                    => 0,
			bar4_io_space_5_hwtcl                     => "Disabled",
			bar4_64bit_mem_space_5_hwtcl              => "Disabled",
			bar4_prefetchable_5_hwtcl                 => "Disabled",
			bar5_size_mask_5_hwtcl                    => 0,
			bar5_io_space_5_hwtcl                     => "Disabled",
			bar5_prefetchable_5_hwtcl                 => "Disabled",
			expansion_base_address_register_5_hwtcl   => 0,
			vendor_id_5_hwtcl                         => 0,
			device_id_5_hwtcl                         => 1,
			revision_id_5_hwtcl                       => 1,
			class_code_5_hwtcl                        => 0,
			subsystem_vendor_id_5_hwtcl               => 0,
			subsystem_device_id_5_hwtcl               => 0,
			max_payload_size_5_hwtcl                  => 256,
			extend_tag_field_5_hwtcl                  => "32",
			completion_timeout_5_hwtcl                => "ABCD",
			enable_completion_timeout_disable_5_hwtcl => 1,
			flr_capability_5_hwtcl                    => 0,
			use_aer_5_hwtcl                           => 0,
			ecrc_check_capable_5_hwtcl                => 0,
			ecrc_gen_capable_5_hwtcl                  => 0,
			dll_active_report_support_5_hwtcl         => 0,
			surprise_down_error_support_5_hwtcl       => 0,
			msi_multi_message_capable_5_hwtcl         => "4",
			msi_64bit_addressing_capable_5_hwtcl      => "true",
			msi_masking_capable_5_hwtcl               => "false",
			msi_support_5_hwtcl                       => "true",
			enable_function_msix_support_5_hwtcl      => 0,
			msix_table_size_5_hwtcl                   => 0,
			msix_table_offset_5_hwtcl                 => "0",
			msix_table_bir_5_hwtcl                    => 0,
			msix_pba_offset_5_hwtcl                   => "0",
			msix_pba_bir_5_hwtcl                      => 0,
			interrupt_pin_5_hwtcl                     => "inta",
			slot_power_scale_5_hwtcl                  => 0,
			slot_power_limit_5_hwtcl                  => 0,
			slot_number_5_hwtcl                       => 0,
			rx_ei_l0s_5_hwtcl                         => 0,
			endpoint_l0_latency_5_hwtcl               => 0,
			endpoint_l1_latency_5_hwtcl               => 0,
			maximum_current_5_hwtcl                   => 0,
			disable_snoop_packet_5_hwtcl              => "false",
			bridge_port_vga_enable_5_hwtcl            => "false",
			bridge_port_ssid_support_5_hwtcl          => "false",
			ssvid_5_hwtcl                             => 0,
			ssid_5_hwtcl                              => 0,
			porttype_func6_hwtcl                      => "Native endpoint",
			bar0_size_mask_6_hwtcl                    => 28,
			bar0_io_space_6_hwtcl                     => "Disabled",
			bar0_64bit_mem_space_6_hwtcl              => "Enabled",
			bar0_prefetchable_6_hwtcl                 => "Enabled",
			bar1_size_mask_6_hwtcl                    => 0,
			bar1_io_space_6_hwtcl                     => "Disabled",
			bar1_prefetchable_6_hwtcl                 => "Disabled",
			bar2_size_mask_6_hwtcl                    => 0,
			bar2_io_space_6_hwtcl                     => "Disabled",
			bar2_64bit_mem_space_6_hwtcl              => "Disabled",
			bar2_prefetchable_6_hwtcl                 => "Disabled",
			bar3_size_mask_6_hwtcl                    => 0,
			bar3_io_space_6_hwtcl                     => "Disabled",
			bar3_prefetchable_6_hwtcl                 => "Disabled",
			bar4_size_mask_6_hwtcl                    => 0,
			bar4_io_space_6_hwtcl                     => "Disabled",
			bar4_64bit_mem_space_6_hwtcl              => "Disabled",
			bar4_prefetchable_6_hwtcl                 => "Disabled",
			bar5_size_mask_6_hwtcl                    => 0,
			bar5_io_space_6_hwtcl                     => "Disabled",
			bar5_prefetchable_6_hwtcl                 => "Disabled",
			expansion_base_address_register_6_hwtcl   => 0,
			vendor_id_6_hwtcl                         => 0,
			device_id_6_hwtcl                         => 1,
			revision_id_6_hwtcl                       => 1,
			class_code_6_hwtcl                        => 0,
			subsystem_vendor_id_6_hwtcl               => 0,
			subsystem_device_id_6_hwtcl               => 0,
			max_payload_size_6_hwtcl                  => 256,
			extend_tag_field_6_hwtcl                  => "32",
			completion_timeout_6_hwtcl                => "ABCD",
			enable_completion_timeout_disable_6_hwtcl => 1,
			flr_capability_6_hwtcl                    => 0,
			use_aer_6_hwtcl                           => 0,
			ecrc_check_capable_6_hwtcl                => 0,
			ecrc_gen_capable_6_hwtcl                  => 0,
			dll_active_report_support_6_hwtcl         => 0,
			surprise_down_error_support_6_hwtcl       => 0,
			msi_multi_message_capable_6_hwtcl         => "4",
			msi_64bit_addressing_capable_6_hwtcl      => "true",
			msi_masking_capable_6_hwtcl               => "false",
			msi_support_6_hwtcl                       => "true",
			enable_function_msix_support_6_hwtcl      => 0,
			msix_table_size_6_hwtcl                   => 0,
			msix_table_offset_6_hwtcl                 => "0",
			msix_table_bir_6_hwtcl                    => 0,
			msix_pba_offset_6_hwtcl                   => "0",
			msix_pba_bir_6_hwtcl                      => 0,
			interrupt_pin_6_hwtcl                     => "inta",
			slot_power_scale_6_hwtcl                  => 0,
			slot_power_limit_6_hwtcl                  => 0,
			slot_number_6_hwtcl                       => 0,
			rx_ei_l0s_6_hwtcl                         => 0,
			endpoint_l0_latency_6_hwtcl               => 0,
			endpoint_l1_latency_6_hwtcl               => 0,
			maximum_current_6_hwtcl                   => 0,
			disable_snoop_packet_6_hwtcl              => "false",
			bridge_port_vga_enable_6_hwtcl            => "false",
			bridge_port_ssid_support_6_hwtcl          => "false",
			ssvid_6_hwtcl                             => 0,
			ssid_6_hwtcl                              => 0,
			porttype_func7_hwtcl                      => "Native endpoint",
			bar0_size_mask_7_hwtcl                    => 28,
			bar0_io_space_7_hwtcl                     => "Disabled",
			bar0_64bit_mem_space_7_hwtcl              => "Enabled",
			bar0_prefetchable_7_hwtcl                 => "Enabled",
			bar1_size_mask_7_hwtcl                    => 0,
			bar1_io_space_7_hwtcl                     => "Disabled",
			bar1_prefetchable_7_hwtcl                 => "Disabled",
			bar2_size_mask_7_hwtcl                    => 0,
			bar2_io_space_7_hwtcl                     => "Disabled",
			bar2_64bit_mem_space_7_hwtcl              => "Disabled",
			bar2_prefetchable_7_hwtcl                 => "Disabled",
			bar3_size_mask_7_hwtcl                    => 0,
			bar3_io_space_7_hwtcl                     => "Disabled",
			bar3_prefetchable_7_hwtcl                 => "Disabled",
			bar4_size_mask_7_hwtcl                    => 0,
			bar4_io_space_7_hwtcl                     => "Disabled",
			bar4_64bit_mem_space_7_hwtcl              => "Disabled",
			bar4_prefetchable_7_hwtcl                 => "Disabled",
			bar5_size_mask_7_hwtcl                    => 0,
			bar5_io_space_7_hwtcl                     => "Disabled",
			bar5_prefetchable_7_hwtcl                 => "Disabled",
			expansion_base_address_register_7_hwtcl   => 0,
			vendor_id_7_hwtcl                         => 0,
			device_id_7_hwtcl                         => 1,
			revision_id_7_hwtcl                       => 1,
			class_code_7_hwtcl                        => 0,
			subsystem_vendor_id_7_hwtcl               => 0,
			subsystem_device_id_7_hwtcl               => 0,
			max_payload_size_7_hwtcl                  => 256,
			extend_tag_field_7_hwtcl                  => "32",
			completion_timeout_7_hwtcl                => "ABCD",
			enable_completion_timeout_disable_7_hwtcl => 1,
			flr_capability_7_hwtcl                    => 0,
			use_aer_7_hwtcl                           => 0,
			ecrc_check_capable_7_hwtcl                => 0,
			ecrc_gen_capable_7_hwtcl                  => 0,
			dll_active_report_support_7_hwtcl         => 0,
			surprise_down_error_support_7_hwtcl       => 0,
			msi_multi_message_capable_7_hwtcl         => "4",
			msi_64bit_addressing_capable_7_hwtcl      => "true",
			msi_masking_capable_7_hwtcl               => "false",
			msi_support_7_hwtcl                       => "true",
			enable_function_msix_support_7_hwtcl      => 0,
			msix_table_size_7_hwtcl                   => 0,
			msix_table_offset_7_hwtcl                 => "0",
			msix_table_bir_7_hwtcl                    => 0,
			msix_pba_offset_7_hwtcl                   => "0",
			msix_pba_bir_7_hwtcl                      => 0,
			interrupt_pin_7_hwtcl                     => "inta",
			slot_power_scale_7_hwtcl                  => 0,
			slot_power_limit_7_hwtcl                  => 0,
			slot_number_7_hwtcl                       => 0,
			rx_ei_l0s_7_hwtcl                         => 0,
			endpoint_l0_latency_7_hwtcl               => 0,
			endpoint_l1_latency_7_hwtcl               => 0,
			maximum_current_7_hwtcl                   => 0,
			disable_snoop_packet_7_hwtcl              => "false",
			bridge_port_vga_enable_7_hwtcl            => "false",
			bridge_port_ssid_support_7_hwtcl          => "false",
			ssvid_7_hwtcl                             => 0,
			ssid_7_hwtcl                              => 0,
			rpre_emph_a_val_hwtcl                     => 11,
			rpre_emph_b_val_hwtcl                     => 0,
			rpre_emph_c_val_hwtcl                     => 22,
			rpre_emph_d_val_hwtcl                     => 12,
			rpre_emph_e_val_hwtcl                     => 21,
			rvod_sel_a_val_hwtcl                      => 50,
			rvod_sel_b_val_hwtcl                      => 34,
			rvod_sel_c_val_hwtcl                      => 50,
			rvod_sel_d_val_hwtcl                      => 50,
			rvod_sel_e_val_hwtcl                      => 9
		)
		port map (
			npor                   => npor,               --               npor.npor
			pin_perst              => pin_perst,          --                   .pin_perst
			test_in                => test_in,            --           hip_ctrl.test_in
			simu_mode_pipe         => simu_mode_pipe,     --                   .simu_mode_pipe
			pld_clk                => pld_clk,            --            pld_clk.clk
			coreclkout             => coreclkout,         --     coreclkout_hip.clk
			refclk                 => refclk,             --             refclk.clk
			rx_in0                 => rx_in0,             --         hip_serial.rx_in0
			rx_in1                 => rx_in1,             --                   .rx_in1
			rx_in2                 => rx_in2,             --                   .rx_in2
			rx_in3                 => rx_in3,             --                   .rx_in3
			tx_out0                => tx_out0,            --                   .tx_out0
			tx_out1                => tx_out1,            --                   .tx_out1
			tx_out2                => tx_out2,            --                   .tx_out2
			tx_out3                => tx_out3,            --                   .tx_out3
			rx_st_valid            => rx_st_valid,        --              rx_st.valid
			rx_st_sop              => rx_st_sop,          --                   .startofpacket
			rx_st_eop              => rx_st_eop,          --                   .endofpacket
			rx_st_ready            => rx_st_ready,        --                   .ready
			rx_st_err              => rx_st_err,          --                   .error
			rx_st_data             => rx_st_data,         --                   .data
			rx_st_bar              => rx_st_bar,          --          rx_bar_be.rx_st_bar
			rx_st_mask             => rx_st_mask,         --                   .rx_st_mask
			tx_st_valid            => tx_st_valid,        --              tx_st.valid
			tx_st_sop              => tx_st_sop,          --                   .startofpacket
			tx_st_eop              => tx_st_eop,          --                   .endofpacket
			tx_st_ready            => tx_st_ready,        --                   .ready
			tx_st_err              => tx_st_err,          --                   .error
			tx_st_data             => tx_st_data,         --                   .data
			tx_fifo_empty          => tx_fifo_empty,      --            tx_fifo.fifo_empty
			tx_cred_datafccp       => tx_cred_datafccp,   --            tx_cred.tx_cred_datafccp
			tx_cred_datafcnp       => tx_cred_datafcnp,   --                   .tx_cred_datafcnp
			tx_cred_datafcp        => tx_cred_datafcp,    --                   .tx_cred_datafcp
			tx_cred_fchipcons      => tx_cred_fchipcons,  --                   .tx_cred_fchipcons
			tx_cred_fcinfinite     => tx_cred_fcinfinite, --                   .tx_cred_fcinfinite
			tx_cred_hdrfccp        => tx_cred_hdrfccp,    --                   .tx_cred_hdrfccp
			tx_cred_hdrfcnp        => tx_cred_hdrfcnp,    --                   .tx_cred_hdrfcnp
			tx_cred_hdrfcp         => tx_cred_hdrfcp,     --                   .tx_cred_hdrfcp
			sim_pipe_pclk_in       => sim_pipe_pclk_in,   --           hip_pipe.sim_pipe_pclk_in
			sim_pipe_rate          => sim_pipe_rate,      --                   .sim_pipe_rate
			sim_ltssmstate         => sim_ltssmstate,     --                   .sim_ltssmstate
			eidleinfersel0         => eidleinfersel0,     --                   .eidleinfersel0
			eidleinfersel1         => eidleinfersel1,     --                   .eidleinfersel1
			eidleinfersel2         => eidleinfersel2,     --                   .eidleinfersel2
			eidleinfersel3         => eidleinfersel3,     --                   .eidleinfersel3
			powerdown0             => powerdown0,         --                   .powerdown0
			powerdown1             => powerdown1,         --                   .powerdown1
			powerdown2             => powerdown2,         --                   .powerdown2
			powerdown3             => powerdown3,         --                   .powerdown3
			rxpolarity0            => rxpolarity0,        --                   .rxpolarity0
			rxpolarity1            => rxpolarity1,        --                   .rxpolarity1
			rxpolarity2            => rxpolarity2,        --                   .rxpolarity2
			rxpolarity3            => rxpolarity3,        --                   .rxpolarity3
			txcompl0               => txcompl0,           --                   .txcompl0
			txcompl1               => txcompl1,           --                   .txcompl1
			txcompl2               => txcompl2,           --                   .txcompl2
			txcompl3               => txcompl3,           --                   .txcompl3
			txdata0                => txdata0,            --                   .txdata0
			txdata1                => txdata1,            --                   .txdata1
			txdata2                => txdata2,            --                   .txdata2
			txdata3                => txdata3,            --                   .txdata3
			txdatak0               => txdatak0,           --                   .txdatak0
			txdatak1               => txdatak1,           --                   .txdatak1
			txdatak2               => txdatak2,           --                   .txdatak2
			txdatak3               => txdatak3,           --                   .txdatak3
			txdetectrx0            => txdetectrx0,        --                   .txdetectrx0
			txdetectrx1            => txdetectrx1,        --                   .txdetectrx1
			txdetectrx2            => txdetectrx2,        --                   .txdetectrx2
			txdetectrx3            => txdetectrx3,        --                   .txdetectrx3
			txelecidle0            => txelecidle0,        --                   .txelecidle0
			txelecidle1            => txelecidle1,        --                   .txelecidle1
			txelecidle2            => txelecidle2,        --                   .txelecidle2
			txelecidle3            => txelecidle3,        --                   .txelecidle3
			txswing0               => txswing0,           --                   .txswing0
			txswing1               => txswing1,           --                   .txswing1
			txswing2               => txswing2,           --                   .txswing2
			txswing3               => txswing3,           --                   .txswing3
			txmargin0              => txmargin0,          --                   .txmargin0
			txmargin1              => txmargin1,          --                   .txmargin1
			txmargin2              => txmargin2,          --                   .txmargin2
			txmargin3              => txmargin3,          --                   .txmargin3
			txdeemph0              => txdeemph0,          --                   .txdeemph0
			txdeemph1              => txdeemph1,          --                   .txdeemph1
			txdeemph2              => txdeemph2,          --                   .txdeemph2
			txdeemph3              => txdeemph3,          --                   .txdeemph3
			phystatus0             => phystatus0,         --                   .phystatus0
			phystatus1             => phystatus1,         --                   .phystatus1
			phystatus2             => phystatus2,         --                   .phystatus2
			phystatus3             => phystatus3,         --                   .phystatus3
			rxdata0                => rxdata0,            --                   .rxdata0
			rxdata1                => rxdata1,            --                   .rxdata1
			rxdata2                => rxdata2,            --                   .rxdata2
			rxdata3                => rxdata3,            --                   .rxdata3
			rxdatak0               => rxdatak0,           --                   .rxdatak0
			rxdatak1               => rxdatak1,           --                   .rxdatak1
			rxdatak2               => rxdatak2,           --                   .rxdatak2
			rxdatak3               => rxdatak3,           --                   .rxdatak3
			rxelecidle0            => rxelecidle0,        --                   .rxelecidle0
			rxelecidle1            => rxelecidle1,        --                   .rxelecidle1
			rxelecidle2            => rxelecidle2,        --                   .rxelecidle2
			rxelecidle3            => rxelecidle3,        --                   .rxelecidle3
			rxstatus0              => rxstatus0,          --                   .rxstatus0
			rxstatus1              => rxstatus1,          --                   .rxstatus1
			rxstatus2              => rxstatus2,          --                   .rxstatus2
			rxstatus3              => rxstatus3,          --                   .rxstatus3
			rxvalid0               => rxvalid0,           --                   .rxvalid0
			rxvalid1               => rxvalid1,           --                   .rxvalid1
			rxvalid2               => rxvalid2,           --                   .rxvalid2
			rxvalid3               => rxvalid3,           --                   .rxvalid3
			reset_status           => reset_status,       --            hip_rst.reset_status
			serdes_pll_locked      => serdes_pll_locked,  --                   .serdes_pll_locked
			pld_clk_inuse          => pld_clk_inuse,      --                   .pld_clk_inuse
			pld_core_ready         => pld_core_ready,     --                   .pld_core_ready
			testin_zero            => testin_zero,        --                   .testin_zero
			lmi_addr               => lmi_addr,           --                lmi.lmi_addr
			lmi_din                => lmi_din,            --                   .lmi_din
			lmi_rden               => lmi_rden,           --                   .lmi_rden
			lmi_wren               => lmi_wren,           --                   .lmi_wren
			lmi_ack                => lmi_ack,            --                   .lmi_ack
			lmi_dout               => lmi_dout,           --                   .lmi_dout
			pm_auxpwr              => pm_auxpwr,          --         power_mngt.pm_auxpwr
			pm_data                => pm_data,            --                   .pm_data
			pme_to_cr              => pme_to_cr,          --                   .pme_to_cr
			pm_event               => pm_event,           --                   .pm_event
			pme_to_sr              => pme_to_sr,          --                   .pme_to_sr
			reconfig_to_xcvr       => reconfig_to_xcvr,   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr     => reconfig_from_xcvr, -- reconfig_from_xcvr.reconfig_from_xcvr
			app_msi_num            => app_msi_num,        --            int_msi.app_msi_num
			app_msi_req            => app_msi_req,        --                   .app_msi_req
			app_msi_tc             => app_msi_tc,         --                   .app_msi_tc
			app_msi_ack            => app_msi_ack,        --                   .app_msi_ack
			app_int_sts_vec        => app_int_sts_vec,    --                   .app_int_sts
			tl_hpg_ctrl_er         => tl_hpg_ctrl_er,     --          config_tl.hpg_ctrler
			tl_cfg_ctl             => tl_cfg_ctl,         --                   .tl_cfg_ctl
			cpl_err                => cpl_err,            --                   .cpl_err
			tl_cfg_add             => tl_cfg_add,         --                   .tl_cfg_add
			tl_cfg_ctl_wr          => tl_cfg_ctl_wr,      --                   .tl_cfg_ctl_wr
			tl_cfg_sts_wr          => tl_cfg_sts_wr,      --                   .tl_cfg_sts_wr
			tl_cfg_sts             => tl_cfg_sts,         --                   .tl_cfg_sts
			cpl_pending            => cpl_pending,        --                   .cpl_pending
			derr_cor_ext_rcv0      => derr_cor_ext_rcv0,  --         hip_status.derr_cor_ext_rcv
			derr_cor_ext_rpl       => derr_cor_ext_rpl,   --                   .derr_cor_ext_rpl
			derr_rpl               => derr_rpl,           --                   .derr_rpl
			dlup_exit              => dlup_exit,          --                   .dlup_exit
			dl_ltssm               => dl_ltssm,           --                   .ltssmstate
			ev128ns                => ev128ns,            --                   .ev128ns
			ev1us                  => ev1us,              --                   .ev1us
			hotrst_exit            => hotrst_exit,        --                   .hotrst_exit
			int_status             => int_status,         --                   .int_status
			l2_exit                => l2_exit,            --                   .l2_exit
			lane_act               => lane_act,           --                   .lane_act
			ko_cpl_spc_header      => ko_cpl_spc_header,  --                   .ko_cpl_spc_header
			ko_cpl_spc_data        => ko_cpl_spc_data,    --                   .ko_cpl_spc_data
			dl_current_speed       => dl_current_speed,   --   hip_currentspeed.currentspeed
			rx_in4                 => '0',                --        (terminated)
			rx_in5                 => '0',                --        (terminated)
			rx_in6                 => '0',                --        (terminated)
			rx_in7                 => '0',                --        (terminated)
			tx_out4                => open,               --        (terminated)
			tx_out5                => open,               --        (terminated)
			tx_out6                => open,               --        (terminated)
			tx_out7                => open,               --        (terminated)
			rx_st_empty            => open,               --        (terminated)
			rx_fifo_empty          => open,               --        (terminated)
			rx_fifo_full           => open,               --        (terminated)
			rx_bar_dec_func_num    => open,               --        (terminated)
			rx_st_be               => open,               --        (terminated)
			tx_st_empty            => '0',                --        (terminated)
			tx_fifo_full           => open,               --        (terminated)
			tx_fifo_rdp            => open,               --        (terminated)
			tx_fifo_wrp            => open,               --        (terminated)
			eidleinfersel4         => open,               --        (terminated)
			eidleinfersel5         => open,               --        (terminated)
			eidleinfersel6         => open,               --        (terminated)
			eidleinfersel7         => open,               --        (terminated)
			powerdown4             => open,               --        (terminated)
			powerdown5             => open,               --        (terminated)
			powerdown6             => open,               --        (terminated)
			powerdown7             => open,               --        (terminated)
			rxpolarity4            => open,               --        (terminated)
			rxpolarity5            => open,               --        (terminated)
			rxpolarity6            => open,               --        (terminated)
			rxpolarity7            => open,               --        (terminated)
			txcompl4               => open,               --        (terminated)
			txcompl5               => open,               --        (terminated)
			txcompl6               => open,               --        (terminated)
			txcompl7               => open,               --        (terminated)
			txdata4                => open,               --        (terminated)
			txdata5                => open,               --        (terminated)
			txdata6                => open,               --        (terminated)
			txdata7                => open,               --        (terminated)
			txdatak4               => open,               --        (terminated)
			txdatak5               => open,               --        (terminated)
			txdatak6               => open,               --        (terminated)
			txdatak7               => open,               --        (terminated)
			txdetectrx4            => open,               --        (terminated)
			txdetectrx5            => open,               --        (terminated)
			txdetectrx6            => open,               --        (terminated)
			txdetectrx7            => open,               --        (terminated)
			txelecidle4            => open,               --        (terminated)
			txelecidle5            => open,               --        (terminated)
			txelecidle6            => open,               --        (terminated)
			txelecidle7            => open,               --        (terminated)
			txswing4               => open,               --        (terminated)
			txswing5               => open,               --        (terminated)
			txswing6               => open,               --        (terminated)
			txswing7               => open,               --        (terminated)
			txmargin4              => open,               --        (terminated)
			txmargin5              => open,               --        (terminated)
			txmargin6              => open,               --        (terminated)
			txmargin7              => open,               --        (terminated)
			txdeemph4              => open,               --        (terminated)
			txdeemph5              => open,               --        (terminated)
			txdeemph6              => open,               --        (terminated)
			txdeemph7              => open,               --        (terminated)
			phystatus4             => '0',                --        (terminated)
			phystatus5             => '0',                --        (terminated)
			phystatus6             => '0',                --        (terminated)
			phystatus7             => '0',                --        (terminated)
			rxdata4                => "00000000",         --        (terminated)
			rxdata5                => "00000000",         --        (terminated)
			rxdata6                => "00000000",         --        (terminated)
			rxdata7                => "00000000",         --        (terminated)
			rxdatak4               => '0',                --        (terminated)
			rxdatak5               => '0',                --        (terminated)
			rxdatak6               => '0',                --        (terminated)
			rxdatak7               => '0',                --        (terminated)
			rxelecidle4            => '0',                --        (terminated)
			rxelecidle5            => '0',                --        (terminated)
			rxelecidle6            => '0',                --        (terminated)
			rxelecidle7            => '0',                --        (terminated)
			rxstatus4              => "000",              --        (terminated)
			rxstatus5              => "000",              --        (terminated)
			rxstatus6              => "000",              --        (terminated)
			rxstatus7              => "000",              --        (terminated)
			rxvalid4               => '0',                --        (terminated)
			rxvalid5               => '0',                --        (terminated)
			rxvalid6               => '0',                --        (terminated)
			rxvalid7               => '0',                --        (terminated)
			sim_pipe_pclk_out      => open,               --        (terminated)
			pm_event_func          => "000",              --        (terminated)
			hip_reconfig_clk       => '0',                --        (terminated)
			hip_reconfig_rst_n     => '0',                --        (terminated)
			hip_reconfig_address   => "0000000000",       --        (terminated)
			hip_reconfig_byte_en   => "00",               --        (terminated)
			hip_reconfig_read      => '0',                --        (terminated)
			hip_reconfig_readdata  => open,               --        (terminated)
			hip_reconfig_write     => '0',                --        (terminated)
			hip_reconfig_writedata => "0000000000000000", --        (terminated)
			ser_shift_load         => '0',                --        (terminated)
			interface_sel          => '0',                --        (terminated)
			app_msi_func           => "000",              --        (terminated)
			serr_out               => open,               --        (terminated)
			aer_msi_num            => "00000",            --        (terminated)
			pex_msi_num            => "00000",            --        (terminated)
			cpl_err_func           => "000"               --        (terminated)
		);

end architecture rtl; -- of pcie
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2019 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_pcie_cv_hip_ast" version="18.1" >
-- Retrieval info: 	<generic name="ACDS_VERSION_HWTCL" value="18.1" />
-- Retrieval info: 	<generic name="INTENDED_DEVICE_FAMILY" value="Cyclone V" />
-- Retrieval info: 	<generic name="pcie_qsys" value="1" />
-- Retrieval info: 	<generic name="altpcie_avmm_hwtcl" value="0" />
-- Retrieval info: 	<generic name="lane_mask_hwtcl" value="x4" />
-- Retrieval info: 	<generic name="gen12_lane_rate_mode_hwtcl" value="Gen1 (2.5 Gbps)" />
-- Retrieval info: 	<generic name="porttype_func_hwtcl" value="Native endpoint" />
-- Retrieval info: 	<generic name="pcie_spec_version_hwtcl" value="2.1" />
-- Retrieval info: 	<generic name="ast_width_hwtcl" value="Avalon-ST 64-bit" />
-- Retrieval info: 	<generic name="rxbuffer_rxreq_hwtcl" value="Low" />
-- Retrieval info: 	<generic name="pll_refclk_freq_hwtcl" value="100 MHz" />
-- Retrieval info: 	<generic name="set_pld_clk_x1_625MHz_hwtcl" value="0" />
-- Retrieval info: 	<generic name="use_rx_st_be_hwtcl" value="0" />
-- Retrieval info: 	<generic name="in_cvp_mode_hwtcl" value="0" />
-- Retrieval info: 	<generic name="hip_reconfig_hwtcl" value="0" />
-- Retrieval info: 	<generic name="num_of_func_hwtcl" value="1" />
-- Retrieval info: 	<generic name="max_payload_size_hwtcl" value="256" />
-- Retrieval info: 	<generic name="extend_tag_field_hwtcl" value="32" />
-- Retrieval info: 	<generic name="completion_timeout_hwtcl" value="ABCD" />
-- Retrieval info: 	<generic name="enable_completion_timeout_disable_hwtcl" value="1" />
-- Retrieval info: 	<generic name="use_aer_hwtcl" value="0" />
-- Retrieval info: 	<generic name="ecrc_check_capable_hwtcl" value="0" />
-- Retrieval info: 	<generic name="ecrc_gen_capable_hwtcl" value="0" />
-- Retrieval info: 	<generic name="use_crc_forwarding_hwtcl" value="0" />
-- Retrieval info: 	<generic name="port_link_number_hwtcl" value="1" />
-- Retrieval info: 	<generic name="slotclkcfg_hwtcl" value="1" />
-- Retrieval info: 	<generic name="enable_slot_register_hwtcl" value="0" />
-- Retrieval info: 	<generic name="slot_power_scale_hwtcl" value="0" />
-- Retrieval info: 	<generic name="slot_power_limit_hwtcl" value="0" />
-- Retrieval info: 	<generic name="slot_number_hwtcl" value="0" />
-- Retrieval info: 	<generic name="endpoint_l0_latency_hwtcl" value="0" />
-- Retrieval info: 	<generic name="endpoint_l1_latency_hwtcl" value="0" />
-- Retrieval info: 	<generic name="vsec_id_hwtcl" value="4466" />
-- Retrieval info: 	<generic name="vsec_rev_hwtcl" value="0" />
-- Retrieval info: 	<generic name="user_id_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar0_type_0_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar0_size_mask_0_hwtcl" value="16" />
-- Retrieval info: 	<generic name="bar1_type_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar1_size_mask_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_type_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_size_mask_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_type_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_size_mask_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_type_0_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar4_size_mask_0_hwtcl" value="16" />
-- Retrieval info: 	<generic name="bar5_type_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_size_mask_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="expansion_base_address_register_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="io_window_addr_width_hwtcl" value="0" />
-- Retrieval info: 	<generic name="prefetchable_mem_window_addr_width_hwtcl" value="0" />
-- Retrieval info: 	<generic name="vendor_id_0_hwtcl" value="4466" />
-- Retrieval info: 	<generic name="device_id_0_hwtcl" value="57347" />
-- Retrieval info: 	<generic name="revision_id_0_hwtcl" value="1" />
-- Retrieval info: 	<generic name="class_code_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_vendor_id_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_device_id_0_hwtcl" value="10337" />
-- Retrieval info: 	<generic name="flr_capability_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="dll_active_report_support_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="surprise_down_error_support_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msi_multi_message_capable_0_hwtcl" value="1" />
-- Retrieval info: 	<generic name="msi_64bit_addressing_capable_0_hwtcl" value="true" />
-- Retrieval info: 	<generic name="msi_masking_capable_0_hwtcl" value="false" />
-- Retrieval info: 	<generic name="msi_support_0_hwtcl" value="true" />
-- Retrieval info: 	<generic name="enable_function_msix_support_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_size_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_offset_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_bir_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_offset_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_bir_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="interrupt_pin_0_hwtcl" value="inta" />
-- Retrieval info: 	<generic name="force_hrc" value="0" />
-- Retrieval info: 	<generic name="force_src" value="0" />
-- Retrieval info: 	<generic name="set_l0s_hwtcl" value="0" />
-- Retrieval info: 	<generic name="serial_sim_hwtcl" value="0" />
-- Retrieval info: 	<generic name="override_rxbuffer_cred_preset" value="0" />
-- Retrieval info: 	<generic name="advanced_default_parameter_override" value="0" />
-- Retrieval info: 	<generic name="override_tbpartner_driver_setting_hwtcl" value="0" />
-- Retrieval info: 	<generic name="enable_rx_buffer_checking_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="disable_link_x2_support_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="device_number_advanced_default_hwtcl" value="0" />
-- Retrieval info: 	<generic name="pipex1_debug_sel_advanced_default_hwtcl" value="disable" />
-- Retrieval info: 	<generic name="pclk_out_sel_advanced_default_hwtcl" value="pclk" />
-- Retrieval info: 	<generic name="no_soft_reset_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="d1_support_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="d2_support_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="d0_pme_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="d1_pme_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="d2_pme_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="d3_hot_pme_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="d3_cold_pme_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="low_priority_vc_advanced_default_hwtcl" value="single_vc" />
-- Retrieval info: 	<generic name="enable_l1_aspm_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="l1_exit_latency_sameclock_advanced_default_hwtcl" value="0" />
-- Retrieval info: 	<generic name="l1_exit_latency_diffclock_advanced_default_hwtcl" value="0" />
-- Retrieval info: 	<generic name="hot_plug_support_advanced_default_hwtcl" value="0" />
-- Retrieval info: 	<generic name="no_command_completed_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="eie_before_nfts_count_advanced_default_hwtcl" value="4" />
-- Retrieval info: 	<generic name="gen2_diffclock_nfts_count_advanced_default_hwtcl" value="255" />
-- Retrieval info: 	<generic name="gen2_sameclock_nfts_count_advanced_default_hwtcl" value="255" />
-- Retrieval info: 	<generic name="deemphasis_enable_advanced_default_hwtcl" value="false" />
-- Retrieval info: 	<generic name="l0_exit_latency_sameclock_advanced_default_hwtcl" value="6" />
-- Retrieval info: 	<generic name="l0_exit_latency_diffclock_advanced_default_hwtcl" value="6" />
-- Retrieval info: 	<generic name="vc0_clk_enable_advanced_default_hwtcl" value="true" />
-- Retrieval info: 	<generic name="register_pipe_signals_advanced_default_hwtcl" value="true" />
-- Retrieval info: 	<generic name="tx_cdc_almost_empty_advanced_default_hwtcl" value="5" />
-- Retrieval info: 	<generic name="rx_l0s_count_idl_advanced_default_hwtcl" value="0" />
-- Retrieval info: 	<generic name="cdc_dummy_insert_limit_advanced_default_hwtcl" value="11" />
-- Retrieval info: 	<generic name="ei_delay_powerdown_count_advanced_default_hwtcl" value="10" />
-- Retrieval info: 	<generic name="skp_os_schedule_count_advanced_default_hwtcl" value="0" />
-- Retrieval info: 	<generic name="fc_init_timer_advanced_default_hwtcl" value="1024" />
-- Retrieval info: 	<generic name="l01_entry_latency_advanced_default_hwtcl" value="31" />
-- Retrieval info: 	<generic name="flow_control_update_count_advanced_default_hwtcl" value="30" />
-- Retrieval info: 	<generic name="flow_control_timeout_count_advanced_default_hwtcl" value="200" />
-- Retrieval info: 	<generic name="retry_buffer_last_active_address_advanced_default_hwtcl" value="255" />
-- Retrieval info: 	<generic name="reserved_debug_advanced_default_hwtcl" value="0" />
-- Retrieval info: 	<generic name="use_tl_cfg_sync_advanced_default_hwtcl" value="1" />
-- Retrieval info: 	<generic name="diffclock_nfts_count_advanced_default_hwtcl" value="255" />
-- Retrieval info: 	<generic name="sameclock_nfts_count_advanced_default_hwtcl" value="255" />
-- Retrieval info: 	<generic name="l2_async_logic_advanced_default_hwtcl" value="disable" />
-- Retrieval info: 	<generic name="rx_cdc_almost_full_advanced_default_hwtcl" value="12" />
-- Retrieval info: 	<generic name="tx_cdc_almost_full_advanced_default_hwtcl" value="11" />
-- Retrieval info: 	<generic name="indicator_advanced_default_hwtcl" value="0" />
-- Retrieval info: 	<generic name="maximum_current_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="disable_snoop_packet_0_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_vga_enable_0_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_ssid_support_0_hwtcl" value="false" />
-- Retrieval info: 	<generic name="ssvid_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="ssid_0_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar0_type_1_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar0_size_mask_1_hwtcl" value="28" />
-- Retrieval info: 	<generic name="bar1_type_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar1_size_mask_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_type_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_size_mask_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_type_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_size_mask_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_type_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_size_mask_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_type_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_size_mask_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="expansion_base_address_register_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="vendor_id_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="device_id_1_hwtcl" value="1" />
-- Retrieval info: 	<generic name="revision_id_1_hwtcl" value="1" />
-- Retrieval info: 	<generic name="class_code_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_vendor_id_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_device_id_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="flr_capability_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="dll_active_report_support_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="surprise_down_error_support_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msi_multi_message_capable_1_hwtcl" value="4" />
-- Retrieval info: 	<generic name="msi_64bit_addressing_capable_1_hwtcl" value="true" />
-- Retrieval info: 	<generic name="msi_masking_capable_1_hwtcl" value="false" />
-- Retrieval info: 	<generic name="msi_support_1_hwtcl" value="true" />
-- Retrieval info: 	<generic name="enable_function_msix_support_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_size_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_offset_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_bir_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_offset_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_bir_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="interrupt_pin_1_hwtcl" value="inta" />
-- Retrieval info: 	<generic name="maximum_current_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="disable_snoop_packet_1_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_vga_enable_1_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_ssid_support_1_hwtcl" value="false" />
-- Retrieval info: 	<generic name="ssvid_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="ssid_1_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar0_type_2_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar0_size_mask_2_hwtcl" value="28" />
-- Retrieval info: 	<generic name="bar1_type_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar1_size_mask_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_type_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_size_mask_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_type_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_size_mask_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_type_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_size_mask_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_type_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_size_mask_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="expansion_base_address_register_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="vendor_id_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="device_id_2_hwtcl" value="1" />
-- Retrieval info: 	<generic name="revision_id_2_hwtcl" value="1" />
-- Retrieval info: 	<generic name="class_code_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_vendor_id_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_device_id_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="flr_capability_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="dll_active_report_support_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="surprise_down_error_support_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msi_multi_message_capable_2_hwtcl" value="4" />
-- Retrieval info: 	<generic name="msi_64bit_addressing_capable_2_hwtcl" value="true" />
-- Retrieval info: 	<generic name="msi_masking_capable_2_hwtcl" value="false" />
-- Retrieval info: 	<generic name="msi_support_2_hwtcl" value="true" />
-- Retrieval info: 	<generic name="enable_function_msix_support_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_size_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_offset_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_bir_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_offset_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_bir_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="interrupt_pin_2_hwtcl" value="inta" />
-- Retrieval info: 	<generic name="maximum_current_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="disable_snoop_packet_2_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_vga_enable_2_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_ssid_support_2_hwtcl" value="false" />
-- Retrieval info: 	<generic name="ssvid_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="ssid_2_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar0_type_3_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar0_size_mask_3_hwtcl" value="28" />
-- Retrieval info: 	<generic name="bar1_type_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar1_size_mask_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_type_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_size_mask_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_type_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_size_mask_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_type_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_size_mask_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_type_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_size_mask_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="expansion_base_address_register_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="vendor_id_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="device_id_3_hwtcl" value="1" />
-- Retrieval info: 	<generic name="revision_id_3_hwtcl" value="1" />
-- Retrieval info: 	<generic name="class_code_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_vendor_id_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_device_id_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="flr_capability_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="dll_active_report_support_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="surprise_down_error_support_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msi_multi_message_capable_3_hwtcl" value="4" />
-- Retrieval info: 	<generic name="msi_64bit_addressing_capable_3_hwtcl" value="true" />
-- Retrieval info: 	<generic name="msi_masking_capable_3_hwtcl" value="false" />
-- Retrieval info: 	<generic name="msi_support_3_hwtcl" value="true" />
-- Retrieval info: 	<generic name="enable_function_msix_support_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_size_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_offset_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_bir_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_offset_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_bir_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="interrupt_pin_3_hwtcl" value="inta" />
-- Retrieval info: 	<generic name="maximum_current_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="disable_snoop_packet_3_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_vga_enable_3_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_ssid_support_3_hwtcl" value="false" />
-- Retrieval info: 	<generic name="ssvid_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="ssid_3_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar0_type_4_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar0_size_mask_4_hwtcl" value="28" />
-- Retrieval info: 	<generic name="bar1_type_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar1_size_mask_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_type_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_size_mask_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_type_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_size_mask_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_type_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_size_mask_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_type_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_size_mask_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="expansion_base_address_register_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="vendor_id_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="device_id_4_hwtcl" value="1" />
-- Retrieval info: 	<generic name="revision_id_4_hwtcl" value="1" />
-- Retrieval info: 	<generic name="class_code_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_vendor_id_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_device_id_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="flr_capability_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="dll_active_report_support_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="surprise_down_error_support_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msi_multi_message_capable_4_hwtcl" value="4" />
-- Retrieval info: 	<generic name="msi_64bit_addressing_capable_4_hwtcl" value="true" />
-- Retrieval info: 	<generic name="msi_masking_capable_4_hwtcl" value="false" />
-- Retrieval info: 	<generic name="msi_support_4_hwtcl" value="true" />
-- Retrieval info: 	<generic name="enable_function_msix_support_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_size_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_offset_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_bir_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_offset_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_bir_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="interrupt_pin_4_hwtcl" value="inta" />
-- Retrieval info: 	<generic name="maximum_current_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="disable_snoop_packet_4_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_vga_enable_4_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_ssid_support_4_hwtcl" value="false" />
-- Retrieval info: 	<generic name="ssvid_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="ssid_4_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar0_type_5_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar0_size_mask_5_hwtcl" value="28" />
-- Retrieval info: 	<generic name="bar1_type_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar1_size_mask_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_type_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_size_mask_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_type_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_size_mask_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_type_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_size_mask_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_type_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_size_mask_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="expansion_base_address_register_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="vendor_id_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="device_id_5_hwtcl" value="1" />
-- Retrieval info: 	<generic name="revision_id_5_hwtcl" value="1" />
-- Retrieval info: 	<generic name="class_code_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_vendor_id_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_device_id_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="flr_capability_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="dll_active_report_support_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="surprise_down_error_support_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msi_multi_message_capable_5_hwtcl" value="4" />
-- Retrieval info: 	<generic name="msi_64bit_addressing_capable_5_hwtcl" value="true" />
-- Retrieval info: 	<generic name="msi_masking_capable_5_hwtcl" value="false" />
-- Retrieval info: 	<generic name="msi_support_5_hwtcl" value="true" />
-- Retrieval info: 	<generic name="enable_function_msix_support_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_size_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_offset_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_bir_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_offset_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_bir_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="interrupt_pin_5_hwtcl" value="inta" />
-- Retrieval info: 	<generic name="maximum_current_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="disable_snoop_packet_5_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_vga_enable_5_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_ssid_support_5_hwtcl" value="false" />
-- Retrieval info: 	<generic name="ssvid_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="ssid_5_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar0_type_6_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar0_size_mask_6_hwtcl" value="28" />
-- Retrieval info: 	<generic name="bar1_type_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar1_size_mask_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_type_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_size_mask_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_type_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_size_mask_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_type_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_size_mask_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_type_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_size_mask_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="expansion_base_address_register_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="vendor_id_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="device_id_6_hwtcl" value="1" />
-- Retrieval info: 	<generic name="revision_id_6_hwtcl" value="1" />
-- Retrieval info: 	<generic name="class_code_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_vendor_id_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_device_id_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="flr_capability_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="dll_active_report_support_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="surprise_down_error_support_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msi_multi_message_capable_6_hwtcl" value="4" />
-- Retrieval info: 	<generic name="msi_64bit_addressing_capable_6_hwtcl" value="true" />
-- Retrieval info: 	<generic name="msi_masking_capable_6_hwtcl" value="false" />
-- Retrieval info: 	<generic name="msi_support_6_hwtcl" value="true" />
-- Retrieval info: 	<generic name="enable_function_msix_support_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_size_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_offset_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_bir_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_offset_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_bir_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="interrupt_pin_6_hwtcl" value="inta" />
-- Retrieval info: 	<generic name="maximum_current_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="disable_snoop_packet_6_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_vga_enable_6_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_ssid_support_6_hwtcl" value="false" />
-- Retrieval info: 	<generic name="ssvid_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="ssid_6_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar0_type_7_hwtcl" value="1" />
-- Retrieval info: 	<generic name="bar0_size_mask_7_hwtcl" value="28" />
-- Retrieval info: 	<generic name="bar1_type_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar1_size_mask_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_type_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar2_size_mask_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_type_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar3_size_mask_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_type_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar4_size_mask_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_type_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="bar5_size_mask_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="expansion_base_address_register_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="vendor_id_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="device_id_7_hwtcl" value="1" />
-- Retrieval info: 	<generic name="revision_id_7_hwtcl" value="1" />
-- Retrieval info: 	<generic name="class_code_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_vendor_id_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="subsystem_device_id_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="flr_capability_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="dll_active_report_support_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="surprise_down_error_support_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msi_multi_message_capable_7_hwtcl" value="4" />
-- Retrieval info: 	<generic name="msi_64bit_addressing_capable_7_hwtcl" value="true" />
-- Retrieval info: 	<generic name="msi_masking_capable_7_hwtcl" value="false" />
-- Retrieval info: 	<generic name="msi_support_7_hwtcl" value="true" />
-- Retrieval info: 	<generic name="enable_function_msix_support_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_size_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_offset_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_table_bir_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_offset_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="msix_pba_bir_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="interrupt_pin_7_hwtcl" value="inta" />
-- Retrieval info: 	<generic name="maximum_current_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="disable_snoop_packet_7_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_vga_enable_7_hwtcl" value="false" />
-- Retrieval info: 	<generic name="bridge_port_ssid_support_7_hwtcl" value="false" />
-- Retrieval info: 	<generic name="ssvid_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="ssid_7_hwtcl" value="0" />
-- Retrieval info: 	<generic name="rpre_emph_a_val_hwtcl" value="11" />
-- Retrieval info: 	<generic name="rpre_emph_b_val_hwtcl" value="0" />
-- Retrieval info: 	<generic name="rpre_emph_c_val_hwtcl" value="22" />
-- Retrieval info: 	<generic name="rpre_emph_d_val_hwtcl" value="12" />
-- Retrieval info: 	<generic name="rpre_emph_e_val_hwtcl" value="21" />
-- Retrieval info: 	<generic name="rvod_sel_a_val_hwtcl" value="50" />
-- Retrieval info: 	<generic name="rvod_sel_b_val_hwtcl" value="34" />
-- Retrieval info: 	<generic name="rvod_sel_c_val_hwtcl" value="50" />
-- Retrieval info: 	<generic name="rvod_sel_d_val_hwtcl" value="50" />
-- Retrieval info: 	<generic name="rvod_sel_e_val_hwtcl" value="9" />
-- Retrieval info: </instance>
-- IPFS_FILES : pcie.vho
-- RELATED_FILES: pcie.vhd, altpcie_cv_hip_ast_hwtcl.v, altpcie_rs_serdes.v, altpcie_rs_hip.v, altpcie_av_hip_128bit_atom.v, altpcie_av_hip_ast_hwtcl.v, altera_xcvr_functions.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, av_xcvr_emsip_adapter.sv, av_xcvr_pipe_native_hip.sv
