// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OAzxmfAIk1RXMi50ABqSM6IUvCYg2uzNq36Es1CeZAYt5d5mbq69YSDv/0I6KjDQ
s8gob8jWTGVUp4UG9GhmHIBxagxyDVH4Xfqu2ZMD9hOXsLyTOOd7HnlJQlQRQdjG
OLaLJWpyWGfNuy6aH/d/rLLQBbroU/hUGAualyLj3nE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 174144)
df9fP7zsDxj62RhZhGwJHm10LGguGA0NkiKQmXgW/G2A5E0yIPha1QaJQSVnRM2H
mdd7UbjbJODoyishCsSUNV7wMH6RqqWACMS+3HKWz8e24myElA00D0pGud6xDj0g
wYy0AzIQEcagbnK787ru0n/3g7w1l7yMIi/D3R2hAhlU+Sk5kg7e95UfBzSDzcZm
XWhoMTxdPJ01qeDn4u3Vs+QfoUbVLIcEiktWUokfGQvHYppHbMH4VwJzvrJ6synZ
2K5BwqdVADCz+dlcNfdM51RNav7vFIzz28kppjfKR6M2hX5RdCpTvYIkwzDG9SUr
REE07u6l7ZHGWmndaQkEBwwqIklm2j4pPNj7g1iih8RBsKimf36Xxm6UtaGFtbSy
4uB/FU1i0E5xWJP8I/4f5eflw3CQOkBPcnFojMmB5bBtiBmc0aCXuf8jy9W/fXki
Ezqyu/kpsZLugZ6R128XJMoTDVMF0pxW/CPJfQkZJrEiJG9QHdqultJQmY1VDvKC
U6KjlI4Tb2cDI7UoJyvTcqUesfbEa7UQTJ3qPvj1xcik1hEUIvbE71Z3AvakSUnF
F3FTH7Cs7dzx5gv0IZgUHIKaz6BA8JCtZMxD7AcasOstBfw7rEhoPlgOoGQTSDDg
EYg6uVaZfSPgJc3NOsOCYwKtzOcm95KVjpNplDeoIyYdXjmCEJJiQ3mu+hYACA0A
I2Pe5f6ONEk4OSabjpzxcPX+XBtc7NiOpkq/32b/SBSBZBMHSiCT79lCQZnGMwod
98pTAldvj7R9CJUIeADW4fCJhKI+Nhsk6wyTxM8ZJok3Y+LoDHI60bg+XR3T3OBs
J9aCtMdKkn8+X8lfFTQeZucb2YzwFbytA0PZuMGC7cTnNDbrC3hJcBDbCMJN3zRr
rSDy7oZSasTY082q2tKtAGtlrZO2XGBQLVFPDuxAAHj3nxvjrqBhPtZ4WoA7Fch3
AhrsepM67+SUmkmFceZt/19HhGMkHN5oczr8x8B6b4LBevlIKR9pWmtQYIZACHK2
fzD3TTf28QF5y2nOR2yLwKxTdNuKeMLu0OrfSxLLqgUc4P9GE5To5NE/ZWuJvMfE
gbTo7hElumYSTiQ8fgK6HiBqlQHhubGzfG+oPt4rAezduD7f4nH6wp7HCWCQx73c
xl2EEALLGjPx1+an6CUORl9WIgETK+VXZLI/RVpOPcRFF+UofH4Vp2WQGX0jpFqr
0E9UJU4mFchAMIoQdpByYPNnp4Ovrqrvt6rr3/HhsXruAL9vnFYgAnn1JxYMmTst
mzXYrwQ34t5wUwWp3E802NlcJ8P8L2UycEI0xYfe3oLeYbQwbQ2lpDX3t3LGoJqH
7MiJVlAVcxJcF6zXK2qghlRiRSiNcSE0ShR8cXJgnXIDl1KsY41VVuLDG6yfWv+E
AgUbiMycfo0C3dOJrkaXJ5dqyXq8nIfwQb+S5xb7d1Y3fb12+YVeRJ5VGr0Ybjf8
vUg8lIyhEI8azmeXy7/LD9khZrX/5ecyGdGVI/m+IGymGrLFXw+bN//urQ9kP578
TrQIVQVtK3H1JCfLOGWSXb8hQ1EgHYchZQH7JturK4DYtc9DtA2mC60OBDIdyDAg
TTsrSUG3Eu1AbHWoogiOK4W386JoN7sURSpHVcGHl4AI2d72nYHZicdus6uSEbBk
4xFX9eD5ebt4jKvi3vLu90YGt2et+4necCNBysO/u7/eumC7pASIER7eSMZCBiUm
ZTjs+WNPIl6+UN+gJ+nyM1DX+F2u/MUvdFD39wpso1GvlXgxMU4ULFEahgVJ9HxU
kHO2PcW0Ov+L0uAz5PBI9ywWyKkIWC/XLA8LPsTjDlKDqFeSqjWyc5GIIgB7d/Bj
fv8reYydGTpP3/nklFMLrjF12209pBwf7GE8ee7SQrLQp4ujGEY7xi+wGuVzwcDl
58ac51/XLCC9fMIMtvVvd3wuePrBthwc5z8cPeXQKgBR3Sd3UAfB/EvEjOsb+h2M
YQMFHc95owe54YcHDLvmUV1LsqRop2OrffAhYBZi/BK08pX5bFD5F7336/WrDrCI
hF+qt2xN7f0ydA9AWoxHHZss1uyj8CoVmIF8/DAKlGUO0XnG7H8PokDCeQz+N8DY
o2LA9fAklUx7KlL8hJteo1TsRaEPzO+ZTj7+7QUXjgpSZGdirTOjSP98y4eC5K4J
hbI4wJ2JknT4u38df4O+lCTEpDsHQMOmnr1FrYbPXDBYQQvAmhCu3n58N+M4fZE5
k0jihQUD3EBFU7qAzy9SxGqR8A5wrNfWUFzCgGQzlHmulqIdrI7mOUTVgextHIdE
OZx02OMjCJ7lgBUCevT5jXDFw6XfzoDmh9vj8jjL6CUK2LqEAvLIrozhmUVuun1H
LKD675Yuc3q2++wZc0LlAdN74GuzXRl7K4gSyBqmDTIs+QwcvjxzKhDlw3EN4q/P
D7t3gsrboDFKrlANeY4eUpt58GVSI2BMTitWr/z9AO6V5IdsVn7dhOgAOAT2nKGg
BJ0RY+RjIzwihnvAEYCNOooSziFbr0k+iHKpoxy4aieWExAl+pSWZSWN6D/IKP9T
Dx12UhPkxmbbSUOB9K60bM3nAK4RVXZ7zD7gxTxbAzscUh6vpaDOoGVuckUYP4lT
rIOZz4zscEKlUaQg8conkv44W2WbyfTFVpTzL5ALlUlQMKi9lNUrVZ45E/P2AzbS
Wefc+eD1WGWNu09rLEpN5Ld7Ci93mdC8SqS/MioJ4Us/R1U2vs34ICaUpcTFWDsC
RtJErCvaXgXtkWEiZI9ByNq1kCGGVXNB5qLEMNyCnkIKi3oCBqeRU6vzq8ooC11W
IHIKGTcUo6i/yrYi9a0yNbrf0jfKN00fkmTiWW0zkfwHLNGMvN07eOaeMS5wsOaj
kQOa0D21F6mja9zt4L21h0Cc4yUwm27RGzPErjLPrwmboc5635+cnJp7L1jc8MBv
yO0TjI699Erog3Hqrub3g2QUwVEOaS7qgpa1opwjDuuoIMm0VqN3/XSwPUmAhKUp
wr1Cg+pX6FbYbk0jk/fqtVIXjvxTuTOB/Otn/NRfTi3Kh/SypbTs9LtaYOfwqsd5
hS0+S4TqwFkcJl1pqsW3t22ISdqhzd6B86+eBkK/Ya048V7+A3VeRTDNZAtRZ71p
sQqEuAjLu5R8tRzweF4ehzo7ZPJkR8UpDKPwAaV3g8XH8170IoDu2SDgwGjp7tuz
2iDs7Sb2hU+wcLO+ui77nKE0/bsh6qxMduxH5RVylp0UntLtxU2SRkH9gRLr0J8C
sw+RrvtaIi/lPI3fmqRzI6l8XpjdUgJiKE/3tHSDk2jRMkc+z8xXvMZXIqS+evRz
HHBmtI1LJ33v+ReZt4sy8wlKpafG0JexRUT1I3pfiZO5RCXzfDj1fBpO9tA0X0wK
u+A0YZJfVai9QRUi5977T14agRtaJdELKrqJXtIP2AfemBUXzc6EvaK0dq4yqFSj
RVRzJv0Qp3z+5JAjVPTiT1s9O4N8ygRuN2Qy8wJSxV6BiZDKG0aq2NO0DwsjS/Br
mht0U+UDU4LBxxZlzL2LqX2XTNCepRW/lbkLAk9Z5KhJJ6OnhkCgOSd+7IQOYwrc
36CgV66CFc+GOiUL8d7NpPpq7cnDdxoSVXTlC5BLkaQ31tiLXyDnMp6vaOrwsaUR
r8n7QDv+GAWVlsgMHX+JmpVzEhbjJenX8UNZF8gTDK6U8s/3BmeDo3r6pEOYb6I9
p0kgEN4FysR7jv9scNuCaPZXMBMfm9Vnt14R5hUZG3yXGmvT/dx6c/DHDd7vJ7Km
N8uIOSMZ/+h3lJwydeiYUfmuHfpWbej6M1cWFJ6Hz6vSH4rjm4/eFVjFfzd6+cDc
ZITsz22m6+undlof7HBVbfFuyzfc7jaT3KSygE3URoz9VFluO2pp7K52Q1tmlEF4
7FEiA+0pPCAKWexgMnkS/FWfJM5IMQe8z5bjvxzJDWnNqbZS3TENDkw5PCdxUtCm
QnyXx9zzWwOElL9UUDBRkrSuO7XGm85OFTSLbTYVLg0rkSbPTBEZHjkDw+/m4L7O
Ld0N27L94IXP0WOON34DGr4kfQbBy4/pbphT75OexHzElrJMw5kfxv/+ZZCGIw+W
NheKsaUvDGai0NQVGKzL8ZQhx7Q+LzICfmEahM9SsdO+lhmhaRDgUZotXGucYsrA
b6LHXMJJzUjLxrITehVammoPcQ0mkAxVx/yNTupWLXDPWzOJuxxaXDbCj3uDkviq
c+ciX2SyySYyg+ywGqrHbIUZQvTv9B5PMPJo1pxLpECDXxI9zi5CqNqiZI7EvQNG
poiHAOpn8ghqzyyCDguuN2z8e84iIRGVqpumW9LR81llgLkT0y3omxqpVnbx3A0b
y3CC8/VGBX6p9CBSYPLg+bjVrwVjrj5Pp8RjIKxDQwFVRlAX6DO2b5t3hjN6gBAg
SuFYRD+ebUCWAW6MRjwzvXGd19+o+k4zYDc0bVnvVoEhymM2tbCVZUJnMikEMe7d
WmkVg6jwOpANRTEU9SBQB6PVwtTDk9codzpDh5NhCRcx2WIivvCGFG5SQaEmkTjo
3htr2K9PsBNAnnnwzKGfrsQifp4rM9ifv/f5yy0FlO+WPsU3XZQ360acmP6NrzDu
9pyDXzBJZy/seM3+fpxOm2Vf/8FC1Ia0PBVfS2SJJFDRckRTDzLj6sfxnYjouZul
1olFLCP0/aMnCKWaZWQcEXOFxdj9FWBEZoSKoAdVSS9RzvlIkDwOQHQDRy11vfuB
FneSFuGQHkKcTDL51tmQrbOFojE2vWteXeN+XTxx5vh3lB9Q/H5FL4gd4HMj6WqF
p3H77HJqV4atc5hMwjrACTyPan3iteK5jZ36HUAjaKWqItNXWIHDnnDw6QNlooDm
4EeKCXP+HUEeMrTTFTvIUScHftk+s/Re0wvJEztGMnvI10o4eFQyY/lo0Ur4ITn3
J+eJE+1U8gKLfAt5X/0BODwczXtP3pDX8xKFSTpRJEKPLps+4i2S768nYKJwrM9/
bqba717i85vo6J7np+pNCpPDyro7N0lDy35vxasFeW3UFoJUxFY86AG6iV7Z44/P
NeV3O/fG9o+QHPim2hBOvS3qB/049dBo05kOjgpoFEh5T4GKpzcqaYeMq2aCEFKk
cnIB5vyPA0jVpDpRUkN9s27jvnaXXOa/QJkq1rI+BLDLestL7mIuod8DDNJXJr3x
FlNnU+CImumJ1fquT0y3kAd7v9LdqY/SF0mH1AyQulM4D4yIg6MIx1/EPWTpvEj1
ctiKq8ReKas0KNyI7soBRW1pKP0+Krjdq4MysoBuPpeXLGC4dFzyLE6/Izizptj3
D9cAQK0aCPFsg+kOD0pwc/WlE5TzYNG7BLRMOPQ8rlDHyE/4H0w/rAeE5zQKi7ne
odeC1Na9Rb9Rn2qutuZ6igvplU4K0ID+0G+JPgnDHLnAStwhBRe9zXLHn1WKtvjr
4v4/BoAMpy0hyRB66IzyxVeMoW/P2b5bt2e0RY+2c0ZQG2yrOr2hMNMf2JTdwKY1
hap/qu3s1Ww18TjnMIONb2X8LColjdXZ0weB/ytY3bPprGUkVC3y71EVqLx1WTng
Sn+Rvw22kkrH09Zm79Ti/vEjHt3sqJbWtgMWLskMIdSH6po0kyqh8H4u1Lq5soX9
yth4BnRG79cz0dJtozAAQ2qhICUWAdhAaSGTQoNcB1uTYXEO1K++67lZ9JDLL/HO
QIJZkUlvQtkg7YYW2d/dazfXCthJs1dFvP8/ssrtuhOrv4U8Mp1dWSU37jhm8Por
t+G5YdXnp1QFy8530cp/0PN2qfb6WEE9RX9ndjqV/kr59L1PIas2oKpS/6ezmEh4
JE71J5U+a6JLOSM6HLwl34CnL7vDW0fsSjZxOosmAU4AepsNaX7yJRB7N7mTh6gF
HAqPxR2eFxTesd9qvnZPWZBtxmdElgpQhJyjo6dFSWwmXCkkPBCswn0IVkyPiWHZ
+lvX8wIICxl4QisOydAeCxOue+BUT4v1miXQok0dJ+ir+PEiJGJ1J0XRdRCjvOvL
j3oYFKa3YCf+/Cu4FOEcxYgxnrfg+0/xQKpKzbnanVUZfvv/cYTVttDLmlZg682H
BI5cpmwmQi6JNVRARQkx2q6K+O284TvMcT2SPCAZ7YOmC2vvcHqjdims+48nDi1J
bXtUOUI/3wt6jYR+/KiWw94pcBdPuaTec48g6cG83E2rhceibFidWVnRYMPI68zE
1mMMqETD+eXjIxA32XMJJHPVMy+SdWClR1VHj9gzV5jV8GctB2puMihEWMeetnmt
0W8aMb1IgYaiDQiHflStO+wqMopt7reEaJQoqw90EQpdzchZ1in7j9nCfe4/gmbY
q80jg2OMAxYa7WyQeSWkUBPFW5zBvDM6GId0jpW05xp4fzbA6+zcTh23klJSOCdC
zhZUC/VqzWhEBCc9tebN7QA7Z4V6ztORr6w5f6xbizQX4DI8d/ASPp7D3Nb3ixxs
SZTuxQpN2cT/rNnZKuBjh8PcdnRKdb1eX1NpE/QvEhlSNb+UHigO5WZKFi8iIAan
CFfqYElvMiLc8t6ir6GDkxrEJANY05OxAger3a+DVQ9tnc9DlyS5pAxfdPuj/sVT
TxjaRnt8L4JYHhNMJBFl1sJlRJrF/ohkOQdy5eKYEJv3RPT3NAwuMFTGE7VjZzRP
cRtMQtB+xTki0ODQ56xzAXOXbBbE/kpUGYqEGvSO7R3empmeI7qTEhHJIeHUhb7F
91SfnJiklBYU/rRYJlHE9kw1Rvxa1AUUeLzsOokojaCv9JPaPbINBn0D96Ixe8xj
6ar6tzi0QH7YlpY56hiPiLA9dUYoIYuYXF80Q53/A7nsSMqIqQBeZ/nm5slXrLoE
5owSMN0uX4BzER4W4Nqu1ajQoboIwIhYWa5Z/bkeHIi18p87G7aeqymfWZd7NtfI
PZKFbeOzU4bPHsHDBzykr0bwLrthuRhZS/i4ZObUWWUWCJG8xeZvcuTFBvbzwFqv
qczuppL1BHN32UMfFxg4FOBcOiAPsroj6aiqdHlv2lMkepMWZmpw1ui9KX2/WRmi
stSwwdlX52z8j26ZfXe+bzPsMWavsJEFs3VLPwyxQiJqKqRigZXWflVTo7Pipovd
WHIxR+ebQ62KrA0/XdLzQSC40vUltcBVIYtdXwR4r2xLf+fhIuyVSBghJV/fiwXd
nK+D/C1i1pUOyYMRwVL3lYQmN8RFEBdhZNYJic+efsPFvAVJoBJO679T3vfxdyDX
0ff5QcQyQdPkBh306AgMM0Mkm+iTBQIRUlEwMHu9wJIYHDmIuKc4/mrYguk6UuN4
TxI8a+DTEMH3AO2AK9byl7qU+qlzzquOiWVph0RKm7JmIF74DGsSXf3AiqTnA8Qm
ILWJGaEcbV7lmwRmM9xKxccB+qethD7kEr5qXUHOkzkj38TkjTgKlgbrjeK5kEVO
zKEtjKV1Yp6ieqxl0VtQLFp+XaENqRMPq/zGNmiIwQkF0K7aABKoA8gWicBsz/zH
xHDOIPKn4M/8bge4AD+u0EXNWcoUK3w10j5tlv6+Y/1YmaO7b8dwn8Lqy7/1AQFQ
5MoEUz1WT7tFudZvodt9PPGt0v6epzz2eEcPXM4EbtqZ2OoiIHcK+t36R0wd6q4k
7wJ+DUSp6mzz9nyhH9QdpYzXYYcKR2CdOecwmI2CI4PEbHOFN7I8yKnD9yoJLVY0
r2gBJeW3lFgJ7blsJLjGCS1XJq8nLt6OdUiOFaCQ1WCX74PuBqnhLdrIAIPF3Z9C
oJiM7hMmCRn16GHQxLrG8DSAAde/Xbz+Yyh6ykzuji5GOATufLOgwgrwajtiE3BL
8Z5TL7ZMrKDUxKrR6zJ9mQkLMN9f5LwQeBotYVUEyG2n7A9Vag0wHMwhKgrw3Bst
UxqjFHLnr/EBgOxa6MFH74+hi6SfyyBLie67EaD50ai01mq6e6PqJoRw5bS8z/ME
8C0Po/di7H0WaW2fNMO4yGEvCYJptS1ZCz5N07bRgk2SKPkdcYCV8wqrVr9jszLY
JMSpl0wwKf3p2Yi1lmATWHUOsUTia+oFIv6FIj4JJ8HnQJ3GSt9wn64Oz3W5gZk3
hIuYA/WX4nkjGZhwyeSO3wFL6X2H+27zGCdn9k1zkrjvHpEDEKD54MrKHNESEp7X
BOS+M8WVNfx2lp2OCCqAQisrGXQ1SDKO1M4KABRVqf2KGwF7vqdtyQL31WM6Pr74
BV7yuYVJPpAAAHqyb9FJ7OSZW03AW89u0UwYJuNJeGyxOaBy9VGRstkz+o0UDxlH
9E89Cc+gJ1e4LbSpjOdZO9hllMQtGeE5xHBOZtQ1irIjKEcQ/Dlwk3sTruT6C1dB
5ZQt0p3DWXF3cccKCahFWggE/+PaPa7vrOfSaYUrW2KwvIHP6aXtaJyWr62XNLTc
2sJ9u/6FW3sX1Q6KMXYwjd7/bbECo5EmoxFITZcthBIcikAXNJxYhFK9pBEbqz4C
VRFBb6hsSQwMP6MSE1QfLxaFHW2Mdiny77MBwV2OVmhk9R1g0O4WzrQM8KvUinOQ
4auVYrUtZu3JLDe7CQuJX0AyJbo5KGFog/cb0slq5W2zbrMSjBnMhHl1+K3rXnzO
haHMLmNASnNEk40v7csZ3ZwzaIWOYUSnqiZxFGRI13LEWDcwem090wJSCI1O5lHO
hxbQspZM1PKZITZWzyB8xSi2/0zNCb/q/SC2AawuB5Yg5xIleARRfQKpKKWYz2RB
klaQqpznMd7Z0qafbUP3DXDO0MPFbM8eQtYuqAj6zbo1fhgnbt4Hpm0BkdsHjx+V
3Qg4NWL0RBAu4uup0+d0QSCQdJeLL6Ew0RhEB2jBV++LVSQazfm0ThzPKU4KUgur
7WPOIsHJymkKh/0Fdhm0hr17ZM00uxWYKVmubC6b7t6fjdPqCndP9B0U4ovMA3Sb
ADJfVsmhDY4VHvQOAnVD9Bq9yK2qWtxdqFEQ1E3xNX+4Rxx1w9zSGUrXoD7uk4B4
30IoQUJnpLPhm1zd3wvzV9g4tPMffiWobuKGQGokyui0wKOTttZHrfLEc9xsXEkI
AkZSQYPvUzkhm7qQL4gKLxkdOATrsSPLic6JI4LjvlST6Puedxj7GeFb/HMQQIsO
OvdiS+SkuiuyeSYOjOW5W/9NFqX/KBcJ07sezVZgJ0q6sxDS07PNhXquDyTNSpXm
8CeAZF7OfilsTCd59X8D1YBTWFDxolZWA0OQRdn0geh1jHEmkCrIbqkSTXtAARW3
JqJyOZiU6Xv80iCTAciAM3Vz6dHWePuVIeqOPiVm7PaT8VhgSWTdXXT3AIlBgYpX
iapGyN648vdw67vJ8K56SRRLfEUKPhcccJlbtD8JS4YW4g4YoVzAgmwL4M5D/C+R
bpn0r5KfwZzVljDNMgFdOowJs8MJHl09dDcN2tDYli3X5qw2qbcgcN9q+8JwPt+K
bGVpIoLW0fWvJV3sz+Pn25UR/CeyRwgLg8zEEsi9lVTVC1u9i+EIknrY652vpeyI
4rM3ihi/g+fqzrvuC7oHRROB9ExNkB4CkAi9Qe5v1cu4ewwHUWTxBGVdeWGS8qjH
fDfZZLqnQLjlwrkNMHt1eQQ3fD9T4hlDbd1hNjV/hC2ok8YY2ZMiyGyW3i0EZlrq
pMCuqCdrOOOZ9CLOANpjAYIrE21U4N9rtYqRqDoIdennwO/s+1F5FM9xIitS4DAy
Blyim9y8piB4S9b8XXJg7e0yGjaBPUSAJywW9V0MNWnnwyZA9/PePXey9XGK8+Gl
kGBDHHTjd32Eg6xWCHZSzfyQDZF3AcM0sh2UqjuPNvpCNLseBXC4H361lyBZDlFe
r/8yb/REMMTpmLMLFCWcxb+H6zcp6D+9OYrukwHh7zGv1oo2Fio0yDMdECYX33dR
WWLyYKf44S6DHCGHIqFQO4cQJC7atimHi39vSEbuz0Z3LTZcF+xPGblN2JiNfTnQ
ncLAVCPLy4AUWzVm2QkqUr7FdntEk54hoKivlKUZNfNo97BpL7Kp/sOtOArfFeVB
FwPVxW9I0ns41yDlPtcCgulkAyVbrHlSPMEgV802GyZWP8iHQoL3BMfGnktulBij
GnFndRbPp6ummMZUBpDQwh281+RnyLjWPyAACQkAUr7eKrVSqxaFyZ2gORPEXFTc
L+oI807mY4LecC3Tg9rPfIADFmiMv0VsJn4+7vTe8O6BcWk+DujDJ0/kgyhdNzpq
UWa9r5Uqmz8prZVc3YyIDyvMwL9fP2ESF90sv/XYrO/lnmdnFwnkJ8YhrXiOlZPd
bJNQLv2bmHhmlMtymS42KhZopkI1BFoTCDEFbVwn8wT5jvJFb8q4Ep5EKheY06Wf
jV+N8nfhlvhRsHmiXFv7axnSxGB30mJwEMqkoKd5nfmdkm9LEzTbcETIBflIyBcR
GL31+qJSrwZqRlRA/g038LCzWpKASiZprac2mFP/AQPWC0Vx8goibBIq7CWzNU03
rrxvnPKZZhmT/q8XbGRB8OL6T7BAWRcKPrvzPtrrk1iqr9V85Ps+wN6OkEzwr9lS
i+99OVXfTC1WFchWcEKos9OKeM6Be0Q2aTU8vTPN6QSdvE3UdnT0LwY6jOuUwBfR
iBoN1E/cSjBclWe5h0rI6GJLRPamLlqG7omIt8KFhKLB6ULVayb6a22BOyLfW3DG
TCShrkpVinvo2BZbBtRNPAUxTg1h7GrTw/6ln3h4X7Z6MtN+yejgHFhKBVZ1LgmH
m9plYyvprnvAgvfT2Vwj3Z54wJmRCmklxmze6O5jhe5jsdLpHI/Miz8KryXr6hnu
3Capp3LNGzhx34+YTadVnq2JKbE0GQ/UASEdDRuFJtyHYsPKLfCBgEHFhQel6VaI
T0xOvwhLwu5i6HyxZMrFAjof4gxnX4SQDzovmnGM5qySFDFibtfZESg5z2NmA5Co
lu6ZM0wsKmjSQLtWD1zTm2puXDH7bH1iNe+hi3Zk/KdReZLIg2eGA0yQuFE0lXtV
IiG95q6pQ+YfurJSu1KBVM+fXhTMwGnV0O/AQpp1T6gMTNUUQTD3/PK8X6qAPwz+
jT3PASVnwpE75FhimJlKe6eBg38+b9g3vkO8lS2kyWetHM6WEi/o3db3OrfawDeB
L13VfluezJg1LDlFmWx9XS4XlpshrdbyXQSDPeYfdZ4zGEXMpdSp0kOVukkiGOFh
hI2jvEonoAsalE0+40ddRJf4KuDyr24GbudeyWkXRfUk3Vz74CgIaLjm7s/18h1T
D2OKy2lnf/ODqio+5tqcydCypdZpvzELcbygWbc/PKIlmS04JNcAnErJp9vRJnAN
/7BpzpwsRNvZcvsOflKEssel+oA2d5J4NC1kEBBm1qQ5/8YwRq48s1IWREBZDCxR
q4WhQg0yT6pxB6SoeG8PYXSKikEsiDoKTXYs2FF9vtl2XuHVAgbnMyZdUL/ZwW0M
M6F3m0FNCCpBXbOsVAC3hiDTWccFtgFuzXMaqfyrlJgn1jBr4sbg37kO4zT7i5bQ
iZ3Ryj4sr1kMsQgosD1DNjVBtL1LFsU4VZyw+POsmJy9EVr/EWFRNOQwwLPvzNI1
wXMvrmWziaj7jHZeGZb3SkM/hAB72laPdotaIArRb8QnD8C+BLEuUEU3USrEj9DX
6PEtgP62hc6klSfptdP3nAG7ZmwKZGvLsKi3WE0qvPqnHji83p46fTHN8bayU8w6
Sjc3YdbYdUrZFaGYKUr4jHynT2Ltglk5AH8WX0PLOvSHLLHuajgafwXBVVjstMgP
h64Vc8wyAjAP60pePbz3PuFHwfT0mmwJozAaOF5KbW0bX16+PsQYhMTfPIEVUao9
5oPyIPtDnZ0YBAsH+7A33pEuHx+VnN6EG2GF/UT/H+BYzFxRam2c8VaY7VH9Pd/V
MuMJedWqnyoGfNFiTZ4cgW8n4kH5cRPmQEv8XJbFLgimy9IzoX5YufXldA8I7VbN
4Mh0Iw6Hp3BAWDP4fw2LIVXP7mPkPkDHBFJUooi89fATySr79CTogT8KRD01rxbC
JMbtKSTBTMsJxbkm5VY6Pb7HFLafdoeBu4EJ2rw4deczyyugPYvFa0n0jnpg85y4
QmG9i+gIOUIn/IxnmQGUX5F/z3pZ4BzQAqnbWFmt5M2dbz9sM6gBlH6zTAMl8Cc3
cnpRDxTYFFnBVfMdYj2AQJCFjT9e8s8WdfmuMO1EOpRBHpc6W7gMFl2ZePb48nSv
h8kl07bQeXSzbhrw3l92MJAAsSbYiYIVgI15lNiJUa0AbH+pgLA0HsdyQ6yd7b90
+FVFN7tdMufj62iKhE1vN1isgauYQJftBri5gSpnyamS31PkdId1JRb+3r58XwOq
VpJ/o2/VTR3/y+taX6GCxsJN82ZQ+b/PBKyyrhB6DufFxRjTU1VX0illnNS0tVKM
5nnxbMvLGiBAETfx5DMIPa1bFZ38v/kdzdy7KQ2sGTlH0hzEOSLaBlGtiYQ8HcUO
L5J7r+J/NzX55paxOyowqlDL4GIbTElp4XYpHipCpOgHhOsgrYtI2l1TP/B3k8DB
nG73YKoHaHitC0B6XiknAvhZaQDFUl46hqwuL0tQvWZph8uWV0xOSskntfiINWVL
UB2BS3piOoOfNXnBvS5Gr1xz3dhteLOKiLMVgd7fMCnHaf2DJkCBDL3HvLYzsTWJ
mFbtMTfLpmqAr7lKjhgxcp3L2HDtug535E7vedWcmFSTuTn8FM+HsIfQRxK3vPXE
9Kv0KUPsoMgcM/Ddo5G+rcc7YUAxITliPodbO1eymKEKy8JlqSdFeAdMBtRQiQi2
jbTdv30ghFJBZrQEUfDg/zZ7GPOufyxBhMVV/eMjXquXNn3qsyUSx+oowc7kE0mR
VpC839McN2YJ7voxqRu0rSqjZhGre43Q8MdEXikAdu2xXdUeGhTV9mZsdi417/kR
j0BwhCqDaQ5BCnmgMgHYHdQEFF6qlt5Ez2/cs8Mcy81oOYEeRaXda8GaGTWG1rFQ
3F/raybZPgd0Fl6GLbWrM3hpBI8cD39l7h6WDhaKu3gycmGVTgi+XaIS7ZDSzT7O
NyaMxJu3nce7JSvFauc4rPMXkMSkOzecXZ1ih/0uV/c1qdhWsMir4uKSQ7awu0Z2
Q34KoHtx6pCPm9g+9n9/rsqOuOvkFLttvUvZvyqUklylLUPgtMwvkmCPzeRjcBXd
pBnchLAD7TM1/j7KK6n8XLxVzLyIjWY1TQ6YXx/jxAMMru1zztk087lnaUVCqhdL
nzcuK8dXp7f7a67+ARf6+bHVZF7rL7T8qcY/wrp5+OtTXwPH0kxxYR7U3C31CV6F
kk8b57afreRyOxDjNovPaPyr2jJIfiCYwis4q+Yk2Y/ZdEog3L/HCqwVBR7T05CK
F+ndWqeodiEakITCps7XZw6VS3/IV9VacSv01EBF5/huj91xyIpTFH0a5k6DpTT7
e0gWEtv0eRjB/2WoJzElb2PxFkN6hETrzsX92Oi1O69Qk8s0FnrtW8R/suLdQAco
eV2GI93+JlsjZie59i+u2xPv8RYiJzxTAJVuYNydSmtV2q45YlrwJHLJOJPbAOIe
k4/26abXagxjeKY6Lb1xl+Ndyp2uN5RQ4nuEP3acuoXiG5PxUmAN4hZd1+a59L30
hJC0d2KS0PA66pWxdsMpem+5e5SwPp9Z6gsb/PnTX3bxnC2QbiA8qJfFDjldhd9v
y3zCq5hUzMZasTrxbW31PpbqIsmmVhDx8qTb4RhiSVhQoDVuhRninExsNWyVdAQ3
il5+VnzpKduvJ+7KulGaczFi3jXoo9zexKD8tpscinfLWnmn6gkJlMM5MOWipAab
jAgt9y5mrpDcd4d7vxJU7n15mMt7Rn5ZZ+qypmn8Z+dycN+OlLq6Z7fX8EIuDOkY
7i6UvPL6Sr4FLjOsOjrPHFh9XFw2P9jiPYqjJe4lpPEzQNiTXQ5jPSH+iwwENFmf
X5ZFozU15Gn9GBXoFUHCJSiXiiwVwbM8rfyatb4RezgZgqOX4ZOA5eD4eD4FUSaq
PwgPUGAiqtipYjhb63qSssYR+BzSqC01h7nlaSqdIY2OODNAahIhwPaUwHd1j9v5
LE0qMdBMbBGS02GhJCllD3v4c2m875DlB3Gg3gIDOmRSNdOy8np8O8Xv4BorzPQV
xnOvB7jLunVbW1lGylBZVKmAqiOqpNNiz2NThK8E65LMVin9zX5IEDpok22UzdLs
b1luSrM/kCHPJOArHnXOfwW2YJh52/oLoIw0BYTWHos5MzZVdRX90aM1NlQvkRq1
tukru/N04gAukmlUc4DCCPXXa6UppL2FViVWKnbfd/I5q710FyJnh1NcEdupCUtd
TS5mPKxBxwnJ0ESwTXNlr4UJ4YZBBbWRPzNeTzAnBWorv0o6weNOyz4OpTPgJysv
pczXF4tF0N03Mh89MWZu9nocr67xBmtB2+tZfyH6fLcwFUSochEgLphrrRcqVHiK
GYlLSHeyqVWHdd720QAvz0gHGsP7kO/u5AjEoePk7mn9m+pJ9dnZC1ryDtQCojm9
hd0LRpeTarxfI6Sb6TB4RZDLCo/wZkVKGaorKLvljzRkSRYjBIIgJaAf3iTn8DRo
2XWctON5QKfekGnpt942KALi39PittkD86wvAXiahFEzab6Z4z7+vbSQA7n7cRj6
c5yjX+qQ33CfmDX1Q3g3bIEA1HIoESZJ4xob7zrTjGdNC7k2QPanKlpBjIQTExEO
IGp68L8ZkxcJe8KIi0DOuMZn3FBR9C9RVNnobO7monmq1KzZis0YoZmXc2DI44/6
kRznZB42QSYkzYLuGDIN5U3NS41A7dp7XQqzQW4hb5jJRHs0o+y1YzdkzCjVIYap
yUoGEGE685STxktDAtnH2qaCi+FKIj1BbNHZy2cAQgORbk5AGsMUs2/5uEdBHNeK
G/TYVv7A+UZbk+Ch9hrgIxydk5E//A8/R/dMOvDQ5gNQ7FI9lAC1lL6DaS+adrRg
37h7eM5kY9ojouevis7KPAv0ThZQypF1e7W4IIvJxHdk3nbI2nbm3bt7T8DttSqW
4nQ+p9g/Pscnee7jZpOPW4pIKF/NqHlBC0/8X+9ihai9gDtQmVodkWfvtNeXg9Y0
Gpw8OwESfu1cG4GOS//+G+11MxoAcLujmRqNRfOPC8ZdPYXWl07OrN7LbvODBPQD
/Pqq/3200RK43Zt+UMJCO6l8QaCdGgx2bfzlbOP+7aqiSY+i5dBRYXEss98An7VO
r7GLiRm5ViQmc3o7g19Rbl9+5e1ZtY5OA2js4BWMcofKkci4HrAsQT7oC7j2egWS
oejoTGVBnRe4hGRZW4826vBctJ4PqDFxh9V2TofqFgfNj+9ItKqRS8EX1M6Dk7dF
RisB3v2mt/AFx4AFCotBLfjJe3EdcYYTKAySyjutbPg3h8ceVhch6nN1Z4qnu+RI
Z5uJ68k3os8qi5l3q14C0lZvbs10gfRCPK5PH+2tFOrYv0crfJY9wFsc9B4nzJk/
yDVSqpQAj4isjDG85Bz6PcgKoz4mM3f0kLKksvyhio+8p8oeRPrpYCLGQBqDDr/u
qtIXMQ97D8knSUBzTtrkqUd2GRN03focL5NbghMBwotmrUVETFx9vtNyJwfq0w9Q
C+J4YzS5tyjC/s8ceVT8LLJ2RHHVYucwJU5bylfvJhxJzu/5Hz9JxI6GzyFL2qh3
EhVQ2EXT4CKc31CZ3O/4YL0dgqSWznIUUTpQJBUpgfl3eMoKjQK2VGA60zBH/vk7
iqKslCIHShPzbYs+sdCO9Ir35t0wsl9JgzopKOyIxDU8XtaOtrna+/77YG8uJSdR
99IUc9jFk6Ybrd1JUMg245bGWLipGj/elkueQ5Rr0STUkOtwtn3pd2LIR80b7Qmb
KLW2zcHPuinl+pppcKTqhmxRqXvQ4g/AVjUjXy6HMMALuFVjWKNIG94F3GHM9nUX
ps29DZSq6mFGeyim5Ex3dlXOxvpwa23SH/45p6GvxTcQObGGqxVw4cQ9FAoAaXyC
O5Ijk5AgJwu3ApBp4WylyddR3VB+iivzvCyQXu4XnSdLQ0hrNTvzTpC7mkvfHeQc
66+7U/Ws0aBCHL1gvpKynrXZbclTaAKIoS6KSKrXvgQz/SX/QWezgzlDJ71H5ZFJ
37qssVbN8lJxM/mYRfcddrck1jbbJ1c1wjWkhcQsFcUmRwAA2C2+qmcn9ZQqmaO2
leIoDPQAGoabPuCKqvdsM67vljlOe8P4VXI/OcTVbLWys+oFndiRQ2E9HF5coqMQ
WV8HouUMBM4ovWDnHc6VtR36AFDLGTLvzhlNoNzF5Ei0Wj2D5VczTnuxZF40jndy
ZJFvzoN1tAlRLI71BicBDfY+wAcebivC3Qp1ebJkErPsqe8TLUbEkU/qCwOH9xYo
Gv4Kd8c8VO4XvF/7DUMhxcsRMghZ4BzXMUZDfjOoUP4ahkp6Wdtk3HXooImPGMYw
iOJR0dBzYgJNa9RCTIy5+kmtBALp0Wuv+OpTL2y66W02QCig6MUe8zp9rVRNoFts
EGU/ytl2ZKm7USa3UEwKxzOrTGsbvzsjQBxm8uDW0xHtx0ifRmhzRdz5aKQe5Nr7
u5dttJu/YCLNAHQi45VM/tHIF4mTKLvXLSQYWzeKI2bYFKMXlJ4AD9n2YuRhrJdd
f//yHFKJXa48JXg8WmY03OrO7cdXDr13IPY7K8MT9VOajxPTWc3zU5wXBChVWd1u
bX3eXw3USG+fcJPwRn8Xa6l9e6OSiRn49JlWmNOrfpCSriVkwzC6JW/G2xmUdczP
FToV2KEldE1PoxKDVhGQBN4KnfsMSD9AMPg2n+3ovJwfpxfOtCP9Ul3Vd1p45cf0
jn6Z03TOlvOqeskAqWLbz4z6VY9Ea2++baXdmebjDaDvxul8BixoM/5syGKoVf5D
zb0iK0aEFQKWkkpyvIK0+x8d8t42M51gfm5mLjwSfihvr2THco/KKC/9PCBuwoee
/WMGXkQX+efmxITaHrwlaVVzNve90TjhIfgZD/M+wU5OFx0LL1T9/AjiA4xu2Bel
cDUFGJcxh447BKe0U+5VZfNfqfA/z/QL1UjGCmKRATL9XqnKWqoY3Cul64S57Ik7
blaZCCf0tJf7eMmqtfiS6ViJP6IQ615EuRbgGhyU/j+6u9ekWbef4dSu/hr44mt4
eAwa+JPpanQoVXC0MPI7GL+KPXg1xWr862zjXe/cUPgcnukqrybcR/KTivfJlZZ5
SrHe9wvXblTjeS85Kq3T73f+ZlddScd3C+k9Y4CO1WTwsagyXpt2VYuAxKBb3t2Q
KlsZ+Ea2KTfzND3RdjZVT4i5695uJWQ58SBG8Dxcm8QEwGnGEWuEPagHMK/E35Gk
Sbj/GrNa9voZNEkv5KE5oEhTzjwoOLtcebWPItT3bZbpHYsqG1PY54Ky8R/Ah9dE
v4EMVF/eGqS4Mfwn1MCgPsCVH78On5/+Sm68ebtX/NMnk8N4YP+Q2I/Bp2pCL1Pa
SjWkXpaqnW1r3LGM7ZnkIAgmVcE/KY49kio5yyTVJbqdWkKYsewbKtCHRXxQwkR3
HTmX44ZdqcUDWDGqan1/b5kuhtn4Oxjn34WGx7BcQjudTHk6Nn7dgl1W1smZDGOa
aSrQPAG1TJcc3zxNN5K1u0SPxeOUdWl8sLzkVXcjFaazT0ZQSH1El+UkRHN6Hgey
x2pXi14tiyJKgYs1kpnid4wEiFBnmBeaOIbkkdghK85XQlHCZKcR8A77ZKgop7Vi
9bc0gYfvES1QTUyvqcTVli1ryPdTySKUsz/kmE9xIUFhZAK++xmNHYqtXb/tqy7z
07oDAttCK5urRIJ5BrHtMPA40xvDDg6n3/KFH+3v45+k2Ev1YYurChGg2slCz6uM
d8m3ptLXYRH/ht0dI3E/8hAd6/TUIt+GGWNdDp8uyULf7MzBCa6cCDQ2EJf3kDcU
QajyDjb8XO5C4g1YoOBJi9wiBoKN5R5IyKI3j3Zil71hG2sp8jW6QDq8qkOGv424
d2A78RGIy1oSr4K0Rf0IE2NVJiAvCPlLHpSxKnGDyIKEWWYPPv6Q0ebrW7l0TjFs
k0lVl/0r4JhVXXvYIaPJVYOoZoFuKAPXlYrEEyqwxrZlJbQ+zYPSyARyp7zGHsUG
3jijRRiRwjYxLPC+oS97nvBJoyTtMJRHgRGcJCI9OQD7V72+oeM+FX8c/nAmzu8H
1hVnCfI69gRnLdOD99H9rGpWuAwoKELTP4Uyw3Ycd8VgIaYi05qVHxEsBa7etaKq
ca8Km4qbwBvFTyvAGH4p0qVSJbc4MlBUeJLtfs9oqxaXV+Ql+6C60xerqEdJ/nNn
QO4lkdZPMvI6LP8WwO9OEsvooMWq7J6hPR+lcDtCjbVC2edMiq3xJPlvihaPNEz9
66p4dYGAZxRIqQxOhXJ7Joh9jwvKZ5BimbmfOhuvwe1PXx84AjHAg4Oh3AEtlOrY
855y/FXJEdySdTQTYFXxIk6u/gQCIkLJH2xjZbiE0DEsaSMSlFqW1QYBsvBZUKiF
q11sZkb7hqehzmc97LcHnoO49hMwZ0cFZiGH5zbDsjfdlAGZ1YV0WLpOdK2tKCfj
Did/t1mU8Sjx2gMqUtQBJdRHaMMQ57xsqBVEuAjMYJLQggafTNJF/Q9Aqux4J06m
EeNjwrBDlM7iQzxuZ74Hm+KQ8KFvMfiAl8MODsAAFzHeHurxSOaundkS/4VtzjFd
DSUvxvgqNXwRIoNOieFNtTHoHI0flqPzKZNvD6gPRVPhplA8TjnTAgQvBnKeq+jg
eYMzMjsILWEWgSjwYDsZP/AA6FyybOpGRaot7rTh0SlU9vhWbwSxLQ1jOsOKjKeU
JLpyE22J8AzO3znii+wtd5IK+2XBIcwwDjXzYdRy7NBhGL7B8VpEnz4KptJxlXeh
TVyQVivvaMHQRbwaA0XvJDF57qX2+PdqPWkB6lAWIWu9Gta3wYA0Z7izk9Vrcd6r
O48nMD7zpHmmHxb4S1UU2IIdfbCkATY5vB/KSBPO7ywyNAWWvlHeaTBXP/0OKbHs
2NdUgkR1dQw260prVREqB36AqXobTif84jFARkW7TiaUXmWSxt3eMYvnw85FcfPq
mKOIXV+nYYGkJ5e9Hwla0k2oXYxkHfZbN1jBCTBfmb06+yz7hGj4E2sOyg+HHMwQ
e+V5KyDSoKlrkmo3jJniosbZo4l1qMMgvUAPQm3iJcz98UfNlL/v2yvI4wcu6qm3
ahAxGDkueHLFO+rUlBoXb5pBfLEVo3B5s1Lv1cEijlpHyd62NZvjXk1UyJBgjEbR
xHIkl8M5BUeSDURA990STInw/u6ttjeY/FfpiNlSqoA38732TQvcy6AVEnAQAMt1
N//4JUBpjavKlQ0NkfQmgCpFHffhu8vTl3yivHHt5TsNMFvyLyJezFvn0DcI+Y/J
VhBl3gTn1BOFiOX6akvMo9iqkXgbabvinGvahNtz4A299Nga8odv7adZT1VkDYQJ
xR3jzhsJhrCzUZNSytwKgBaiFuLFK5DZ1AWxfcOUs3+8MONyz6BdMc7wtI8B2mez
WYWZ2AktmhjeDhQoViWFyNzwp5koVAvO5LmkrNIRQ/uItxaanLZF0jhaaqZX3Qn1
w2h17y18C5KSKE6rulWv5ysdX52Gp7FSmBMaez0Lj1XRXSncEbXozim9K3C6s+1w
b1uKZA4tqXg1KJuPkyg8iip/s9udwZkSYaw6c6SOdognCaXFPpHFL40fr0vLFPji
oqYzrjEf2xpPossalnMFLe7Jd6E0THRKK1f4eeMoObFxu3PalbUrFfubrB6IIghw
ALfGzrArRkyYpF8R4cLBGHFuusQ0FkBSYRJvXxzFF0vCMxtEswGaoOHFpUPb4p/u
D6S+PF9/jBEAIrad3yJrZWRL14O3FP48yS1PTeqG6QW2R+RcRNUjwkizcu+7cvcF
sbj2ercz7IasB3PmOB3dhxqygppbyvc9/U/Pv+Iu3fwgK+A/i3vcli28G8rsznx/
2MxEjKQQFsZIh92xFJLR9/3IHqq1MuOkIrU4xITSXZwrxXshkwHXFgP24IaYHY1l
8W9CpGdEkxAGSnKqiS9Io9ynRHgaGe2XVw2sJsn3iRH9/7PPAf4hlJkhYBIA0Jwl
smG9SLrTzmqzZ8jSqQJeQkLMZAQo1fhuoWhwFQHA9Dcy2gvhkoDq+tPI5Cm/tY83
fajE0DFYAPF2e4EWzcYJMdEdCluGaFmYN1E1LS0LSGCBm1u4d6dvZGZgomhNn5GM
FwcPNoxuBQQX/R2SLMXX0yCmh9+FtEWVrCfP8GCuZN6ATqiBv2U+NxDsg+6HOHZZ
CRfl9VsVbjdk2mCXBF/02DdUWiBRrPrdX1OnuwwvYNiRWr0nvhBHpjS5vwKOCweZ
8ucVp1ZlMq8gWeixuFxwIwKDCP3eA5Rlm39QhqI9r6luFTiz2NB6lATEm9/kilza
ANDyMr0qqHwePSigPZfqvM4IR6I7LbpHD9Sgt3Q6iAH6ti5F9lf73RHH0KtEofGh
TKO1Bpbn02gO7Jx87h7pSUgPwnsi59x1GOGQqfU4QLc3F2nwVKKLkbxQfFCCdfdA
RT08DxrUNdu+MjDVglMQ4P+Li5JmduUSJhfDmvMoP53sPbKUlBZug1jxPQLPM7eQ
pLrpqEGGG5idc2Y6xTPg6kCVwV2yAXef9et3JFrmlI1XEtm59kj/94tdaRbYFgJy
uBLn96I8QHGd7vMjuDvX22j/hlcyzy0afloMsCEmN1XQfTi9wx1u+W1mdtdIkn+I
XxaCoWltZ9d0MEnh91AVwxeqDv2mHzc/rZ3oB3XhyFaenMJDsDkDrEvjzgaw593v
EnwYRxTpdd5U4w5SKz1ZXd/6/ysY3Xu6mGJ3KrtJBeBmC0QgzIMGA3C4u/djtzxe
vMkTfQ8X/2K9YouwWFAU+/7kSodsXqFtt1B/mS2bkBPe8Aiz4/Mol7fu/FGPz3T+
W9w2WVXyGGwskW8suR13g7j8a56Qr9GJf9dpbM7FS1U5/vneoo6E43Y9MqJjQfgn
8G17gbVTul69Z4kUa1u7TClZdDLwLBXnJGzA6NAq3YX4To5+Qjk2dmPnk/cEmKfM
GNc6691L3Jeyedw6uB2R1DkgeNWwIXGU06zkudxARX0dpMVTF3PVBRqyiWiudTNG
L5DVei+qGoCcwLa4fsCGW7SfTnQdHX/Wak1/6E4wME3biH8RibehnlvpY/iY3Cu2
YrCoLXgWvrlM2tvvEc4L1znOjsPBC8xo054c43WAE/MxiPEAm4noD7rw6imaXNza
W0l1oVb9r5QvYJVNtyFDzSDJKM97sITjFPeXpp/Tu6dcdlp7rjWPPSMyjKeIl1uL
JTmyXWvVxlNLChvflrV6m3SsbzDCNUFXXiPFVk3YeQrhALKlZtPF7ykiZyeFzylo
tGcSOUFh1as4F/MV1ptib0ZINWXL+G9d3KzebHKbFlbnCz6OszxgsWqHiVtH9PO9
6q/XhfaEUKZ4ja0ujK49w/VLoGnou9FBc4EU9fYjIjDyFr8CsCshNAr8oPEO3DiW
65L7P5uskNg7TSFP1X6l27OrhMeqGwFU9MP1hRVzsqGG1YNk3JeFPMCDJltKYDCE
7xsPUhoMDKx69zKERVzOPmnh9D7RkuO7BMVDnpxgKCaXwb98nGiAthiUy05vJ9k8
r3m//QSBbDSPRW08/e/Recad61OiLs+KwmRdN5DVCY0XBIqziYK3RNMzbK8zAPGe
/OWFyYdzQXCqhN3q3wJkHviHK0+Y1/jY5QkOpKcZrGAMn5l7XQnkYsTtxRocvKq+
znI7UKuNhpck0uOarHKB7qJIJU0azSkpHLwnXxdWhhyB6qWlSQqOkLuJfO/tn+im
5jIgQHYYfIpUf9HBaAS1VIOM6LGkH0ub+DoKkoGaOM9LWpWH9Yk2ZnjWppzbUatl
erVz34JMY/Z2psGwClf4vwHYk8kdCxc2bgjhBB1oYU86Nx7GJEubasL2fiZHnB3x
drFmx7zr/8N3pgQBLk3VumHIITmy1PESoQ3SLoJyBSzQHLscuPbAl2rZFcT2I1/L
1Gbq/ik/mkD38k7iNLRCxRvE2QJIz1tIkZF7+NXjYaS8hdF+ECTMD1H+RRlllwC7
R6viXlmKb/6O9G8GpLLtgchorGq6TAZcXLobWChDogA4Le5dWb8Tv/I416GLCltq
+uYWK4zAAmQZj6b+TfhwMRy/SqswcChvZMTeZL5AhrZrILNgPYbfZ4c8gG8b7wGq
Vrne4m9lAASYroceyfeXtIk40y9KH/2Z73urz2tow72mwIQneF6PK0De3hVt/5kk
kQMAX9sLZGEYeTSa1UAP5lnSZQX3pfKnDkLI1/mIKAtvYb/cRBhrD93gR1VpsO1j
uKe6k7KqOdItqZ5lCyavoyTBLVpUVSXMwN8qAnLpG0dYX4RAM1fZcElleYXSmWc1
QqQbBgjd1b7PGDLRshd+j5y2EHITDVFwCruFePdSGSxVhyBqzp/TgWQQyXBq8+l/
30xXcULRBcyJ4kunKHvzKZfMsNqz7pd7XkS1zVqOO77DJPcHoWkZLxb86/+jO+QQ
xa2wx1PwJ71lBlp90685gZ568x5AXJMuXNVqWrXAj4Opl6EMoT1mOkRWc3ej5pnc
cJGfBQ7FJJgur87Xv60Z50OlepupWEf1bsVsCDmC7Aa/Bqhdz5M9pV54bQylR2ox
BgXwft4Zw6ks0+w938lSsvlcmy3mysfRbhjwGVaL0Ac7zw68AAVI1u5QX/yNMtaQ
ELozhIVbfS0jZNgrZkGrudDbdwcMP2QBhsa8z/iRdRr4hAfRBFiq1+OLUKjmumrQ
HY1+Q5iLy8i7gUR81CqyFmPzuJDk0umMku42sCQUX3s0K96dSSzSRIP9QM8QPXK5
qAmxBRG/ImYEEThRUvna2CVYGdiOlJmVaRLdhl3Hp6o18VHl7GFyQuyD91qTGIJj
X452vHlltQP+Gd6g4aSzfKviPUDXl41fH0l5lNoj3Cc/8Q4lC3yZbQnnp+6R4OuK
+dla6fzu553KEtDYkmtpjjvJ3pOVI12pBljL/EBejN/+D7n+lp/V/aeY3J/y8Fbh
LqPpTNFIeMCoaUzpTIMKZUkFXNOjMFQHP8Hyc2r/LLlP4O+l+UaOEMU9/LiMssBZ
CPXR0Gv7JJTk4uMwePzH32kdwdohoSf//VtE8D+kIvpru3t2br/AZNz+ibJjmOxG
h7wW1v8UbAjGjgg1e0SwKJDdIs3JZUq8DM7N92gjSpxmCmTbOY0LeC1kDQe0JggF
9UXrxd1zHazG0LOnpUYCSBEb0mbcDmQooOA+8gZQ8sCxblaJ/Nkyah/Io05CY2bY
didFQYqKbE36guZWaHZ7cDpcuF9GxDYl4jcQL6dTUCi1FKSxrV32vuOZH+DZm0tK
NaivAPX8KMbIh0uCBNNBZ+hGp5AqTwKNLm5FHRqv1zGEu+XYIw1BNLFbnrqW8lCS
sP9/gky3njllodYMMufcUfuSMHdS+Lzf3N1rNWqOEBuyeZcedXEEhw5hdjkRbKpS
S4hHlTQiSyvgykEaEtcs6d9QUtjg/O7jgwMZY9gL9iPgEqwaL8fmr1lNcILZ/HAD
3qnrVRHTYc7MCG7E4VMbYlkrR/jy01IwHYzjJQ8mb4zwHFnurm/SZq+bRjVswUPz
+2q0qURRswzvryxtOqH8eIkwQhOBfGlz0ZERu8/59kcMo+zIjuI4POZG3kVEUHz0
Rnf8mjAJ4A7vnjRMCBmDd0Xp/UYbLo/G4mTsZRVKzkXKD+yhKeCC38h79BizMkcP
Sgiz5d2Mdz+vmWZdsFC3Dd8eMmHn6L+kCD+wUPG+wY/RdmgQvbrk3+ppVxBYyG0Q
pHqZBeIC5K4SGC+lx2ftV1KEM29NvJcdnwAgOTrnljKELeVq2IER5XkWpyW5AwQu
t8zDdCZ42OBQ4FHsZR20JP8REx5qi+u85Fegw60O07SgROvLcIgIlmFI4nng+JUq
5DnWP4hPnrssjuH2y7g/7Ww7rGC3WD8/5AS1HNvzpOXN0+7sXriUV3rEEDDhhCDb
AhNf0JrwvMFWRmcGfhcJvYtTmE8akygzbevY7rKSUEaZ34vgVcx1zo0RYD+63Ykv
KG19Q/8PYONHY0x5LbJ7+Awc4xmRcMrppt9YAJ5X6pt+gq98RtZxQhxuB/7gGwsS
/n7Lf+PVM3JUjUIsYS22ydEbb7FZ5Hp1wzSwdRF4FLJIiAMBZSaKiC8d2ZZuZrHz
dSbPFC7zkFTSNcnYHcs1+G0CTHhkmtqbnTGC877SPEifkz/+OwX4hqBcAI6kkps/
sPMOHLBwrMH4fSA+xG19GNA7kKAR1H0rlbiHwsZlB2oZs5CNSSoObUxb0q1vGJmk
Mec4LYuTSefYTpv5aesk35gfbA9vCzMgvxJqhC04oNftbCdafMARxuJ5KOe/TNHR
LrN5sFFfhdpkXUUhu1Lx1fq9HVpmXCrAwRuFqnneeyo0LLPlpkAIQxMvg6HTxPIz
vyuq3++BEZ3ZGl7JxwAZIs2fhDAECk8dHlQ26xB4V96zh7ATMu0mYjNPdRwvEXDP
M9q/odeTbOjH4mzw9kTZ55BTS8Kg6y9K/Nhn0JvdWp306IREgLuynFb3UdBXYFmB
UF1fFf/IA8xycS9yUMB0AJKmck/t0/t65WvXu4dv/RY+3NQFLMiSHIGLvFOlQ2tz
QLCoXn2U9LL2n2svq9YfuM7nB+NNhSxI7thZ7MWu3K6WJK0+EDCfr2cUNqoROjeU
Z1nSMzD2vmkhUoAaXc223AQgIKI6v/w2eL2SH0txjs3sAUyxtPD/KI4Bmp9HqI/C
A50G+xKVkFQDFPxWYM8WAS258Zv+rLJKPkz698iTtQCphnbUl1CdTm/kJ9gBiMei
TX5bYFiu/Cch12WyOzi4s5Ig7W2lebvrql9kztG79egZZHjeQGRVwlYelDwe2AFT
1dXuicqxqJz6MCkIlvU1Q7WiopSvLu9jS9Uy0Wsxv3JQEYNesdb8epGQDunYaAXV
MebtqbWNx9WLg/+YG9rE8VkaSfUrfLcF9cY9zuHZSxhZDCUSGS7aH89iBwWmJXL1
VOsu9APAw0kIr9UrhclAnppiGMSu2mV/7bFGbPSAu5W4B5SJfCrz2zvZlJaS97KJ
AzgjhK3Wu7JD9TLQscoG5VRITUxraG1Tjz3IA+r5hf2gCWBwsaHiwJvUopYLoEm+
dNhg8uYub+luoTH8pDyiC7Oy9M2figBJj0vXqjGSqNZ2PoZtw7Z/Od5zAbIBCZSM
pUPggPeE4IOtz/fEq7lVZJOyE3oOElVtsWRuzswxC3xBE7qgcsMBx4t0AZ1qbvLC
DWHTNTzYjiSrdPMLHiiEL0L2VhKrOU0Oi/1OcpvW+hhh+DVIokfHesSocWMjtuS3
ZtIQq4kfYn3yBxGRes7YmBWyyzt1AbZjtkp5FdbuzpjjMM6jgqm3vtPLc/fl/a85
fuk/Cd/Y7klIfWuKuZMAnv1S1D6DmXnKyUmgqThyrkVmbTC/mD8LvndV+odrisP5
Kl7rogRiVAGrbZr9uVTTnDrKxfK/8M+nz8+QuGVRDiRh4XB+o31MxPDWEUi/pV2u
1pc7SJtxall91iPJWZrTHCVR056HmECmpCnpXAW00hzx73hKJadyjx/0QtSOG1xG
F/Z7xsnLEc1OrZrwvY7HzkbEq9d26FyO0aoaMGy38L5/8cI/uMjzVvR34oRxzoWK
XnKyW0dU/3euYSUPVE5RkrUNoA6eHHyLeMgEhljF9lq3ij3k1/EXlYZLMM+o/R7m
9FXLW9X1vckepzmrV4+lA5K6WYutV/I+9M+9xTiQPQeQ4wEJzLfGJa2RgVUulZRK
tm3tN6q0OWp8NXd+BZU/nKYwCarddTCH8+p7O8L1wniFeEa1/+IERlMxSbXRDWD6
A6+UEJfov9qewV5/Dp6OMYEoTMIb1FYvgC7hgHF2TuYDjjWSeTCnZuZgofqL61tQ
uVmedvI4hQ1o3VzpHGe0YJq5oZHvRvNu99cpp9eVQaEeEn/Vg9t4EJL9vhAZ8jsa
tQ0W9PaYNYKQqfpNjrNQngAPOkG9V3HyGAeWm3YSyjnxUiegXoRg0+1qIWhn6PP5
Yz8rTNDbyxGXnfxUjOpfAo3t9Q8NLq4bNJpNj6I0c7tNIYKY/D69tSEGOzPT0ppo
1kXFTTZFk5yh/DItpp00ytl5UzSya54tbSK5iQFcEgAlDMb9efgABD1GBkL/HDTH
XO9bb18I1ZvarLHs+q27nP1sdeHg5XqipMlCeHfDIcvbLpRtqi783pqoJ356Ne0s
DK6u+2X9UDstC5Ir2yolyGb7l4YvyW0jx6vF0FB054UKUHyKXil7JJMbSHBheQ8z
IoNe7gNB2ZsBR00e/zrIUFPf0lw/SuoPfL9Zgv3IK4X7V+cFy2RMsXZ7LtAQznVV
4V4zB3T0iAx5+5Up9F89KMzlg+GPOUM18B2E7m5iMSw+izQ6Co1n5w3ZovSymYYl
YOq/5HsiblmahjS6wKVAWVnb7zBmdR+UI67PXjAhprtKC1blWa/Q7wgZNRxcjsG5
+NhtqmoszVyc9p8TdD+DeKUmRFmiix5wCTjK/FW5IGqphwDOpxazWP5w3UeVuAiA
fffHZxi7sjBPyqNy846kygovI/6rskZrl2VWbIpoZMP2NwBJ5caz+Cagh9I3Q0fq
OLuFPkXc4aa4YecqEsKMKjyxfu8iOVAOy1xH8S9iK4vYZ5yJ33UdWgpIAGgaWrGP
y6hRW106i0oHnwTU2iV0Kvy26TjdwyrFI/0YzoXqpeusbUm7mCGc0a992cHiJeo/
Sva/xK4+AZqv9aj6bAfYtI22dZDpO6DhiO9kIleihZU4kI3JSGjmCS2GdLXyaiZw
InWxRsQJHbEtRaTT/x8WHGQWxosctqECTx+USRYPHh9Cbb2GV/BOqLWJDXEtgvX6
CvgTQTrMQMN29v6QZHHsWYvA3oRxfXaGFus6Kgj9djEqJYIgEzWMukQwoQSBOVy0
fATG11qvz+2PZVnJ51Q2kslz6rR4qVowD5/JdJBKr3MLS892OLN0YEJi8qDJJNIl
AobpMtY7l40XSnFOLJS+Lj5n1dq+jXNIAzwhkcLNivIWMg1BhNaNYcCscN7Lr0PU
ZueNh0Ml/wBjE+psOY6Zjvmq0vvfmGc3yo0UWnFm4MBqUomWfHwAgxjFTIYRavWH
MdmBSQD2PLiyrEiy1lBkgi8kdh80Ncl0CvEYt/BoRjiZXrbAM1CeikEn4wFca7yB
ndDJKH85iccrUJ/p7gzgRrvNUpJbyvsaZMCqbtisyqpHmU1cKVad3D6AkO2lKC+N
7IGIupCDOlso5BbT6MdvVc+1Mw4deKY1BWPkTDgJPS9gDmArueDZrQiOx2+pBtvE
FIW7hzAwq4S+CwjirEzXmWX6jyhXSRkRiqFM/8zWX5hORALaAD1Qc6kpvmxf6VpW
RuIeSxVBy/8qi3SaQ2T0gONjCwryV1QldCZ9eJYbW7SqYij8T30GFJqQKPzpeJ3+
fXcR3OH5hfOETcEpi1kRsuf3Y2oMSHykvS7WiAcizif9WAh4yUZBmbJPBBAWLaGd
mhtJg4/4C7CASjtwmNPKhX+bEEXD6iyBS4f2GGJeiks3PWXQML3PHjLq7FH73G9q
S7rGzK/nHVnAmblKIl5BZXOzFdkq1dbu55wxQh6w0PKLt7FBKrY6PbLUBTI6xMnZ
maKmxskyXyApg3NF8G8g8kCMQWISQzbcYIlMtS52WUORErSsTjG1mDI+O+/N6Xyq
gQG175oHqNsmJGsRcJVW+XR4OTjzEjYk4Dhg+e5WDNPzICdNwE/7PhDY0fiBwovC
sTKU0Q6cbVrp0QDPBoFj4uOqC2GFiSsrlEqxRfNK6j9Ya/cMH9Q+7FuCITg5g/Bx
yrBLiu6tAXCF5LOBHl4yPv/osJDA51USf7AldrdMor6PtNR+JYrLbpJpRSTsQIeW
Up544sRo9v/PCY4O6EOzF33DR+uiZWCz44FA7GWu+1IxYSpBKxixIni34LccclWh
4lje0n44sYE0sAOGhjmKUPqQfv1msVMECMMAigVHkODU/ODLeY6E8qdykFdeTp0G
8XQcfnsQnQ9z88R2kKrhQ8UBauAspIxN5XjYxcYAtWWjziQ1wRmWcN5P4ZFSFjMg
m8ui9SI3FoQHhM6p2yC9O7oB9hXOvjzHt7rQrHvlbh8jzA02tIST6bPZQ9WphPN0
H81fWFCI5zS3tGNAbTTivvAOmfadO4AThzAEuIbKb0hb1Hiy7c2ubpDUggorKI7S
dJcTkK00MpJY6qxtiovot7bFb94E0a2VAhOc9cYl5/lci1t2qRPhmFK+bDzvhF93
MRcLyWbM7HG2RdvlN0fpy5ubIv4LOyZbHYMz+NUF9b0SCvLDHg1LQm2Dt/6d4Ldd
WfK4/aTjxxteVNAUC4di62UGrHlg4p1heiaEfih7msuMwZnHi10/NgDCJsi/h353
KFJwVuvEfFPsLfevGdqQkRKeBknBwN089utfyiODm1Ku4e9LgZuwoj9/DLUqiiBl
5HY54O+KSTGaHL1neKLyI2/7lkr1vUBFMQUwG+6Vgypb8nnufaF8bsjRF4lhNJVP
+x06617t7meM4foQitgc2BcavM9lmusqUpZQ12ia9o9AFhnn1Bj+x/tXeW+MGsvM
e4oivSCCfGyX7GXV+EmD393klDpuJTlRIptgBERWFDtehEwNiRT9G1FWbDtulCxi
RzsGyuIuGB5iODDRz/txpK0x9GgBJAZcbkITalESDDaAF1w7sLnbPWpsMQGVbv5X
ZPgqfKAk36duDMk+uYaxwTLtnBoxsDxnpGYjrUpFPCJZC/OTRjBLR4+OvojZnbrh
Q/HzjfIpM6WxWNM+u1IdB1umi4QlZSedH481z5xS/gVZ4g4DikZquUFa96+wlqZx
7t2NJaUYdGSbF0JFxJmzxD7ow4mvals7qbKOdqvg1i952/rJfLak4zYZuBxLYPRl
IhsjH9jnsHRIB72fCO36iA22uduwkZNzRtC3QzxCaujAUrA6Gk1G19qV1pNsIYIS
LVeNPMjCcg0qOsvfHH+RqKOIIYbslO2oDRIGi2ypPsX1NXmZsjQ5t6Hp20so3Cwa
ipuoz9R6zAbRvnYQe73p5UqNwRbVsjL65ImWGtRoc+0qhQVZT6V6fMSj+eYwuuEw
hPggLkpbM9gvTlY9Oc33XWqNGUaG9M3EO882kbTZsgkK3nSZh0W2XhsoHKl3Gl/a
g5yJaxaEo7xM7UTDfP3kZ5tsCRtbxHdR0KYjJFYWhwws7P5pidxlnSKyA41z5zz7
S2p5wF+NYSVI7ZYKYGcT+hjK3T2AasuJKc60sLXcUQ1D7BxshTcCicy2MHp1a7xo
KqaWwKAksZc1P+ijmRZ4XbY2++uuYFLBZTU5J0xYGlBom10d210jKIW+AJqONELI
55Msidlwpm38o/Rp3XIwUVASEPHbfLuEvZZNWBYhh3WLreADDLo4Pqjs1p0AAXit
XXaF6TC6Rqm9Euk/GtNgbVGlm0HHxs5dNc8FttLFwkVVRmXos+h1Udr8tGDzZctp
pc0gq5w2oyQR0ExVE7/htzRbZ/04dDRg7l9nLX8O/PfPwvy/m2L6Ut8TT6kzQMhO
/nu8Oj0WkneQxj4cFgcB/tQEqevad5HJgpsAQCc+VkQBP6EApQO/cCkygnxDKcDz
zvPrJseB2ZbnESzXJ7SBPaoWE82hd6C0+jDh2dnLSgGWPYQ29auc00dI2L3fjUNy
wd+f6Tty8FdvBUeflKdVsNOk9hN6fQL+RLYYJW9/ENNh6vc5c9tTmjgKX5vNtp6Z
5xTtT04mWCMxO0D+aZJfP0c9srJbmUGD0N1v0X8DGOw0bBDZ7daqq37VTiijnAcK
/TEehuDf5ZuYbzkDpuhZxYJiT+0zWPuS8HLXdbcePhlShjs+LUHqK9uRt7WL0sGe
ONQBoZcSmS6PLQBOAUFlIpio6JwEFAqYHYFN2wB7dmzFNPH24YegC2zPdYlsgCfE
toLLBtxXrNkbxHEMt9Qrt4awctp+AxnPnQYSs2S17/wZG5Yhhz7aD9guhl4ZJLID
s8QuM3LhxJNTe/IiW6EoDr76iY8FAYk6yKX7ZSKCXvcH6bLABayq6NeUUXl3nxF9
8Bb6EbpS36AiIs+1Aw+IL5J3drxZHA/BXT1E5KUA5bg/hMsVy4kmVFmqETq5P8he
+aTKBaIu2fEwaN5ZBfCKexkgBEsMPEElSMNMVrS9iPhHcrWkKH71gwI/7PNbqJol
O9y5ElpNBPGwLlKeUOMoFUu6eUD/wqA43EawDmV/UTzJ/DM52QXkDeFPZN1Wt8Sv
SqXoXE4mb6F+/8zcm+UCGdX42a0GEM0h83ETJB34CTVU8dPJQ8XQLQLtiFBwhqPq
hNAxUWEX8dxdMaJjEYGv8pLA3yqRds6sGdvFf5s0D8MMrb2pnAQi7iFS5T+dP+eT
f9G6u+ULf2zf+hmnm8fiVpnBHfQIocGC4EHwzyos6AYRKgwJ1pLhlYF8yJmhAwdN
uJ684f7rEXbgPuSLjirFDKKuo3sXYLhterUBW0THtnYUVgxDZfu1ZSCgFLbzn+WO
1W+wCSTDFKngdejQzL6NLBzF+W2yGUz9+zGc03rRkEkkUNEhs2FGt1oXmaxTdDjT
bOrRF+HpJL9jGseJDxNYE4w1rNBsosq6ji9u2DU3tic8UZD/Cf4o5kHO6PhHkZwX
Ylgg+CN4g9cYrMLXRBcUhoHv2kFM7gDCr7nDUh4+cvsx2TW7I96usEJ/9nabSTAp
CCUyY1xF7qCxQD3uTt4B2d2H/GhqKhAW09b2C0Tf27x5Zt8LFKsDZf9zsnGW0C5R
2fGY5+iDv//x1PxqHkVuVz0HE/FbMOJ7Qma9SfohBysAECuklVr5UQD99Vw2sNMF
f/ON1PqktEQzAEBrTbeoohLUB9iYqxTMF7lMos5Cbivx5qCvzN9uw6zoQfk41P7Q
VElpTGzVhQ0a+H+wqHvRGXIwt2vpfGuaEOd4nJnifZbV1UPHThCjHC4swr/hzsn/
56MIfLXjKK8/BkDLvmX/6t+YoXPhE8vquAfGEXtF5eUZ4sQ37v1M0Y62Z4RT8IKX
L090GcP+B+r7MYvBPTervMPUxYj+z6380dTN7gamL0McZcHQhBkTik5R859YcW3+
HlqlORxPJcaHGjuy44J1xwKR6l04I8iQaekwtDuhmJuCo3lRTMsTAEPce1ljOr6Z
WB2A4ddB9ZS9fjRtlzHegvbdzOtWFEigYokdeveie0CLIGVS/ZDl/1aKmhSsJ001
8Z8s7ayz4x9Dr2PrV6I3a31YbZ59uzjJKFry6bGeooUaomGzA6JIx7vI4Y8MFObq
uzYVAJ2+hY1qRIdQMCoLorkrdG5tvqcv6KwHHzAeK5MqEmmgkSGBbWdzJc4zKBXO
2YHJIE1c7Gh6hC+zvVGyERNCnaKYl4H8q2QCKbuGp4fWNoA48TwWFtC3EejitlWK
rclADl11U01EUlxD82/Yp/k6bWbIj7Klr5gj2r866WTVSyyviFfquCcU5sY3rk7R
h5fAW3r1swkojnuWo3XKcHgzS6FujdANb3d7I0lYwyTBX4i2FfRxu6uAHxOAPYCT
rSZQFsJg3OxnwZwjBdIUf7V5o52g7WueThqEsXlTbB7tK/oeqhhaE7P+idA5tDmq
cqwacEMgSz71CzTayUMvBhAI7UlReLVIUorO2dwyAvZ/3tkfQj585tYdRoaa6SzI
Sc1g6ZYKU4OicjuC4RsaWCAaXr9FRuVJ8s0lv0tFbx2/4euZwjNMlXtMX3SUTpUx
INdpu3XN50PjnWURYuLq/4alFPQmOt48d7x1xmbemxVzksZ2254vS2CPN/aX4Ts+
fT9g9Udc0RngwoyJbO7h9yevvNIGKtC7wc13JFdpmYWoHMcXDc3QM6pJv46X3NZY
iLCUVJ7qUz4s9Cj5o67bnnltc7B/cYFaGqCfzI2/qxuW4p5yRl9frrlI7dBIhqmb
ziTlsGiMwtKmmyS3MTj25dE2ZCaxKxdSAmEplE0vg9RZmwOEf4UHLrvgjQP+3SP5
jETcgYrtAdnz0/r6NkDopBRQjjCfqWWlCQRwYpTAJZ4PS3L9L3+WYabmwvM+a8qD
eLj/BCXUe3wLiWmt8HSS3q3ZWIRL1svslBm4UUNllQURPGgo23ptET1J8/9dtsj5
BknlWDFy4FLkxXRUMrO4+3VQtpSmw0hjRpA/QJ/Y3w/YHAflu/Uez0Zxp8X8K9d9
G5y1orOOh1cihFg8m9UMw+YzLKb7VYzP6PGPYXBUGgKwCfDfOFXpWN0PMds9zbg9
Rp2+SZUDoKNYbPyZdb6NOIKjYSlfn4Y4UFGTuk/oB1MPDgy6JgUAFx8nl3owgDlC
gLfItWKo1k+dgwdv8T4nFZXsRR6TK58hpI3KDw+Gi7EG6O1vTbHpyKvEVrJ3N76Y
dipufnGr1Eqb4O8SYXVGKm8XtrLkNdL29Zf61gGE1AQhAV8xfejhiQaQRu1b0QDN
hwa2BXICU8VoaAaZS3CFMKuaE6MrFaq3BmX82F+102rcr4sReAFlCrDuHcq9+GOz
IvX8TduDQ0R4G2YDihuhBZvSNvfIDbX6N1nQvjpOIWKz0WAfVSjhds1AL5f3XOww
uF7+pClsRMyAD+3V8/8ZEm045vK8p8c9bAKEWYh6IUZsFcscZmp8i58xe8QCCc4S
7BMZD++VTEioTVXzRrbdZ38IQT2drLPTCMxhktyAvXV+kMqddd8TUovcfdQ/CLhY
wKMxGkZO7THbsl4ClIRkOnMC+WwICOgwy/6sAhcEnDSixf/Cp8eb5e2r1x/m64y/
1H3V4sMg8GbVWv7z6678g6YmKUlyzga9Pu5zNYASXQjck0lNbBDcH41QjfeQQAdL
pb5tBXbborEjyxwWYAIiTFaIvH8Z7Bi+Pz8O/vho+J+C14PBHTPXf5fiepIvxKFs
/jbCZdrnyD6erby97SVYiijYZM5oHd8/pys9RijEvv2xqujrnWmjqhxXjjou3Vyt
j6G1fttjAA0T3xB3zZVU/j7QFKdVUJaXfNHXFDwDfZfPqNfZ4ddWtZLKpGVCHB0A
cqrPrU0/rv3rTBinAViwPXLdFKLvE4veIY31auMyyHJ/19Socv90H0m/xp1M9eR5
C+FA6FyLu/lo32QHQSBmRwzyRbN3a++sff1LDv4ZjKkaeXxssZpVQBR0IEiBSet5
CkaGbF0qGoYSydcwGXu8TgbWVr5FZuCAmvlq6F+Zd4DpzyL2HCDp9RrAK8nXlMQl
a432sk9sTRqTa2XaV1YByN2dijWWOowu4iy+vLgMlKRGq9W1TjrKO+nsRlGdwj3U
6KiDu18tKKhw+wKdPtARyTVh5COZGBodM2fXnUHM/2rBoJG9JG5Q52W7nGiAjOK0
MclqltK+Yu5DhHfP58vKUbyGfAuhUUYWYadvmd4BLQQFTmhpQlTkwe50hAednA9B
M41L0CANF7V6trPCdKe/mGG9cqmPcdFxtGVTYphzYgFTe/NhMktjjCsY+WuM585E
+miUO4gRA0esbKIRQ4xVZU2fQOjwsHH0DL2IV6V3RctjYKzPmNvtJKngTdeTW2At
HTsPVDtvjILX5CIJK4MVVRLgDtg6ZNoAHXL5I6/u1ZhwByGCsRa+OWfJOwixwGVF
cyyue3b1N/wbrYsSyt3Q5SiJZcgYI+lz+lmozKnrWQeRJw1i6KcBgky4L1M1NahK
NifBOQpnX/0KNNEnGhFav7T3LwHG38QIYw7ez+rxT7OYHmZgMkgJeRWhRWYQLlrJ
zVtDxVGsqfrqteIioMa2dCZiZoGE4+NEWO1xvEfb3GZ6gi3A5to+lkETYQdaK5Po
TFAlT5uPFLZ0GLbmhV4Lwz5t/HlMgCuzs3P9m1g/vsXXq6PJGrBX04CggmOZciD+
StBCaVwpC6ItitzaWWJtG24YuAvaDEMqmslpO4VUuswEa7eCwyrXPG49jhkMnLe0
7KaOU9VRCDylDbgedG3uhDQtvbjGrCF+1EdQVXka6nQ/Qfe6wamxb1+oiftCj2mJ
Af1NOI87DLilWY2AsC9/Da2A49IDDNWSLElB/dyT8SAuivYi/EvGrjL6m633Dp4z
1j6NUFZQOrd1xSkJhpX11CEIYLTil7gucn4EiIylY4BRy7+t9jpA2eHT+5Q+epVW
zmuifGiJDmeKsRm5Q4rLOjyOBE3NAipxI/6X68cKZvCxXe16PjyHCiJ4ZDLkXpvC
JTk1HU+Zy2raMEu2JZAY3/jsMt72eMWsU8Zpd1DES6qYY37MFGWyF78bqw6alZHB
dL6PlxUuKNwl1XPtJjrtdIeeZeZyDEscFmeIZ7/xhTlEZOrqlwrNYfgTZA5Fd1Mu
DHS+PLB6JqnXQTZbU0CgOY5tVQL2avP1zxiaPnETlOYhbN0r7pB7Suh/yOImW3zZ
JhPHGlq5UNhEpnoSwzVD/H442XC39EHfEd2z2WqV7IL6JZemvuGdqoyDPzgHaESV
FmTVvfhAoA70MgmMzaiD4bP9yoeQQkQxqZ2wfU4hri66o/hHYH/DD8Rzn1Cf11BJ
jezCm3fM0T+qNyKTUbE/OIR/LhdXBQ57KjBGKCBJM5RYmi5P2Rkunu6hvGoCJE2t
J5+HQLmjW8xvl53myUoT3RMSXMiZOxNYFTWAxtqDrkkii2tSyyUca1XJzE/g7Ni3
47DwsGGeGlBbTWP3Gacqvu9Uko6YbhEDG034ciDbdzLmHS1OWnjC+OnrupgMHZSS
fir3Y8t3X7G13Vk0TgoqFHtgCM0UfFhjTYQq3e6Cp3F4GBb0Qd/qpsFslM1sVLoH
EX+WDzsadigfJ7KYWzRaQUEIw6UHNO/tCTPs32OmUB/qGAGBUYX89F5E3J8qS3kr
cl0wYPabHsThgXCkk/75xeGiKV92iIt7WxEKQhsw3w/rs3uJZMXOUlihVwbvigdO
1PWC3tx9FMXLZd/gfQocKmJsRZSvMfPogW5iYK8qDROIb6+qmzRdesTYrNv89GY8
Ex7ps1TGA8NH+9/BkmaURV2/QLacvDdwpT1pQoeTU3ppT0CrAFDDIXQ2GLqq1aJ6
8N2Sqy+QB3KPcFQdWP2WUgwRflzmpA9c8PdfEA7RcAD5r2Vz/Ztq4BqvlAehm6SQ
c3U2PRPepSUS7nA5zuoAJlLq6Y7rh8FVzyxSux+r2BW11kWsezhHx1f4uXm6nBC+
0f8LMkPt9m9bKoctUr8zbNnBGpGkc75cV3MOmkCkZ8LDSIH702zy1uA3zM+f7RyJ
6gcjZH3cOyxicCxBfSuE182YsoW0Ud6IfS58j+0DA8F9noDPTwK49pux2o2kPZ3t
TLviqEu3VYrewb0sFlfQao2cVKtTMvCSjEsGA3uTRDEBIzm0SOPRpNdn8tjQ4Hep
ai8QT0Z+O02GV+F06fI3knAZL2SxfCvwf9+s0/lEe90oiKvO7q5w2az2uIB+GcnJ
GAUnoWEV3SQCVsmznX0oE2BMP/yawHqeSkXmctCjqlRUtdTLfOwfOvsmHqLAsKbF
7qQSEcLNX3CD0nfzPrNuI3I43X5VlrNse5Orp7KZivX/OqmP+OdmfY8MZc9BojK6
zvmdCp8SAk8zyxGK4KQqFZ42VrD7gFm+Y8ZDz65IktSfJSEde8n4BIiqQTOtfWa1
7ZuLRFsLHdl/pDHzfun2IUsFSajSGFA1JbdMlwNUVCKSsC90osonPXPqA3kUbb6l
sxoVFH9WPweDSKn3UK4iBGa751CIpZd8ybH8io+KYcWhwmodvVY04z1Ly+LjP2ge
Znmhe4/0G/WlpLPgHK6bM1DYcA/JTS2/x7zSLLfc4FbLvGhmLiZcYdlik5hTJdXj
rGSRVcR3n7/TRMEmvKQ1kOJty0ZSoyiOVRmtZxB5STtIwEhN3QdXqsF5+2cTYKC6
3lW/9+JUf+h8qicZK79BmTDD3MvR4L12gA13klYX94TR5cHKnZXUZrr0Lj5HgVXM
GNJ2LB61cbcJS3hr6nCDQLrCC8kfWDNT4t9RC66us4DTU3FIwWvs0ztqbqDGfyq/
TYP7Aw8KNly/amGdZOjIi5wWhATEmRkAbkzLCYpwS30pQMpASEFijeYRehsLPc/Y
FjXBfMt0x8po1keRHP7vFwrrkBsvfbz0fw5yINzsVrshbf6Nl0RwGdQd13kMGRsp
RdQjeb6qxpx1/wPUPQsqYYPpyQlDLOj2aLuZU4t3HULEFjCSzGLjagcd6w6hJYFv
n+AG52DOwDfuHDmkvgntZnYOk7Uahubuh44CJU9BqL8Y0Mz+Oh1nnfjyXpDcRwWH
S6NHO6LX42EA4h56kR25l+s+JilVLUlqX/X56ohNlEjbTn7zG93FxlfTh6rI6RWw
JtozPM+QMq6/P4PAl/B30KJ5xf6V51IWOKmGtYGxOmS3yb7WTGJsPnbTwbC4QrqT
l61bslqK5EgYf3KoeZBGLf34SiIwhWaaPVygPD64Hre006dmpKKFU2u3Ngtw4J9m
ym02iuBSVhWoqzWKQeisEhSo9+YK/UeJud11x0XxQsjmQSO5uaYd7QcJKFKPjnA7
ajtHSbuJx1jFX3xX6Fr6/08EMPkR5e9m6pSImodcOBCNMym33jYpF5gS/oR2vdTt
CCnaoePQhvt6uMU9syTvI1eOQ7+lk9BXLmgQrbmefX7k7TOnanDHIbNNSWH/2Izo
q0bfBu7h+SH1JzSNilykC61LHOoU2RGS9MwNw+VLlarxo/c/7gEe4tWX2Omda1AH
xieQUoBSAVetXATIT740o/G+wFIQCUZEhMWAuKWoSnQReh2ctB8goEiRXxyrc9ur
Q6eW4enlbqn0H75y9Du8dNZCnoruhs7CvRAVEogB8HN7PT63BQgKWmOaEJ1EZpjG
ZGrXEbhcSF+61ZWd0/tYl+OE2lFRB4icYw+Fb+26d2m+DCDU8a5brPjcdV5V1q58
UbYcqkJ0Jghc3SHYaKGGlI8G/VwXhnK2Z+JuPzRrk5N5f6wdlr0f6nP7kx4dvdOu
HtRkJ/Flcf0qyBPhL6Fg9A1ZJW28hdM/qXybrzKt/zvr0RjcvULjiGgax/y9rTdQ
PtHU2i2+ZUj/2Njr0ooz2lJpNZGiVwq4L3OhHxuCgUQdcWBJZXWy6Nw2G/pkQpEo
GwHonRed/oC0LPPXvoP8QCZy57mj9f7I4tw+qx1IE5JIVs5xOKXrW+JvyyqXOkix
0F6NAiR0PaJLK7blKpdMBECpELssYW6QMDxshrTChXH0Eq0ei1WWDwndg6OXBYAH
2oFkMw2natqGjNbNRpXP8HH8Dzsd67qJCkCSvyvMOdw06apB4iWlZqjYH2dKHbb9
5Dui17CTGYieg+evyEhJFDPc1a0VMT7ti34NeDZKwkDbffU/pHMSsL+qGAnu0CSJ
fAGK+4bdgOZHi1VIlxKLUSQSRFL9jsCe4I2FWqKNBVsY1yFmQdX2Q/x1hQAvJaNj
/kdNfxRAyq9ynzlM9cYcBZ+KIHTb2gMJuCJYVv2BGXb0ywwJOBs/JcONeXw/xAsO
kfFVDCMG6eE3360sX+gCWmjTzRbvj7hYTsZkH2Uw7YlhxScaJ1041gzO5w2PTJX4
nCAKJ09ebuWepdB3E6KW+EAn1bH4CZ2KSkiDCloT/mc1BWLNTidFT0zKJ45DbX+S
HlLwC5jbuWW/sCwuc5A5db0ue3AEywDcU5k/hzSmyDa5tVJm2rdMOTkEO2YqcXi1
mQWmSiNs8gfUpUnuIgrOwAHfRY/yTsw89UYlURDB7L7MAS7z52K7R6cvZVX3LB7O
wkHDuag+cjMV9FrfItut+GXoBDip8MYwtOiDSB1lPkrTQ1RiKvz+T2mf7L0Zu9lq
9WR6G9yzgEa8of2oksb2ikver55h+FxtcjbJq8y6J+80ZBlxRCe8g7sRW53fAhds
rqlDGzEluJeZabz9Lvr7R/dyM6Q0WLQMLKZhwP/qxQ5MyetcBP1cSQX3hLBGtaGe
jfYQhbzO51Nx1mX63VJ9vqhakxMMAJne7gMRIGLGhp06EzgvH70RG9kodr8656V1
PmyfGvzr0f0OpizpIG8BkqMTxrG3H82D+vVTOghkNyEOSTx7KXgBTT+BAVHgOYBV
oipKXV4ek5ZBbU71N5OrnR/dlE+GcTJJIpq8ZoSP0BBAPMXaO2exWGNIX1AjtBVG
as6GtOmTukjVIXk//InsGh6mX7dIndvJwXop7C1BOTO02DOvBxuojcqWIBsfrZbt
9xsthfcrgWgsBVsJHlbHcgUwQwsqI81zhBdU4fQw3TpOK9Oed60EIwgYwdUNlulS
9Xk0R+/1yy6XNEJ7wkHdHjTDnTrGYVvbfioP2tFZ+ixCFmrP6oKff5E42RWUK9uu
X1YmNJxbz6zrUhFyGNr8Q/0g4CJSkKHDNUZT521KR/5LJ5BHnAtXgQ4aSmJ4ivF6
ZjbFOSpuVuDaIVmCzRLbEsh824NIXj2PfK6Gsq7yNbpl2gaGRwMoKil3FtBihNKJ
V+ndyLWtOj4vqQ41hipY6Gc3MWYoeD97OVw+bj9OP9xliNHMgfSX6wt0Y02kgol/
u4yuOS1gZEo4+7u5xcc529opBLlPm1iNZ3wKhZLcta22yaAb4FLmyjtAaXcS6W/A
/WW8hKs1gxl0+anoD4SW8fhbMaBEWlm6mlZp65gpHcY/tujOWXv5rCZYEBCYNLzB
evsvd5hhj5O8jAwZs452FG8rdsSOnz1Mpyb9apKxhjTGY8+yiXhZkXRxo8GiRjY6
S6maudhXi90CWVFab6G0YbWrCd7A27lheKPhArdcfrUSzKXgQx3HpVbPs4CUwYQ9
QTDap4zepEF/kPxn7Q5iL0S1azD2CdVcN78YfgIBW9tNmcX/9fCe6khWMaWi4zOa
t76+QEzOswuFnctFsk/4vL5ABCnxx0qFLbHuQhPB+6sxMrbl2Mbnj8Ih39ElIO3H
mOIp6apH6Z86lmY72EHf2ilb4Dl069qYSMWqPpclygo7IJTQc/JuhEX+Bskv1wod
xbJ3pU59IcDVAXkl2bZmJDagEBvAjOkeZz3d9weOni0c1eveJVPTWMKeJ5PFMVT+
k8pclNdGWigfs4/dpICf1h1kn6emAygHoqpGz/BSeLWvIUXg62l2vzNwezadf4aU
sFsT2hkRX7XfmZNVDGbgWEon3Nm+NFR8jwMaDh+hhq/O/xTiaPEknjpGKhed7nZ/
GDJdPCbfo3otqkwRlNRyE63mjuCX+/DaxFpVfW0DN8U1AjyqpUC9h2VQzV0iohTa
QdSFoyjN+ZUHGENfS+RK9IXN6HjC++KgUyVX63jspkyFoK1BdvtPJ7qx1qintTRm
0KlazoJybIfl81/rFXer3TXig4C6DSsCHQzk31pLQSbBY7Vw/Miu5yB+Mvj4zzOb
kHthFbMkSDDJr2v15owj7j/lraHPfoGZIW0/B+6afyFvDGd9xccceNm6ZcDQzpGE
mt64rqSsazT+fiiPU9BGER4VtayWAuoaGr+Wj8dLMLFT2N3ar1XxnQaYQ6j1KcpR
liGm+ctNFBuxJLw1yHCDViPcOIknpJofDo91xEssld+S17eXXKvnSVDNOu7u88n7
+Utgmxkvsf8zCxCbYg1g5VxIBffPYOe7dy2/5OLx0xwS/aRJeXj88Cq5WCNJN9bk
+gG/qWGDciKUwW268TKFEm5AtriHKGAwwxJStq0qU7RYD6R69IEonaK0qbpUcHrr
2CPcGrnU0/SjyJP+J8k3coLGvIV2zy2JGf6fjJMMTRiqjGfLvObGkQO8eI3SewBd
kJLc93ZpHg/O2NJZgSGCCC7KnV9BsZS0vq0yS3SaDAAzmIAyJScOE/Fj3m806q+S
CfRNJ46f0y/Vhp1UmjY3/OZWtd9fb3duuzXvKgkTqn9QMxhfruwaG88lFM94spg9
Y8bzixrw0TxEhn63IsIoU2AwRVHyvaP7HoLsp2ewU/8qsoirB/0IT5REhymeV8Pw
UJ3x2SV8bUV02rWSuCNGs07ZFjvFz7T4vE7d7W0XKlpDliRJwb0RoFggjJw/4LNu
yzadw7DiAlqIkB5F2cXDj/74jDluuf1skvGbreq0P07vT0keW/4m5Act5JpD7Ow9
LeYNAVW05kHoBIV9ojEWVVIp+NK9jpr2u+6SvHsfvrm/dC7TUzZpDipMUofTM6AV
1oVLDWWdl8+iwnaBQ920c0WH0utuMFYUgJkwHU7eK+ZAmPdlp5zxDVRWgYNRJ3wq
QUBSnIZAGBsBRIhBDZnBtIWCvFPAq15nizChghL42e+M2mdUKEL6Zx5pm+GNaCDl
H6P0zlxw8e+rj4uXGa9h0NFS2UkT+Lbyk/Bv7US59nNucBkvDMrx7VYn5uVNOTYD
vEbRrNpUKIlTTHEtB5WDsGZV+tTY3Qz/iaxezqlsu4qWkrfu7suT4Z687/7L81Ji
EsNQ1OPaG7kLMvqOe/PqVpvpgsfydlW8HZdWR/DGqba//zpcZi3owWQ1rOiSRJ6/
OYuJKLmw9T0gzD1NMwTBlgLfbuKMclY63V1MVsRTl56ldT8Fv9C3h2/7kBo4I93t
1uae1sQtrP/nSuTJc9KrtEjS0W0McnhMD1JJV8NeW/Wi5QPw33GIClHunLQoWAh5
Ps6QioyGstB5xQYq2XHAQeWPzBjkszYrdgE0nXLyBc7F6chbQ6645mnXYG8ODB1I
W0vLRr5IAOQALPW+1+jG8qJp6P0mA8C3Un7tPCL3Dm0B/+FNwgtFV2vQ5NC9Fr68
lOFHp4gk4fJfAIPA5idNocvBpShwCISR+1uc/nl4AnjIWzS8s1dSXbitAOreGyds
yHFer/RFQuITHA684fg1LygXF2HE7+OONw/gANxChb8rx8JcXt3ozqfu5iDt9RSs
07UsDM9c3O0FjZNh/+3NL1CLc73kpTk1P/yXZqzl5iCvBolqNy47OGf2wYXg08vt
Ox1ERGdxezOd7S3VDSgL+J94u5YqQvGLFktc5vJ3aTUIJFF13kA94khE7jH6mR19
ACU4ycwYAQVifPMjI1pwSyObqj/wXpqiDDddyv4D/GX3OXnL3nsCXB/fODat4Job
JoXSwvjdohVwz0Y6Am7u5+8n2uj8HAEfXZLWs3dCYOB9UqBrvhg75sjV6CS5zElM
JLnmWsHV3QQNfIMhRcPRxyv7SP4H+/yLUjSUJysaYEUxU18arHJHWMS6xC8zHVHg
t4mYnDgvWY1afoLIIbjPKRbbbsrdVaXSqkHruM26OS62v4Uk26wLjzcuEgPMU4VX
sq4mDuGcDnh6BPuB07IKvoS7pjaQnVSltfGBhNDZbTQcbbYptghtTmSAOXODp08a
A8FUQTtEBs2bQLUexItcmmS31wFBjRhog9j6dCWBOVEK8/Xbu2b2/Vbg8x+9IJFT
bEQWrLs61NAS5/Q5w45s7zeU6qNut2YW5eYnc4pnMt8KUa064a24D919YFaOM9e5
QWj58pq87/KpdtbPkk1H9zdUa8eAMiIdbcldtA1etIBDwX/bJP3k140Zk9Zr6z4W
pFXHNTRLN1Zjtr0UOXyXi4GVlgKHoaNwDuOumPdJP/gUPJdNsKN3KO2r6glU9o+J
RX7tqN6LnRcD7ZT6EC27HTzDqfZDdJYOSFR0y+9rs//Axlndp4MYeEexh153YOsM
tXUXvE8QUOPc3dLrNiw6LZWngmFpX6VGDkqyI7hkNFGaXz0IcfSKqEEmI7DS4Gxl
G7y9LOjuDRGJ4OEX0cS8VY+1RfSjXiK8jfLDS9++gG+2RXcRh9hJlQuB69pMqQF2
GyK9xKCluQrsV2nbsQBTLxzW7j34U9pWBRoPE+sO4txclcLVztklk6w6MiHUSNJp
AJB62TpTYGjfcYOlVoDGq7zox18kZ4SSX+nn6/kMknJP2BOznvC0Vud2XGweodpi
krY4vQ27G4H4ED+2cZ4WGDrnlTIKMeVsmD5/hFicux2M+hJkdloww/UARAus4E5c
8bMljmar9sVPzDbgvl/So3V6pG0ulIwSREU+W6rA2g9UrqJsplcvUXs+fsZGScQT
Jhki3WZU0MGm3gxfeLrlMBCkVXKjyK97h0Hym8AD/8tfslZLmoaKXieGHR+rGl0W
EtQAulFhcftcvhvodnFkMKXAtfRK859EdX1PXkZW/MGoo/ZYLN+eRY+3uZMrPqFY
0VvbU/dFm2m5GwvvzYNvI5SunYMfGlx41/s8hQ/beB0ihT0vFKiJX6GjGznRFFVH
Bq3lZWjRdURDj3Cwh1NDyYXavXIsZJZZKl/YsP/D5UHkyc0lOpaPi/XumrosbN1B
UmmqVaqEbx6d5eygL0bckIk7fCRFK+kebZuddxIYpn3m832e5z3Vy/Dg+egZb/s7
g39M+LAt5WbaQe/ItFXdFDNMhm1V2kZ3DELannPv3NGQjV7JCeNcmZEYpog9kdXM
Skp5ibCODWzw/1iXfPxbqfwiKZcuIRRnnQ9bZoS2aK3iIyKDhpAb258E4hHU/GJx
OyJ/CdbGUSfXqoTVE6ijgkKj1m0ejyRyqmEQ79cCQMd7IEuoRvxlNGcQmE933tDN
eIH0CaFEmFZ3qtj4+lHKePu03yLwnYY5pAsR5fyqq6GMTb0jwuOpnYHHBWVUPjSL
28lQfEuBHeoV+YmG99mt1VwPCs/v2u5JMl/dZIt1GwDqNYQbyBjoTVJwNq7fioFV
ZZOo/2r9cafYF7BB1sndwtvfOzjJKt4IJ5BBcWO9OZC7To9Qrgn57mCNmd570MWl
t289dtfb4+bbMbmTHe5k0mhKuJxmJLYD1Gw9+uQ+wzWFD3S/xe7HD77IypOmwbZn
l8beBrkIPQC6rAhvlB66UsNNFj/C9Bv5PUVG9lebRKKooHijHfm17fHh7HqqPpUQ
4Jy5RusVGq90Xex9vVX4nxCPS/H8QANaO64ZizHebUCH9kP78swWKMpsJB2EqNYv
ZZYd52TUGy8+Cw5wavWiv93rGujDcbPdOP7ZSt7eJB7LvpjyaO1accAqWqEpJnDK
4PA98cnQAHKeKnOBJT5vpKjJhjxEUfqSYQsTc+xJCpexYqr7fWaCBdzKbO23wJj1
/yp4EXlvtAph70M2m4aHoV1IWFF/FqQ+a0mnLxJc70CVLHlr2yxd406zRSjD/kA2
aY+7H4YMaY+E7upTE82NC300aNiSEHhuby2uZ0Zs039sTrtWKjDZui+kRnQiZXzF
94PQJ44VdfmDgUrmcbdEcn7bhf4OjSYGkfPjGKb6aJsW4vjo41YVEOrc214WQJ18
Y+MDOJhycfvFlwPIYEmNeJaL6ioZJPGfaEojRp/A1o2nG1JpZbPlY3JS1LXkG25x
eTjzFLZNHwKijHJwEwZU50IXjRaxXOhGXClyzHRLt4fHq+kFSGRbZhL7geSI4aep
LktxolI1duKhnlXZEJmnCxt6x8ncUZ9SqY8C3cIeqMiK0l5f9wQjeJhcVjIqRWDY
WDMMqMhW0k1pUwbTOHFtYTWXywrl2n+Ca7JMm0263WbpE6vF0oLLoGjl6wHa+1vw
iff1ffB/rdavgmibRqSIwqWrXgWTHElNJkArQ8VqnCoD9D9cTKRhfTeaGEgydtOo
lyYMPvyzcLES7tzSX8yLrHgbeVy7bygbIiwfNdJbmNDyc4SxknQdgZo+EM4lntp2
O+aza5er3bzypph4+kBP/iwqjvs9C5K9Xv7Swe4SuHn86tcX7Cjz4ooCBXrZBtBF
iY7ULQWmjiS1wZgjErhTeyIXJtkC0kX/PgpVgWWdb8DgQWm0QNQ7vs7ZGQfqFZJ6
pa17i4VQGsK6lfuM0vRB8zyAJV9YUwuP1t9hl+gN4XqDVhjY8V/XhxMlwcsNhI6X
irKbW4UsfapKVY+FPmCIVali2WkGwBPQOGe7gPGYY1krW010yUOYotguubjIvhzO
kLO6N7HmuebSQTr3w7aJU9w+RvglQDpfrqspe7BxmyOy3ibv1oaQEWBu7f4De1BN
+yuB/yRnXJcBsPUT4DZIznK4Rw9qZbr79vHr2WaYW6YNZfLMoEmh7it8zlYFT4TJ
96msPeCv5mPQ0gcRrdgW13207IgQCgxr++YRn8SUzioPb4YuBIvknMARHLhowjwr
xWtyIdtGHRo/Mv6+lxOek4VR7IMAllTRU7itaVdA8/g01J3kqLnhOPBoFJJUJbML
kt5IoerruiI4ACLnVU7zpfSBtrAo6gr4yRnxePXvOmEVsVKIh0A1Si86GOpm6Hae
n1FO/3wJJ3vsf/CDL2Qn7bhK8SHqMwDZor2ybY3dyT+IkjQuhG42JnPV9NQd0dfd
vRN7ZaLNQS9hD+P/2iVN7uI4RWWmV8i9wImRQBOGPYFTqo4L2kNfG6xCGkrKSBYM
iF820w2mThoWmKLipMVUh6JZQBkA/NMrMPkWzdSIrOh7BSr1dvCZjpb3jdwgx1nB
bZW4+gYppwQGlPkApJZp2UOVH/z3ZNfVg+k+voabhf4ksX4pxjIdZ6xMy6pCQ45q
uzni7G5V1RFu0XeRo/W6KnjNsIzqjD24zxfxr3kGL5THL0U6GIJP+N1ZIzIHPvTF
8PfoU6Ze/hw4gSnqdVuZec9c4nD83kBOSjBp3tH8xWIW80Vz0oPKr9ouwFOFFj5b
O33ueNtp9cd0rvDAJmy/GD7teNebBMn6fUjcT73W6YpPCLAbn7GBav3+Bkue/MLV
dJQifKkHsZ7DYGkxkviJPK0OKGceTZYEcMB+dhJvVqgNozH6WBaYpcOeQ1+zBsPl
VFj2jU+9jTN0EwM+1PAjGvP1l0ousxyJj6dQATss/UYULd8z1Hja4amOQWWyMwgB
9Py2H7I0hyaSFQ2g3fyFo12RPxq2BU73wyrwnNeyzHEKstbhKcTRvnCdOkNUcXpA
dUPy8fWYYsW61X2HtoiXnRUUl3BXJMsIwm94Q6GECWVyoLhDIkonKwSVsEb41fEU
Nd1st3EgrfSoiZCwHrkwjmnP9bB45YFChLK3ad44K5oaAjaIN9npvM+lvsjFHNLC
pYae3aqIJYXXXXUaiTDQIp5RI1cYzDQOewTGrcuchPaPJexOBxHfUvl0KO3EmOjb
fyvelQiohw+Ed2RV0ZKTy/0MEaElUmlChrQnvecbl3t+b6M2HKFlBdd/0Jj0Idpf
mDKQ2KN6jUkNI+uds7oYR8pQwznY5G1KT+G9Z3hlIX5xFfjkEfpET3ZachzlIbCT
FpwWpHz7iSc2o41GhtI9078UtfUDORaqsO1c4k5kjr35YCIKi6Dl2PwwHqp+yRUt
BthBAs9+uCZCS+Eu7MuVT3TvOJjpmfNexpKGDDuhlJlBVRy/9/dOvGaIPfFUMJCP
G4GAUR9RUnoAwj01gvBW2tWBk2Q3tbPWrMR41JRvMufyck8DlCBI0HrrYCPUsrbY
3KLy4ph0WZaQeCAXM6EH4mNeDdXklJg5j/LuQxTpp6knGE8kibSj6yGBj6mOfnDZ
8JP9yK8b2kshzfkLo5MJoC1yUmi4S4fKCISqYTqKbhETs2Hx7Rb3lrBDAfmYdpMR
TFO/0qGdvng7WnPbZNOojRuO0fPzHElkSiEh5ZI5FzL4aWzBtx3q/j5xsrcgtV9G
dkj8ddcJYiIo7Z1aDRTBL+NrdzgfF96FLNZOyBCizMGjOGIa6labb6lAWym59C+/
OpHP8vLHwcuMTUP2Sqj5WLvHZefkKoq7kj3cJh3TBBZzzSQ7uUxomIAM669C3tzw
ixZztSjoiR80NvJON3NpYTgenWyzzl+F7tD7LekvgJ/LbIa5iqPPj2nzmlvTxLgu
Oz0+bmFGb0SCwxuGNlVyR6TqN7/DJSZij5ldZbTHYSL2N7BRnEydJJ/YsrQ/cOZh
F3ePlGO8lxyVgKxFoV/k/0SkajLPG3uQKi261jPjLuxgBvv2J8Cteqdd7HmDCIV1
oecquVmPY7e/QVS1ES34nRJjsxFozW8DNaL5eFzIw1NMN0LqMNzQQD5LHs9iKoN6
IejWu2F+3nJNdJBEpsRfXbQpduy1juuDrf3c2V5sOFvZDzozMtVgrLn25/5B0VRX
AnnuvHnZHG7aGBYZq82F8DP7IE3jzDdu59xN/Jg7qXEVyD1iSmkYbTybJ3YQSG/Q
vvLAQnZeIN0Ek0gOPDvdio6cNbPhqj11P5sARf5XDzWlio7G6lsfcs5TUcAEn/T/
ZOy6gQBEb3TqtiLkMK1EKYqW2vuIDU1AdMionyye3RDFsivcNc5rU3cSOK9qHprR
jhmKFEogaCeeOaI4gPuLVnal5RgP7W9RQhnrZYszl9wHPCwb3bsu3j9CUaFQdq19
GD7RASjwVHDzv6vH8xB5w6MFR5m2th7RitoKV0u6eaLwDzQpEG4+R1+3WZGS1nE0
kkn3AtP2mVdRW6sBDwLpmtC4S29n0nH95mW4scKyV5adpoYl0oiDmVb5dTJo0JsU
AMtkI68d+QZwYBXbLrEKzYw15HQD1zrziTse8MvnaIvyFSO1RLq4Dp98kV3WW+OO
hCX0oqZSIi27xgFyEndPqp+YAlVeEoLaBZaNWxJagSsUSDKylveXqoBcGAaCk8Eh
IjI+egwtq3BUvd8tcn/j8L5gCf6rrZwqX8nGZ3WyQ6atpLFeaRcWMZVpbqtr8SlW
ON5e0zDalcfeaRrZpZK1TdpAGcGzfuuC2zql/h2oIiZIkfEGNPbskvU2hhMtQqcH
ORnpRXbkp/qzukRQ+/68Kxan4vog20mTkz4YAw/IOwHpWALsjhcJGfNjtCVUuQid
j9NrTdAjfd34pXlDMX1cHYNegzrD5xTBEocZFHtzLBtOvtsAET7QS3X2f64fNfvW
smkWaA3ydqC65wXmQr8ZI+iXY0abwnMni9iPCo82xnLG2dAodbsH/B8q2sWnMw9d
REKFiGyEBuKhclwnvljDcyzlxA9V9EXoISYbNOyu4F09y1eGEVUe93Jbgat5jVNF
O+nZcn0wWNrxdKMVTmx3lsZrSBMTHSMLgGzTikvg/WaNq7SbqB/g5M+2jnEmv1hu
u6QIaw6H6GnnHO98dBPuT+raRLFVoeWw8RVik7FDpS3+IJ3X67yRr2BfbD1DjTpc
ZOgutLD7DcvoP5GzNUXWBz1gsN0QVXvxz/PVEEfNM+zs2dCaKvgQYxnr2XTBFNgt
r5/Umc3oMKkgPTgrfLobBFg2xkMP+TJPY8p8FOkBqp1fMBqMbxQbNUy9ykRgHyZa
mx20yhOFNhrxzCQijEkMAv4jzjNbso53mJWfnv8fJqLRdlOHZquT4/IDzjLJLMza
pXqLxsu2LbrKauu66xA7O/qK+lyKG9RTnEINo4m7U91owNfs2pUOP3y2T0sNQ8Gw
5lta/5bBFk8KSW1+Q7ysOtHhbI+DnuLcdi0TyFswxbBqR5ospk4JS9oVQpPfOG5w
tIORQtv1dmrZ8YC1MWSCHbKfGHy4w6AsH8M373gyI8mqEz5GUrvAtpw5GqPFMJE/
8vTW5J8GDQWjRdGR1cDmMsqsZm71kGvPBOOhpubm9NBQ/VFh+PIkZJ3LpTkfJP9h
zmLsH7ekpJDLl+JNgcckdGCjkRC58O55XCoYLybif15dOM+vNhIFb2ILarz++wDV
OhUlEX+/+tmvjCzqNFaCB42hjQOMS7AuoO/G8y8N8xqUF1psVbNdxdvgv2RA0J+K
IaecuPcPgVcDKp7gtPVbcx4kAJdGOKJjx3CLc4zesOtidouvT/o1AjOMnAiZdyVe
zLbyAzhUfXV2cc0n/QivVpL0plpuKKoUNuWSbm3Ccs9K7z8tOuKPH2FGEElTiKW6
q9t2DvpxjcPYUuqNEFOIpdJpO40DqlDwRshLgVZpIWk3reVPimht2d/GLqqkuykA
VGe23RJTSDdhesDCUGDvnkETV+tS7C08Ssd8XwLa0aBnuFudDVmWKRV42z0T46S+
I61OACzDMNYozjStSXzy4KRTN4jwqw2MJm3QY3L6F60+aNkikeVDY8zqaTRWDmNp
C5SGDyoMhaHml2lAoEboa5oVknUj8sG/CRH73vSh7Dz90nCJG7TczGIa40bxBBjU
UJ2ZWMfLQA82QOouwKZu111zzrr22mVqu/OXZYy/rX2iIvnXROySNchTds4nEqvh
d+307aL0mTxpPPe/VRyNIwOP0A0nFVkRaF0Zytz+HBr91iKErtSBbOxZWIBRSifg
rKIlphEmHiS6btddzEUPIsNTz7rJ5GtoLCpXPq02nzPzpM+lnZLXXiJrINCMk06j
KQyeZKTGpJLnwlGoTHhxYb3WNzQf/UcLvbcCviyZVOtvcY15+At2A4ug4hk5e6Xq
JJ7t/OwVRw0KgyeyIe2ShlxALyaQlC06glF4v9r0EOQLkp1wwPwwovg+VoxRvxUX
q4E1Qpb8/5dgQiHhW/J2yQ5AQ1MJmJCki2vgr3HvdDJEaevdfmiVLPUvSJfXovW8
Jr7GNclM4Gj+ZdRv2vDglQGFl/w/S1A4Mx/l0P4Q5d1DzkO85q5BisAsmPyrM5K2
s3Qy+cZH+Ee1gFGesnUjnq525gcst8aRlBAqUaLcgnqF/yrE8cVCMgMQ0kJwXvVD
F9y4fg5WL5sdKVuSYWl7SGqsP8wG7Eq0OfqcAwNjfz2HNS8tWNnNVItVMvJhiJyI
ClNjXQwx5I1OSER+u+4v6s9Txm3cQbsT70VGTkbpQNs8Dg1n45OXQyev1Zxhud0G
Izn2rwemd4Pdrmb6lZmUGtcaAgZIDZGNP1cHrTbJGw+2y/KrEPkPoX77k16DUWiU
xkdZYIZySWaX3IJPoRio27qyNqRAf9Xwgq8JNa7Uj1GxDc1mIoriqPm5zEyJgXVA
E1/sl+r3uD800uY7n99dm77ojjp5vGFartd9XL6ftZgkZGa/5JE+DdPg3Ldlt/ai
UrxTtRjhpaPLAHXYDqWo7BbqXwyRGPYQNXHMk+Fgcl1CGgXtEz+iXLEj3+rL8lt4
4bSZZqKv4rdyPvXsoneZIoqqerlxbsBqo0sHsRPATyYAxxo3CQFTNRV4HCu57W0Z
Qi+mexWXRpqXepxiORrzvkctvXpGultoYADHlicV4SFZMkE7az9MDCOqh3oUk59A
KnmACDdFnodLiEtwDXdXSuzG+Wm5F6+T1v7arl2pbWL5CIatBqrc9NzQi1rUdY6J
ppggQPbTc56sBFplDQcHBiI7whkOx9EXbr1f8KWc90W4+ONO5c0GjE0IsjoDxO0u
D85l/xNCVroQQcXtbd1kO6cbz4pDpA4D9tn10Mlzi/tRoEZyhjWhjlC6/JDRlFuq
4UdG5mQ6RNMWIdLGt1e33e9YKARnLg0xDk0g+prRi/g/VjCMMzIkm06CE+27YvIi
7aW9hRURag9DuKTPtCHiFwcoq7a1jgfMBTrpygRFDAa26kdT9fz/r5fSFPwKEnFZ
4fFowNuyONtvVGIe3gsQnZ6QIfViinfMQ/tT9x/RFkVf05t9M77ps5Jxd/Iq8dNi
x7yju1UIcmaStqaVCKMrln0OXRZhYTL5PdZkwdzkLBuRIM4DzPxJ4v9JTFIQ0EMN
ijYRjOb7XWkG4RPSeyx3ADV4ZD76qEyEccyXm4peBMCds76vOaM9J8/+y6bs+T+C
kYBRslEEHI3vRfxLMY1mZNkElhoGoyCuaEbKlC7MGYDKW5svXhxGMGdZ2q+o76P9
MHpGt2S/+fDqFZ0Zo1bWbBk++uA4nk8GpvQk05/wCq/U711ZEFDfxAJhRrrcPaGw
Kl/vF27TpiMnZ0w34Xbu0WIHAbC448WEe8U5JJzwvMndmgWrUnY6gzPcOUkjzfrB
wG1sWdIjOoAoqj7h8PhUvo3ckDgDxtJs2TY6xuLeRfn0SgCc7WAJyU4PSt8l7UHG
CkNpZmvPLyBzSw+f3by+1BTZvTKm6wrDeN5yaYSbkEv/feEuUYELoyH2Y++ESwsn
sNw1L6etyFxT9LvpZxo762Pvz9hX5DFboTCPOef7zWaZ2lv2uCmifT7vzu8OZhcB
QGQXCPv06dqHampz/69/pMYkVdJLk5oceMGMt45+r6KxbJHxEaVrNt2xx7JEzc2q
Nu7DhcQlK4rPscP5ECgP0dIRzDhRPSY6syFcy1n+U8Cp3ubImpGdUcfG6q7KifsK
6D12ds3OLvN627mZ1p6oOrzgRv2l2GYC/RYWviLZ6hBUnbbt4FUv7mwHg04PcCfI
339XoJ45TuRaOjYCDaaYdFKh+C4JKQJ2MVdJ02HKwylyeVywKxdvUIPXqeOo6M9U
bOUA6j6DZYvBIRfDWF07o0eN56FOoPv03fmil9LYJ+ZD6Ia3lbb7STNI40uSuqyA
v4uyOpYCcMjerKgnywSpn6agqZ/5Aso/ulLLx6Ut+pnjvS7iTqf8YIeMmFObJA8U
xziHfZMElKRgMGsnQ6UmaYj1qWiyIiZ2Mm0TQwJlsr9StugcHDUxuGO9xuLMQ975
4i4KqFAZm+HOLPLjcNlHjObPp2buLGUGlEWtIe3gqprSyDFkzHSSa+nkB8cgmFvm
oAbG+9FOVOxYmw11yMn96MjdlkE3QO/U7Pjtd77IHhJwXTD8ngQ88nAmki7qAtQX
++7Ptt5I3wQ70lbyKWGYVPb2rZp1aLed7b/T9jsvXbWd8b7appSsOIcFSrmxMYOf
8H29ZPQLLnpS9TB+xJurLfJ/gVsAKnU2bIwbC2AYr/BhgP8Y1sMCin7xy0V6z129
48DuxOee/C5xhQAnBRF/lOPtYxoZx7DA+eMI/spF6OBk51pE5Hc7myLQqZPIWLf1
mR6YderyGaD8iTxHA7LFB5NPqeeV2E+tDTGeoC1U+w7XEtg1PhCSYnYWKQwxZbCN
AyajxGcjEkz3kRB5L9ejCMfgO5eHi7oJQAOWIDXFpMzWjyDKx0MdMjd0rQ3SCb8I
OC/pcHanFNyIPLh2KjRz0DyCubE15a8+lvlqyWUbmHJGkHNdLg1eWrxGHB+M6yv1
Tp0IGn2mZpdcYG0C9wsONQ9zIkmEJYIOLmoWanConjZKoj3m6mb3GNafXB/Myy/e
IyLU7vwt0raVa5LYT1RdppiCa4ZomVb5daLx5lZk504QeXHv88c2EpN6g1H1e/lH
m1jpn0dPk8vedMuVL1aJPfLpqQ6n/ujyxw1QiUGRipkBL+OS8ayZI+3lM5THO1SS
/aZ0p9R2eGCPTYk5mYuFmkS4ETFSOYgrjgfzlmDbZsQial8F+mVG2nC3B9dME2w/
QLFHXal0iSn5/8nc1RTGbPv/YoHv7AR6nXLpMttV0FDFmCfrVmOCmXXK0gSegS9P
onkV9GaiothWf2VMNdj5mefK/fWcyTuyrwXQFMYRvupef40Utti+IhX2CidNg442
ndzk491b3mPRd/eQFjzZAZ5Up+/JQGWDBVVAv8E0sh+YdlEet1eOu+u009QxTEMf
1DMiOx1tvmlkjnw0daDJWW/v+UiCRO73ghNUkFXsocKmE1JVxemviYNWVU2dGe3w
seNY5ogHVPekqNWGenN2GPT8BWbOCThVElEFIVKQkZHK83feRVkq8ALLdeH2IiE3
mySn5T1nUjLN1WC9MAd7KTB8vUNlVrjrRjtItqCQiP4yQUd5jFe7hku93Gxf+anI
MIUXPp/Up5wuW0PgMTwzbyAzzygWzea9ZDnYrJar4V2vNCSzvWrmZ9P7hZQ5z7bN
c/obz3EZCC85PS6LTnoTmq19btOHhZ9WAlIANiFJXD8innQIcTxeohprTFK6Qm3Q
j6H1DSnNxed5JrRjB5PgS8AGec/KYVu7ebNs2LUKSAuHppmN4RjNNspKJ1iKZ95x
3IxL0jA6pLEXyEMhGH6GwxEommd+sCAnxujSNBePBw3bPllhk7dW0oUU+fkpZzYo
mBpfOOTLYFPOkRVtoPXsSEWiI2hVnPeTjcNvHu9YhfEd7Cm7ySvEEy6i8RwsJUeD
eL2jUkJFXlwAu/7ZPv3dXTiWVW4cDYnI3X1wsQrUWfpcw+WgJBNy0QnahPYepZy2
zYfTlMZyKc+h4alqBKI6NmlstoVrRWeU3Q3OL2hz28qHitVHz9LwO8IniCIO+bak
A1pHZJlWT0YknqLYtFMa/OeAeCtFKHLNy5mtG430B86VvLPjsSEZs7lhbFIWCPrp
hxbipXCYNDtQhA3ugq+MTaxkg9tx7199G/srPpnaRWHnA55aIcaknkfbf7ppzDjs
hCs7h1vTQmlK1ZX7whp/EWNUWpe6/n2vSdUsjVKZmk+mo3496rRS4xHwKh/dhEnn
yqLgWJB43FY2kzMcGbUKQzBo1zlwk+UqX0QwQT2EasP0Ge+ukZFLbdkcCxco9oTN
BERSXFqeFd09pSOvLZUI0FA+e6Gc/GYiaRoZzOss+X/N9YyThCMTFtgxFbiqZkzn
A19i9fYliL7oS/SXnHTh5PCsFFTFj72KVER4f7xU93D7Z0lj9vcqqwbXkDSPxT8o
2ymqpskRBVUtRi7/FWU1VijCuRQOAfNtB9JBf4pyHz+p5HXLGxL1Ic0Mn0d3PY9g
QqLanC8lLvvOe9RuV7xCrF+JpozEE25thDrQb+/jr60w4TkKKcm6M6S/79tZGv7y
a4SLJ4lSh21HD1poCaFap/UN0NT7pp/Cd9xO8JOIJsDoyPU7gRYv+HWsYCn0Ta9z
f7mUgBTyvrwoL2IcTZkcwsn4QA3YYVPY+v8NWUvhBhAp7WukutNWZFK1IlBRTeAe
tvXftV7hyd+IbRHZ6SEaxmC4GsKlyVc2M1qBbAv6Wxz2686LT88xiwB5QID7LAzt
oUkIsCFubiSNHZY+6SfbFChusa5UVA8KlkR3jyRCEhsHJfHiRUqgx5YngjFhGxMN
6Jcol6U0Se+e2r8RMcByVGawU4qdON0A6RWci9/x5WAs6GtTq4y+Sc9sOgb2DsH9
HeXqdWBQIlm/GZ9W0XTH8uLVxFDitadIc2X8Bz/qe1meq70Fnx7Qjp4NAXtpuWbR
90Z9RYXEWicYS38rHRdXOFIwqdHo7Dt3M3YaVUNflJLCWcFZA1CmKpjpcMJUAsOo
0CxxYCECkntiFAVyywX09GvL/v7luYwNr1TL8kOzycOg1ImVC4tE0LRZV6b0PZyA
cd+FNHDOq1eCQKC1cJlgg9u8Y3Emu6DI8XJ+UYjqcaTSns/NiAHz6Px33VWkNYh7
xfaU/8hAj0WXviH6T4kwLzLUlucX0xrXuV+3Am3JmPk9PqDFY/miz7OpRMOYibFX
snqXJ3Gq5ASV2tvcmiv2s5WvkntuQA+FjJw1FvrYxwrOW93tpfYpImj6OHHG58wE
YgxAyr+ZhHtFe7q7VrdYTorYQae6/hIp0kCCBAcoJ2PME1lYRPcIUZkQCN+iDDkB
+PKkucZrHDJkOADepEwD5wZL0zRq1QemiQJWm6f7IksFIOs0cQn3h+n3scTIbHj2
O/co8Y1d9H1cH7OypSD+mEF8I/XLrJaFgQxVukbkxTQfoIa4bTBTbjsLYKhmwLcl
Ln0N6YoqhTCtQb0C8nW1Vu/gRocVsJDHrm4UdaxhjbdDG4k8Q0psgX76cqrcpQ2c
H038X6hZRd8+pI+nsa8fNUIy2y4FxFlqTxBnlU9AgQ8SAhm54PwMLa1+zr4y4mI7
p/6TDhS80ly9IxUcps/5m+UWuVFoyQvWpMCHEvzkADzJRd7j/W+mEeLTXgvmUI+j
EGDf/qogQm0eyZgiY2hLedsihRJLvsrftlAkc9PGmSpWvQJfKeGR2LeDkxUvuJdP
YOJQlc0NH+hK4MHF8KXTAb5ucKA5qiQoZ+XjJnBdzxv0ZApTe6Kx78HMhNGOoLBE
bWr2Ca2tKNsIOhNuhsMVhTbqCxesaQslp9zl9xqzgHi6k/VzRgNIb2/DaqXTQ1ri
xAhhurA5xQxUx2eTUwjc9Q0zET528RPRiWMVqEkROrG2VPKxAxMscxzXpuUbts3u
JSoTUQmdqO5V7Rl+hY620qe61AAc9GIgYhc5Vofm0PnAilpKa+jwV7+Pefh7aC1R
5dMh9ohqbyaWyNGnEK2dW9itKDCHC2wU0H0Fo1asVbiETZtf8drji6VUdFLYTOfA
mD6XdtQzdQ0CigolQsf6omYQk+JT4tEsBkTv/GtHR1p0XZ/5V4bRg22NcjFPjyyO
dBxqXOnEAK/BrKhOpLZ1sG3KQuW/2c7ivovrMSc4gbbqXAh4+MpkZnfN7deY7Kvq
iQX9AU89pQIM1Bpd9PjxCqpXlo/niYOwodX1JR7FQWeorpHrRjCiMU36hOnZHo+M
bBsl8Om5hA0filZeg0QNhQlXRMR9vwInuqAgdzOb49i5m6s0dc64j0PGmQ0ogsTe
RsFG4/adJJFnoXiFjwDBpNCtKl1PrCOfGZ6+3WKWwtSwulh6gSWgyRuZxq1cmnlz
dWxEEnefpbeC6iOKarvgHWfeIlFXuwMGdImofWnWJ7WrBRb4QJNTjGmLpM/13L4P
RcEKvbHr+bDCxuS+bzB1zkeuX+3iXbyWklUpBr66wsHt1MHyDF8wNsV1/IEFBcLq
TcWehKhCxoXIwm3j+in6pYULYIhcVADfjUPAFmtXi/ssPGD4UKNStZ/pfiQgdG+A
sv98nwwsmwmZcaS3GqxgfEqazSdbh4iUI67T2uAGWDm54iSg3uLXlH1thJF4xqO1
XLlQVm42XQILi2wZbT4xwNc+7Brvu8m9QD2c4y08hTbdrwB1fFMZT9TjKgW/Dsg8
M8e2Wabtr9T+Gx5KknPhEhVkWVhaLDjLkv/se+ctI/H6gh16y3mhsANlqyA3Gk2z
T4h2CV9JC3ZceLwRc/i9TfSJ32TxakYYzL8Nfe21S8Jz611uQj6EfH5VMr7acpl8
ZAPnnPUL4OQ85IXgu8K74Q8Y15pOcHX5Clxy6sSrej19unjQ4woUpTMXHcDSYOIM
JJP+oqkLmyMXpcnUBF7mFhopVCmwBnbj78TqIs/LdoRHq2gPBmxpG2d14XA+kjh1
VlaWNDdtG/H9rup6cLHQWcCtUWyFTWZHTVi8qk6oPxuzjrvA2ScGTyidHYaO7P0+
Wz7oNXwCvxCi9C0xpXjQMaD8a9QGMGOLVAe6oxLTcAye66UE5NOcLNG2gUu4YRvU
wYH9YNfo03bURUajnMM93MRscSo0XRVndHwj79YrCKwnBj+GebV6DH6DUJ10UDHl
ZIid/y5aYVnzZ+geLkOohLVBF3afq4N93kMWIWJiOVmlh69tap/yrCZRdU2c4/F3
19qm2onKCmBmibstIf3tftgkPRKsFoSDW8z0haTjXgZWSGfCu/BiZ4CSk1RZdGkd
9gEyGOy2H+kzROkTw0nKrS0Nc4aOgta9654S9a/lVWWr25oy3kjH6t/hpIbXK8nj
kS2eiKN7Xaj+8vspGsHsCYuKKlUulmrOUiMrtsPET4c8Af4vEbuZmRQWnkWmwZFo
Vqo8vG/IiNcVHPr5sh43w4Danj2j8+MfLnrK3r9HB84HbQkONhAUYnfto2ARoW7z
wwSiCsjVZ0DK91R5uI+lDfCutx6cEmSWXW0+ZRvLfJrKdMGBO1lyrSVi+oBpvwYd
6etghkn8SjHCbJAkL+wglvatFMGCLsRgYDRfzW0zGyKxhvPXrAUHnyz1H5bywrkg
EXzK5UkFJSWew1K2na1qiUAe6jAQR8mdXtJYRDHnw16BZZk4v+a5i1G0lv0CJbdB
YoN4Tk1iP4jgCIHZJRPQLfMVLVS+4ogyxYrTJL9rOzPw6BB2uoV+CwRI2VxYj1No
dDvrE/TYmU02d3TDe+tAe+fII/xgMwUp7YIiWlKWjJ0zI0wvLq8C6RguU/lfG2GU
6/NkSjqDA1oNaOE0eOrqdlQ7IKkItdb9hD9ikOlA6utXFJfxkgHcgfxvjU16kIh8
Ep4ROa7fwRNfgh3myHgjflaZsGclQ7DuOagiG2thIxrPg6u1TGKjcQx2jZmCsN16
OQCBLdlRQa4WDj9v9+C4IWwqmuKyi8+ZpvxqlIl66M1YOJpx4Lzc9gRQAJ7P/z+d
WBwXaFuURqEcpGYWYn9Ql87AC1TytK8aNO2fpF0A+ZmjCIYhIJXhNVebNuE6SHav
XfRsKlrKtgNPFQwuQHyuA0X6eP7eAXigWsjmkxCvtC7BsX54Fa/Z6+HvkCtst4+q
o5JUsDuT+cCKguQu8+9mSf4l1GrJqH3ICbsEzbxPbn6Rqs9O9DXeePBe3WfVFzA2
v5PK2Z+k6wdjU8e3ylpWiyKsUdu8letYq1f4lTSRt9EF37S8GQAv/O21jV5qvex1
i28pc1uWQpcGCRvsQTJV4mcZwUcLPrkjaLFbIuNv7DpPmT01u82QCVNBS98F4o9L
och9BKCSuXDcPK075ATtLX7KzbUU/BdEjUgAAshxLySna1CkIOjmSGCNu23VS/Xe
UoCtES9ZL7scc0yWLnkf0HryFOlXiYmrQTHMK81uOkEhIXaQRpfyydtVuNnS5ssP
9LzNkmDiveMcn7BO2IEw8sxfxG070OP75KEXxWkSE8EbQ4PeV3PmsvfIoRhAVd7b
LuEmuC48YW8I8lnA/awAnyUc98IgOo36Uxhzh6821E4PVOiXYACDLhLKmra5RvZA
aChfgasinioPq/GJVf25T3hnW6BmADESGMtf6LwW8KgSZUV4l1YCRPiQ5unwLeKh
7iXHzVvzUU0Vm21eP7m9EJSnyZjm2Usz5oSY3sbrUSwGn/7zgOejEqGxo2tbPuZj
Lk8jJ438N6m9LB7TvzkOv+81MGMytAf+d/1/PomAL92Wq0glfv4J8GpT0YHtwY8U
Eg6shyXp6DJUsnwbOE9YdouIHyPTnOZ3BuTfEUnXWM2Jqw16M8jiAE15W2+w6ifc
6TPt4/CeQdF+dklgo8UQB8LOB1Mgtteoe4jACo6B/SBVyywdRVl+GfF6lU5hK7+W
PyVEFzvZu/r3a+mgcKfKzXhj5IGiCrdUTqy4PRTiN8sZL6RO6BdX6YujMqgbcbsk
NsULDENv8rrXFYrTXL4ORB8t3ZFx0dyPQqxF7rUpUae+cYuCH4I0Cy1Akx9w4Gd1
F9X2c5so/ZEKK6HyMoI7UJ+iGpLVwQDQVHB2rG8jFPBG05g6tGsyFJN/n6vaO2C5
3whzfSFMqiDh8po0rkEfJX2L+Kl9+B6E7Hvwpx54nj8nNNSn3Xk0oOMrAcbk53A3
SeaUHD7aImAjN6Om1aNuk0k272NBBoN+8/ZKJ9QmMzl8hkjhUENpBuK7VY2RO14V
YBPYpe9LJ1gZ3ys08ORB9e3iNZkPffvrLJs1FVhqvU5ZXucQMX8m9cOFu6NW3v7w
01N556vs/pKg+oGM5GPrrP+MHFLPaeJZu8V6XjO9PWg+iFnD8C63yoi+4Cet24La
+NXIYCGZeDmEEhoEmXpBViyfbKrgDkekeAnjgeO12bKd22L3FZK8O1zwLqPg3wR4
yfD5pM7dJkc0eSnhEBFDMnOi9MAKykMK3qq45jddfC4J44pk7OD1gh0r6mWn0lwA
5rSHD4YuZbllId2lJGrrP4oSVRAav8EzbQfTDmqbAsHQS2mOmY/nGhssh3Ia12gb
TnmcGKsbCDRkN9+9DxjPUbazFyg7bhUKO1WJJvYHWuix79pSy0hjS4M2tUE/1CZc
LHmSfTRMzm+JmPbbICTAzYADpJfhfUeEBDir2GhrgXla/R/Wv8qu/ur1Q+2z29HT
ID/59HH2QN+oCiYp9Xr//W1loXvxCWb+yfU95HmrBxRsZ+LOxCjTix74IOiXmUYI
sjJWUM48m0MwlS6BaB4ni81X0PX3QRD2DZ15UTvbPqbSLzGM53N8Dn0Lb3xBavRi
BBSj3pPIiGpd7idvUHIVsGQOJcjGNU2LuJ3YOMk29pc68tIPti/CMPlBrNA/4qjO
Z5rU2bPbrWByZasdnU938i4w2vuygqxL66EavJINpwfrIfgt2TOTmEdpWCWTN7e3
aFHTqdw0kZe5kEQkaPJkq0um/D7IcxEK6fnt71WWq18EeGcwuT6OB+51df6eFAJI
QALaSKIbeXRK20KxZ2RAh/cNPQCSGATi3gUrJDqjpghW1bGLzQp6EVfAzf6sCmOk
3XkszhURgeNEsFoZCyfu0CjNntxSPcKI6u6NDyFj6548HoLgPRn4FMacFX4h1Cy0
Np198DfIH2Zkt53KZmxVT76XsZsMX9MpYsg2NodpA5uWhEJ4x47vc68txDCqudel
8MwfaiVhqmsILTlQC7HX1dL18rI7TeZvQOkzEWcA+lbqYS7CeM00Fp8cug+Zs4oR
trDtMS7j1YtLTieQp6PYYtHE03+eDts5au+pI22Cgp9w3HI0dcJLAc7Gmd+YQqWS
IYQTh8jriToCTKDjAkLbgEGOmVHbCa+ZNKprNOHyhRERLj04H1XLFnmJSN7g3cIl
gH/mlTQbh0GDyiUOZQ6Xg7cWTtlOfWFI35YlJ8rCZJXm0Jx4LXb/49ujF+oU6xRh
WG7UkOBH/mLwOI3W4X8v6+uN2kRSRsZ3iC0HJtVRp8c7WfJSEd/3hlUFNjy8lpIi
0/14Dfr8kmGJA3ZTl2DRLfy5B+vAPuG8Y0S2lvNcuiv2cOngHZanSol+zLauKg2V
Y0iK7v/TXfo70d+QMvh+383mkLJ7EKhp5rDjpihBaU2DQYO3CytMde6xs31pIP9v
r4MIkiaSybHV0ZLfmupHtLXkkDI3pKY5RK1MJzRKQoLyiCppwPeEip6zQfvMb1LW
1Z8u5RBbDnRTLoDbvUMUCyfmI9xQ2e5tEVHzxNQ+MNJiBg5xx7OMCAHzpC6m2H+8
LuV72SvRC/279N3GSrQoiSEEVDlKWy8IOly0ZkUZIjQ1tzaLLQTMQzZggOJ+5a0X
EHk9PSJfNA10Sp4nApezH3MfI2E9lR/hWbDZ4xpk1xyfsou18/FRBVmFgLgZ0+lK
61SSLzJms8dk1eh0uJ2WkMfeZEooY27+RIDHxIkHu7An+xjjg07oRroEtn+zfOkh
OZ3ShDP7uNvZHio/ugOTZBU6F6f8tMYrbDT5jrz+60gMVYOsv4JVx9GJn6F3jnhq
3WMHb1JTCbfA5r0A1qt4Nkd7pD1PzpdC7MeO04RjGjWp2hY5crskKCXvcC5Y1kiQ
j6ljFLnFJ87/BlQCpXRTDsrGMQIqb0JCwfjvtG0EXKG+d/jYYc0Q9PmoIiqwihLq
5rlNqmYpBhpdNhO1fvHvD9nahN3325CwwvjDNoh2vFJCKqckywG5cj3bmbE9u+dd
NTIqc48vIuICTmD57zBLBFoU/HsiUDwGdIZ2kaUP5sQR+g1uoRtOGN2YZq0aoLN+
4ZPa4osJ06xVegAbVpL8uU4S3MU05q9qzR6anRmvqFa0xGC+jN3Nxa9U8o7bpjtC
dut0h6VVkoJlbDG2efF+kGpvpWGyY+nLKlss6L1ifu0dedE0zmckGDcvs1F6zxDT
uy6lfHtTDAooMXYBafAXzZfBJLevTkAhLyBOQntbaLry0ajfYHq+Iwqh2TvBiNcc
LVPAWdtWRmKxxC/MBWC+u6ORroFmfFREMw0tu/GWffvax03uZevvh+U1xOqdDIq8
zFgpMNjrLtFkeK7VokDeMMouuU5mXHZfFbTBWlmqlPdo07nssqDixkRRtICWZ0GW
9Rq6UDnc599AZmQP9MPwIRg1EWkTVuau+ugqAisS9lXGSl3Z+5KqK+VMHZAcTDDy
cQ0iYvOTz867pRaQlS4ZT7FNbA8y4m6CDTnFlDjXiEuY5IgGOP4XA5yUXaDn1rs8
wWeiFFySXZGEoTQOYWg2n+D8WJXBY4Fhg8jiLqio92/1rPe0x9zpJ2Io9tAhsxG+
9iKomaWO8ThpGoGPKAyyzA/HMDbDVqLOYt/MhhaskanA1OlGelNpg1wBazCklsOz
3VywH6nnrYg/G6VKUTvWpIkzBfWknbjm1gMuZRlXDxQste0YivVs6CmDvIpf+wGS
rZPsuZrTSpt88zCrbqpI0ui1+1YQtqEv1M9P5+vH7eYhi/j79+lDmvbzXR3BNYAm
93X6HTheKkZzcJSlypv2sYQW+g5K0tWxeU1af+ezP+Z5meYuvgtk/gGPmATjhwdk
w+z3ArW2fF9VZORqORiop6wy8Mf6WPP3MFCLX4ZIiPg9/8Fw7P1h4VmwyPcBhF40
iEpNXELsY5hqOMd5QaLRNi17kvzUYepjGnRgX9mjWQV8nbQd/TZqjnsCZs6pCI93
fm5Gd7KU9DJ7bDmRQ/20kNAu00zLdOn0VHkexEW88aPneUaaddRvVi1vV8xDLy/a
T3NFB9ktelSNz61lmRrriy9+mFLZeuipXspKn/YTcNb9DFSGD/AA4cRo0ztANqQZ
D6sw5kYp7FjRwj4uqxwHu7Gnc3n5XnQ6oWomIAIMVKTql1w598AzqV67MV47VRCO
Dc0Rt5WmOrX/qzto9CzIOSzzin/VADT0IwR/SKzUDf7/LJvHh69VwjPP7ULG3W7s
OJzANVTkn7xK6VrjcUsEN1BqriDjCoT1FVf95zfv/EtUJmQVy7o/EYBs+TQ8eM6d
7rpfSul2jx1zYcp0u6fP2r90tqm4YCex92txnsoN6I0S64bYvG0CYY9Nv+IBujEB
mWLoF3kfZJ3LIWBXJCK1iYUzUhd6nl48X7j3k3Tkhz2pa07fCNibqOVYROoNG87S
wXv45EQhkD52+OUiQ85iMwQ3rNy0isd0IzkWlP8ko8OoL5xdmNmE8o6/LxVz2RfF
cPwyOaY+/8ACUSqlT+4ijFThyjmqwItZG+KQ6uwISmSTAJfXlU/iV9gh9dl7Y4cq
bvF1yFHXWX1ZG2I+qdj4Scbp0iqggFllvchnSYGSnZtgQlSnVJcuj9iAvxBzgHoL
+pSo9GHAk+iCbIc7wEZXbWWeeL2lwkyxRb6DcFfLVpq7uQ9LFeAysv5wXQ13ksBR
omEJm+Q2d8274hNhydO2lwGzJl4Wz1qI0qnCDEUJ+FgL0CEQrJVHlWLIiXsRRB4S
/aqHGzXP3o/MstpfdUvdk1+ARPAdX2ud8YzFICS8raBfzSya4MeYPESTARC8C8EZ
tFDkwx3AngFAl2KYPiYj29jZiHDp9lUcTxkX4YKbCO3uVi6TFzzlaS7HYRUNQ2zW
Bprqq6BjubUvhJmb/auAtF7ZnGA+klTmK99R1eIAI8I4Au1LqnTi0ep0S3OfU3xn
8+tUmj8l/IDgWA6QB2oFnV3aGqpweeXbYAIc00OgNKg2pbvb7YpWb+r8k41f4rz0
DHdOyRIUSlCD+LV2jgR2pDN2l/YJ764v8rYUzUvnLrjuIC/dQhbsFeavEvo9E+XR
L2JLIHhbGdbmPqVlo8qRclLRxKCGpF4nH4n0fFPERC4b0cusxAQo69IzypsgERyu
SalqOhA9wgyRCUVE1vJ2Cr4EKqjgb5ycU/cuy6ov9T96OxIbV0jvF+aF59lz3YzC
+FWcaVlSXSm2nPQ/UvASsaa+vib+qNnCIEcvpIZQXQ2g7ZLhgoUEMgK6+FV/GPP/
4wN8dPMRTXuWAmvWxw1TDUDBtTs3RXx5LkS/H+RXE4wjg9CcLGvA8zlaQPJnq0x3
Pb2KsKpJh06big4T7rbNHL0QsDMGAVrLBIqaM9wuy0FqndLerEfh1G37w0ZWeZ5J
LkjvNWQyoiSfZb3N9gBuljt89kK7TUQ9Jfy7oojbdR0w7lCg5aQsu/dKFR/SYOFt
zFdEohMFxC2Hdq2NsnXluSCAYyzYCIclHsbg7HuPYqrQaB0O4R53i9VT4CMep6Wo
9AFkfIBDnUrUy9caCMwwujlVxujVa8VT9S6pKZN9o7D5xWW0ghI9ajLb5LgutqCX
HOnZBNWLcKOw1ok/i4lvNHLWyRh+nfrLYkL7LRllc46sZEs2HamLmZRJYmTsaEj8
bc3/gpoKUf4Xs4+XKLqO5br7i3ol8tzhx6ULm0RaCCJgzd7EM6DDxS//1yiNtk3X
7leznOAY+n5S2gIhw3vxOjIycZXe2cEBs1cCCkrFc/VSeOht4Ti9MPL86yh2703Q
BgA1V4Y0M8CYLzVWkPV1MGVjpAyoYAdrnSg8q40vgV190GVUC5zAahVH+67bcHJS
lv+LrSpc8owTByaKO1grErFcOL+3LUAhNZBDWmg/PucUXcEBtYytaBzH7WI+UrOt
L1sJQTtmaNUH1+nIk9zx8izhdYKtkrcytBxmKHnBU1hH1RQRLDjSIXTaNCx74nlu
I2k2JzeA5KOsuLZW/QxFjCK1d58V0RuvnFIwd7JwqwET6vv/UuwY+eLgAUfI3UbD
8vA/H4i9Fu5WaqIt/Nii0czJTYXvPFF2svjCRGjhyt/aV8zoqrlD9CoFgWa7BnAC
eQXWSH8mrxuvAQidlHSEIQCAYuYCLrMimlF9SGcDoKUn6KhDFyKLm/FDn0HVY5EE
WTW2Qas1qjQPx5O6SlSoSz/T9Xq9deNY/d2sF3jGE1VmzKDw8xSCZNTKDiaXMUVf
H4q+s5NumYGm/t8DzFKchUbQKQ4JVEV3jtf/GSiWmz0gmEjj7DfekdKWNKfyP/91
pjbwLuj8v+JzmnGoMrIQ1P1bg1cIF5cjth4nrv/rbo8fKZBIqiPq6Oj9Y/MCf0nz
DKirzd1EdYdGgmR+53vvCs0AbqrIgbk1IFjfZf9ZR9gLXB7xPv1JgGNKje2xybk0
5u8yFl7csxUjT15u8vslRBKpx2dThkiJo1gRcMs52FB9Ck6m8FllnuLbmeCBQPUc
cJN2cUcd2KKBDjrg5OfvEGMtYwbLD63BG7G5ldqaIYNB0TZkQhtGzZCnjsBvEVQh
g+i2gVwGvlSGzJONFw2u7kVfw9ZbeNISPN4tQaqsES00jYJFX7ghvqXLvoUrrFyu
5XmhWW4QnKAq0yCAq2RJK6JvaqBGZzZNfW85VG+rBoOKduF1BohHcdTeAKzy5R24
3drO06s8dtu0D9O+1CGnMWjExnWzbDG7Zd02XQjRHHT5lxSHXc5foP6guq2uTmjn
H/qON9mWXlVdTZxqERzkeLJL4X03PfTtq5yNhe1lUai17HT5yzTRYnbCCoHBbbvT
I+mJUnbXWddgkwBtwmKghB2BNAg4t6iB+3j9WsJLbXK1alsG1CbgSGJsfSC2RZu9
dKn4VcMlUw9z0FjM+VJ0mJh8CTGF2zWxLfBY8OnIp/hajD20vV61DKsOyhk1FJnE
oalZsaH4Ibysm8owp9HwYT2lVcVV27B5XhUjttmmMtT+yW4v/J9MVQmtNMZ0Hby8
/hvNWOPmF/lyzi7bBOgsFnFWuO9cK5VmnYgi2IQ0U2dojgY2bf/ytkgVjn9/4u6z
Ko5xUiwKZ4lc8sFan5xh1zjFm2veU3jKX75KDZKv75NF77Sw6xd4yjccglGwV7h+
W1b/ZBvAVULrjpah5vYKrc0e4UV+DJKzLnwKpzFhEUO4d594TjdrwV92OVxGFDry
3pEau200E819gKsOjDN1LT540sNne/EZIdUmCJc9xwZ58XdUkP4jxCCJ7Tw+IzHA
N1i62MNcIWuBFLZTrII7YiYsEbM+XwfZTFWmwkOKv2VqKxGhWNTtB+InHEsE4nyU
GKq3bPlXFRmxvJHE9E5yeeOZzue9+MSayq9BkfnSbmlRYsdPkPTtG61CkmbIAZlj
EBkb6VUU1yrRY+B2okCMeJehs7w2FYTCDzy5G3FAlvk+jjZ0DaOiMjGK6yqhDztn
G0ru2k+DGvSVLBHpI4hnKAAcaF3AbhVaIe9Ggb1kSIDWuurm4OPekdfHQGSKEqco
vaY4X+tChdahxlNqr7V99FOybV1AksBe8RMWLErhMbCxIcDC7fIH7XqYBIS1NsWY
+2iEbjRSVGHQVQSjkhQRoecj9UpGEHfR0HURQLSlYieZ0IH7dbWrqg+dER2SH4Yp
lD5AQqJSd/rodqULsMA5cP2He5yf1C8mdZcxdlRZ+NbcGgCEolxYhsN8RIiCInvb
1rZy2uhBZPnCqZCbZYEvTvkVDHAzZtF+AzD4Vw9k3AQJ8eL0T0QqhLC+/3l/6it9
zA6wn7b+1b0ASnVCBPObeG+y2YyKAky3dZuMSKy6nDl8SMNCjMdIjX7z5wKcp6Ek
CAzfgrf8squaU0bAROzbILOl3CqMc6HzUBnhjcjSNMPM0OQxGEWDlqwqOukMeyaL
agnb1zEA4MzkrfmTl+59hYyjGsx68lZgCzWafApPCZzOKh0cuaOueoqnAZqrQK1z
PeGsC5UfWYLU28AlNK0Oc+2LgvDq89dQXY/hvStTZ/cj8/Z0/rrYo35HOWagUNgq
y+naqxHpfyNc+bnqgd3Xz9cmuN2BgJos0MklXlG9mCLLzYD6tUT349xJiL82cinF
QESkJIsx1QAQ5x+0v4Xl+N2JZhLOWYO81W0gk8WIJwGpNYhBohaEcmBqrVdbXOXN
l6fO2dQv9JTz5CjZnzL8wYZ9qx+1V7z/iL27KB1/aYuFQFk/4xgkteoiILGottXF
fL3SScsXjrnQidUaDI5n2TbUEkSEoJcQeirc+3oaBZqRnRk/1CliR+vax8xkR4Gz
ebmqUS3QJS9uh5dP7yV1zi0Vsmbnt/plg0bMG3Q0k+zSQU3IcZFVnSfX0GH3NTVs
tjeuclViULoRFMFUECrUavnWGsbCWCNHPgxlcc9m7Utsu7plecR0ad3BpH9GzHDr
k4K4chAkqqP+1uLFYrC96wxZdsRzNeDrRth+rAIJlPmpi4x3LBkxUB730CPP9mFV
Ildtr8kE4kXEHnnNrNdjT3a1zr+UxnJlapFr0QFF630VEU3Z0KzRmoWXTRQRRz3e
Bxq2Fw21RnkeRK8PAOZJ6O6l4EWPB4GU36csUDrEOd1El34tgg/5WjcM3xzjBKNt
r8fd3xPK6ybapdlzm8hPQ5Kt68I3jzkYEnBTRHCcjakyX8lD97sscKK3OHe8d1tJ
1j/K0a6fxI0KuVtD7zL7WIurSESnCP0aqaM+luNW7uDyWm3FMq30lvP05MDvzdH5
J4qvo8v35U92MN3tzjLug5yJL9lPF4bNjupxpN51DccVkDnzZNTX1k2/c6Tydnyk
JDQRMebR0r6a1SPhVSh7iHxIHlV8uRhA9MNifBLpwfdPXimIaZm0pca8GFp1B6B+
dwEV2B6K5VpF3IF1uaRb8dkvPaXRqroSVVatSthll+zv2N95xLp5d3QSMgOBFcYo
2sb3UCQzHcPUbuYWPyAOuzb1n0EnmB/YX+z2XGoO8Amt1RQDScJ/ui3jB2WeCg7j
X2FghQZAxTpgicN952usHeINCszMdhxnzxWRIN8GnEl3ifhIblR0nrZPd67DTR78
2YSexJkG6C8NwyPx3orzR8io2sqAKHuVIhUtP4pQSSGhNSgXLo6o6+VCIHn+7ZaN
FW8IVcXi3cRlmkmHZVkWekOuGEJvMjJrFaAUj8cJ02PCCFnmv99hbFzjQQA7T0o8
QWnChvMqUg6DiqkZy9BQ6fgAEqVJfs4wDp3fbUm0knRrDQwDgf/B3TIfe0rXXYIw
wPVKzY+s86twf0XUXqvwXsoU+l09VpqvY6qha3i5wx57BMD1eJe8TA+rf8uT/C5g
VJ6nszVEzN6IGSxsIpb8bPKCwxbQ4CcayQs6z40AQtFDmftU09YfM2vfY/myExwe
HK9kHfTGZjiMpDZmUUoJGCp1nlxdorNQ3DigN8k9XpbMdn7bSaebz0pkt88DRT4s
SuLdQnIt+3jhI5IdrQlDDH7E+t5EGd48tTQiRzk5kmnalSRwsW9NDvOREOkMEEpW
wi/GIAPfhIgdmz1pKnqnK/fFK/wlXwzqetbxfpvYqLc8n9z5RO9e4f9DhH8QLRDQ
II9tyYelqeFsj0VzxIE0QrUxp6qqMz0epwH2O9+BKv4NZ/sUz3CnSdv9vTaUv8xY
2/rLRW2q3BSbdjMHkEk55onXHUY+f1RK5KY5mfr7Gmh1cVz+D8CMLy7UIEOBms8+
NiyjMuX8DAiEG/O4+lzPl2wkM4rY8WJpp48EC6Q/KXgbQky0sMeMJth4C4JWgqsB
xlqvd+An2dHcB1OvwFYS0+vkyUcKpB+afajla96HZ+6SLgm+aKX2sGp6Y93z6WLL
g0Ind2eT7NBBOduVVOtKLxQdikoTAMpnM27tBF8K8mYa9blIMfQp7Hhdk1SmOniw
51gIbixwsGSIi6YtZpaFM3h5PjmJzISEOCYyIAatito/Vkbo7gmGpat0AzIDu9eI
4hGJp8Irl0uJzPQYVACJy5evwcFXy5hQ2i7wrOaPsS/cR9NXvk8DsN3AtCdWS/UW
zD6hd9deD55jZitHHSAcvfLMUMw+XPsE4TdaKXObTYMvMgKVQaFeqZBdhplX0gDd
Bn8s05pQA1rYYbisNKhNIHhL2Tp4Ersos2reVYNMdudwOgSnhr9QJX2BUJxzywIv
Dtfe7I4oi5jSTpTgRZUyfRONw8kN9R6ZavG3nI59q+P11xF8moyRFdhRhanPeK6D
0XTvKm+RN2h+JxpXUM+98DmTpcXm65nh+qj/kDhGsWq0KknSHIsrthkwlHov46jP
jr+OcGQT1mles/XRSFddrEkd0oI40vwgKv6jCvyJAeKi+vzbUaxAGyO7m8w8jTPQ
exPQYG/46/Pvpz4hliuqeGmc5y4HX/4BI0gbEA/25ex5TXkOgNngs8z01yLOxMGs
DB/X+SlNJ0uNLIsH2F3cqT87D/xO0/jmdUj8jy/ZDJLsY1o1RaRPEBSGp1WjYVSw
OKOK+ofRu7vDxiCwdya1XpducS+/2w2mMDxtIh735cL2uq9AEDrac8Sjw3GTfDFh
8egghcCFQZB0SRgoBsEBzzHEpE7QZxycxScvqkLo6byY/3F5TSESuBUPQuSMq7tG
oWUOtR5kPiQngnuUhYsN9dDlqJv1D/PzZGwdMadXyf4QXl1cFowvbcEIko4deVPr
92Se1+OYonBEM6wXocuc8bxluHBz9I+ueYVtEjo+yFXdJnrNuEfn8Rnk8r6aMoXu
iV/8/AnVE3ae4TQUdDSoZf51HOsgdcdyv4if0Yn1boa65XbevGMy1W3Yilu2wAFz
aKguUTcA+woMBNUkF+AeK+iFcAez0vuai6JtifPJgrWyIbBk6ZHzuugFh0C+FtDN
QlDNAFmVB8D4ZwmMhK8ZQJJ5MUeIu+3cjN7uO+hgHs7Rn7HzFvp/WuUVXsXlBfiD
8Yo/bW0/aycvE64jNHVQTbQ6i1NLvYknmkg7zUEUeY1G1hKM6EgcvP11B3q1hLwU
v6Jb5RIuKphYK5iECvU8T3XbDUlK7+j7rlJ72fjdw2opqc4xHUU0iw41oy0G1ky2
G9tu1tlheKxrnTEBaSwGmRJ2Od9S2LjUXjJsdGVEtRouKpeY3lI/pV0EbYB/wIW7
+jKZ1o8A18ORO1lb7tfUlTjZ3T48vYPbMwRd+dvR8U+s+cw7GjXf7ThUmmvFozNK
IEK3MFgc27neG2QYM0nyzMg5org0JrQUHgFEivFN5iPt0VpD/ZWIYT4ns9YSJyLP
kfxT4uJEzzdUJlY0IVePf3fmpmM2Px0p3NqZG50uhwNLQ7fmJm7YuUUNb6nMDcAw
b1K1b5g3gEeCqsIjkt+JQuIV5haw6/eYAOFM7lDErmAlCgEG48lvW3VHBKxgfONx
IUcMyHdmAmfZWB038cMAfkLPnSx4X1PR79hKBNgRoUdHg2oul+HrWVcJOG4PFcqG
I/xNwgC9yLJAXHNSitxlOZ6U3bRsynSr0SbzR1UsWCDkpYUQoaCWD/kcvUq6glIk
BvtygpDzER1Ep0CuLArDMReJeJRlzA1f48DxQBzrmM2RBotW/YTL/47pNIQzFto8
Ump+tOfzBT3/umBElmETB+H+uIBoHTNtGf63+eNfPQF0iZILtc8s0UApZcR7K6d7
M1kMu6I0NvHLG43tflVxFqMmnFBC81iD3O/9LFICi7yi7PjLacNwhszmDCmlRw6g
pGwkGPG/UZBn3lwkh1gi/zxZ4Lbj72ZkuedmxTWjAAG6/TUuw5XSCgBqOAuXAfIZ
/Lcb6F+Va1sDBq4ZLOtrFNlGrBsNkfbprU1zy5KNUNoqhsHsv95zFciSS+iVvmOC
MuQoPi/01HRZ9FKpS3BM5cMohvghOFloXy1rzO8UboWriQ/jXy+hnjecSVQEYRjp
pQdXAXv2NwYaUWuFIiI/Oym0jKBcsuJb3UBleE/Qz1jovJirijrOJzcF9DtvjfuH
clkFGShH7I4/oXnFQC0wFtq6i2+YfJCffsuq8mB2btxLoR+FTEEwA8nr+qV8arqY
DG5ALE1y740VEXO7f15Yg00EcrcFwvUfQDXd2HidFe8DfFZP25PBYqWufMG2qamt
UkrLd1M3A8kKcc7RQKdyHS6xqZMSRwvYEzfnGUMIRveoekXT02pb+b703R0DjwvI
k8DvWxEwAI7FZyZk+wWRAKb+LdsCTEe3iEm+/5if4bSAvdCdMiIPMeKJGWmv1llu
qgnEwFZXb76GxmVHOISyxMX789Cmw7I+eyZFte9jnRkWgEjIE87dVICZQ6H3+xwd
dgJuur8VJHZVVuMbTZigUyLd1H7wFpdhAcS5JRuGUGLhwLuK/TdEMfqUjc8nrerS
mj8IfDePfqJXB6SgrjJg7MsZRZzd4EFnvv6FJZOvTltS2PCY4ANM4KJ4fJ5uz6r9
jfas3lgrdDyMNx29pA4Al/TxSwaXAlkkp5AoAzQlfX1Ss8RDtFcPAogQ+fGwI1Hc
c+6d65Bzef7KQTQTHNv5kVEONwCO4BSvu1bvtIOr4nk6EADIRpXJP5LMaiOLcK4R
raMSlfCzMZQzhyAebzDcp6OBUcgMb2c5sV203wU3f3uqpl7iLFWDFWTqPb86P0wg
vBFiRen3aQMSNRvKlJHN+k72kvmmlx4v7EdaXWq7PUEfulx0W05oW/TFiip/5CPo
Lz1PPOeSdPM9mjN42tj33yr5VVkPBxgbmwKQxt9skF/Lx79idZ/gdQrNMh5MmmFH
vQl1K3B8LVCaC3Vj7oxnxOI6FoevZHno4Qd9weurJVZtXpcvrVM7sjuviZwgo3Gk
CGIupOy87VZvHRYUiVBK85EWR4+9bwq0EAV+uBcEl94wxTaANdq8qbIEFISdCVBK
kNpxHqbl34wzvNM9JOaYZR1MHlTPMPxbIcPfbpeaI76ihA2k/Q0Eui0LV8rDXPB4
dgCVUFrjVj0/5OTl2qxdGS6nIpSVm6drBHHOJzJXkYPzSAtd8zVHpBJ9lw/g0MDm
2kisQSIDiMYDG3sMc/mV1Hw8uaLJZOmITMJD1xRXy8clCXgNnrgeAJpdf/6ZlWRW
1xDfqJX7alMi5g/yGZ0ntWrjgRk8M3GoAblMbCFtKr+A5zlRakFxbQnHwayklygt
8HNqA008D/KwAgOmeaSj140q4gZr7ye57ztG/cyrjnUou49uLiXSC5af9BxzeTNl
KjtcJYVsfiX3WkQUzpyfQRIFpH2cOcpgPKaaFJTZ1bE/p9lH6gnEO65Ao+352Nhq
26KRsaEMvb/vdumVFiqObbriRUFage9nQUxwlm1VmLxqDfkl+Y8MGg6QN3kEfJ49
Icy/rJkghWOTxAHRua7ql+vFrJmLrEXx2KO9baZOUrdD04lZC6wfGO648zSwUVs5
S0lEMnGJyUyUX2ZAMEGPKgLOLCiTPUGN10HJMMoBXeTg9rCKun87Bg+dd8wYfhPX
qjdIM1h2ZTOybJkOTL6G2rlJYYHK1unFVEZvDXJdAZvcYGFGMgAR0E8kPVWcIDDe
vf82HWjpR7ADJKqCc4y2GqPag0ZZuz51ihlKH/RGj5rn365cF93Pc0kxLG6PoMoo
gzSfCH9M8x6us4VCTUIPx8M0ftlZStk5ov+5jrhN+RB3wHeN5opJTYYuOCNQaTcI
HZxuqTYHviGhs15v4t1SPmbY6f1EgJu0fFhDJGguqz4Q7528jk2jmWd33fkX+O1+
WwN9AyNBZY+/NbHLsQEAjDn8h8TctRyiAfVe8iYFE+Py8y8/G46UscnSGNlnUKjN
lh/5c7mVzv+uN4ia64IBHM5K7cn7K59fFN6xaWAaXePzLIAWCOJ0cLX5LazYyDHF
AxYQbf2dB7Mxt02hVV0tmIcuopeuFY7rW37HkjZJxLGw1eARSXnaU2t2T2LTjbdT
sYYRfUcMig4e44rWw0rldqUColRjtc1VF/BPCxlZFx/wjdmCdnXlRPzQ20PAM8t4
prK+14Jb6OHw7SwvnS9aYzCH/o/QJY7cxkCJTNMGY7hxQ0xW9FuKNZBocBK0w2Ib
oF82GAzvTUqQQI7UKTdJJv9nume0jK4rVqsSznKnjAFfresuAGSENjKn5bjA0KT9
sbmIhwssbylP0klMjpOEUqqknnQdo9zaEBv8frbgKy6jOllM0LBJzUoIUJsTcdl0
t7MR3htPJTsHnKs9jVJFh35CFerkZFVfJ3pTxljXAdjQa3nkzxeMzTm9xfR1LgsS
bST75ol+V681ghyjGQNmAcMl3XGEqKQ4dnCG+ENIsp/G/Oc2q19vdM8cj9aDzWmg
qGEbdS4yIkyxFdplb1t6QU9hogjsVxqnwkM439hozNl0XTwnHzagNzV80mYidM6j
cmHqPC36YeGRX6bL++uPhEdhhHLFwlIcjjMkQbqd2CWhhOkYeV1oCLnIrbVb7aB8
PBF8miX/uxNy9yVaLalVT6131Bu9lTGYXzOe2y3fbIjv4fobM/MuGRToo5Pnk4pY
cj3s1hVlAZvFYW8BYEgNOR/q87ZM5o5M3HZfzxqmp5Bvvym+BTjfaq0DMjcbWfR2
8IBL13WkpuRtlkF7PLD7n0JnVDH741pY+V8nOW4X3+SoIJEhRVaUvpQcumo/Yoj8
v2UNWDnJFpJ36cEHKymvb7eGqQIc6ztH9MOp8nEFcxqV6GV4hd84H2RWiBXLQAqB
RihsPkKYroPZiGVUzAIFz16M/RPTMok/rOncPpg34btjxSIuxCjMlbyiwH/DyMXo
2minFV3xyUS7beAPf57qYJKQVv/s6DT0mzYyyAumfpy7BJGaYBp6/L+D5AXr3mgm
vEf/F3ErqcmJEnewlCcjxb0tL7G87/nFZGOshleptBvTAkH8mcMaushS/Air02fA
o2RWdc5Ahz2yU4eKtGDShWQoSJN1bBaG/8TRXSusu5wyx4YX/GRDmYDSJOL4nQ44
7HYvTiFy1/nUYwD+IxQQY03/EouKfcagnoNc8Dvqsn6uU0OwHrBNzDsejMX4FMKW
ncRZ2a4YOFqnqWpYS20S5FQn21vmH+y8/drohImAbbPRq4TgIn0axXcVDt2a/9oZ
sPPG70QoX2sAo4w1n01xGOrMSGgjBRfS0qERsfVLGZwm+b3khgUF8b3kgRIwsfyF
jLpGHnzFYmWc7reunWvY2D/LSGxObdAeNM9wp9L0CTt34W8nOaLTs0tPkX6KnXOl
1v/Jzc32nTbDeiMJsdRyAVrVmCYojI4ULob2grr1qO02OF4gNOw1Dghh+33vOjXb
aY+eEb895U0vil6gS7s8/QYb8smNBw1a0/PLNaSwx8+yA0/nhu95P1/yyaSfDQdP
A9K+NEKDWxSSfa+/0z26Yf0vTjLrPElEcv4QeDGR/5vS8xAl8ZVugaWq9d0oXeWg
q0EcA3tw0Srk9oC0z2c+fhglJvkTM2vgeKSUOQNe5rpbDl7AQJUvhxfxZN4k9sEO
19r2Rg/23DavnpkNr8Geo/QAyO1fiL1wMU8qSyzdxAQ4hLXDxJrtwl1wbV8HYkOk
dkCcm7FRk0daDTrFq892xEaSe1oSqPoDe8dQD/OoaRQs1AVmhRdH4PBAl4nabvjK
34gKtL+A8SxcwjHbcFgGyqMFvloNIxH2TNaT14HzCnfad9OX3RC0FDxSLgGcrrIb
85VtcwXHj1Rf2JpUwOfOS9e2qKDsjdq4Hj42GOmrUDYWur4Ik2ZFu8o2h9G1sipf
lijrGwtJT7R7D9qsNmRw+CizVYcGSoXXngfD0YLSfRomvqvtl9VnSNFXYWfVfvu1
71CHDRMC+RNQeBV3Qbg8KzBOvCnFVmdHX6/p8DeJxLF+lshg+u1xMRVvjguUPh0p
3csq9IO19AUTQJxDRWZxqtWlA9ygFJ1SU+Fcz4jqjKzu+3gBg4lAFjfKTCzmJ7W+
eTz1XJatyJ50LkKXFQ+8kUwCLg92tVwg+5p9TC3p7WrWTfbqePirj4q+ARetkGEw
5KxjcA3XANG7HysP1rf3RdKgWBgs1zz2x+HqN6dEFxUM+IqpWaqR/FP9Nt110/dj
6yV/wAqdG8qj9gPhADbMc+A9DxiC9dATUygaHPOG8xC9ap6UQHvvEfVllYux0jB4
YHvuYODE/dZsDqmUHfG2992zWyFjuMweynoV7J1BDMNx3Cg+hMpoJd8B+Nb2Fs6o
XuRE6JBuqq0iiZvZD1Utt/GVhD7yRVtEvjNg5gHLp2k70fKUbuVFebs97itA0FV5
PRRk2cVnu3gUTZrTe4b5YBCk9evx0N6o2pavq9YHG7Xm8LfDHvnd4l1sYs0LS3DP
i6H0FbefCYPazWEIpeh+9eL+XJx4MvAABveLptsPiCyBy4XHngIJBWqrx8vYgbEo
eZdJ5nI4qJdJ0IRWVq+Kn/6bHINSxQhpO/wCoF0qlQcxXAGNp4NxHj7LurtvODZc
jr+7r4Q1xLbt2csVnuEyFUej2GP7ysTLwvuNn6b53fPPxJ3FwH6dM6bbB/Jw9c8e
KbFn1HjQm5+2IKFdEhMiZBDFXt6bVmyydW/Gi1GzpAXFJpZeEBtJRfc3kEiHSxvX
axwHj0KZ1U467Rg2TgofjbRRyz4mhlVuN/tOcw/XKxThO70lQC/6meYiJdfJpnUU
U6mIuW+cKe+cK7ZVcAJ8P/YL6dfb2IPkODbfy5YIGIvtbDwgXQDQqODwIZxIaig9
JdNRrx/CMXpHv8W6U4Hv4oDYjQwi+hazv1NcmQTepnu+O+Jke7ehzewLwAUYceXx
qAtOLWSA3YSFa8JtO9A4JDUUX5YJ4ZHs/A4ji3PLo7AbK0olnnquH2yLaIs/UEg7
II9qOFrmFxFRo+ovda2So6Q18OP+wDrwMmH/TTlz2aLVgtF2TDIriH/6Sz4DVuby
hh86jNaXl5yrutr3FTFBHC8o9thDzqGgd9RxmY1kxDPom+ntwRE9vTI9KgzJDuUg
IhfFdWqwYdW6Ckgy8uI9ru4JyAwBoAnGreFospsQQin0Re2woMfdzm9/rFTsJtw+
rH+Toh5Gj68hUeJEH4dsQouxSQJhUYD0akXqcwD9C8Y4RE9r1jZHYCgboxvpqHhE
8FiqXSqoPadm+HS3Fzcq2/XyUy7D3GbcZJTCJ5jbD4x4sEd6X1sY02XJaecwABb7
Dwq7oX4xg+SIiV8syKpEzdOdNBP3uSz3iMNFKLPfCDr9yeeTU9IVSN3qX/sroEXN
PdvPpyiLE5SycMd9FBfnIyv6/4HYMLAAHgm5vt5zVWV8mGXYcoIA+sbppL9O53gI
UKLYRJgRWMuw9W0Qr+/fLCdna8qZydZHfPS5TtUMBstIFFkbblmcVRQBhsbP3A0x
ptol1H5TfQJ3Y+odSAdXCJ1Kuow8TLEXmyjgkrBHU81Wj53BHgUTEQK7lohJhaXC
vZbwx1eBTdSmKL+dZ2IgsTnc+upw6xwBrA+j5MMBxm7H3CBSHk2ZNK1qw7dCbhtR
yJC+zcvFQQVHgX5bpm79t6/RCPFj3fYGKEfXHwUSmiogLXx3mi0TlFoJVpHb88P+
N/NwC9u1nlve45mS1FzubWYMRmWg+CHCXFVNh1iyhL+VWJ7ymzl+xBIoFuMDkWLc
bFDDX1jfsqGXmJrs7ehDitUjRE81EhVEGtDNxYS2H9tnBWMPwPOALj9z36PTcNgN
4YpUrSCjxu1glmNghiBp8HjrM2TV2ZCkAcjl4PoBl/28s3tJw0yu9Llfqwzv/mWq
sHdFybfHvvRSOjluW7vMoC4Q75Zc3dM8SACNR1InVK1BQ9Mz8pN3R6YPkRZ40jSZ
mQ49ZdPZ5ltSSTdsjGC49hjGMX1ROT9LSjoy41bP8KRC1IKAx1rifmr6bxomQdEF
gChFWnbwzVGMpRo51dYZUCCqAhB0GNBAypuKfbii8n7RYBbgz2YkNwSokVNxaC33
RaECr1b/oopDTtrO21nccnXaLx1ZzPIs0dXBa/PPKK6FLZ+XSIeL4uFvzyBbrbIk
FsR/iGptPJrvxvk4EXvSHBFNbPidlOa8VybiKlpwkkJAzbhntapuEO65VVxjZc6V
jXETGuKVoolQMUDulKMaJP7AcLejTYgEurOG8wSJq+Ypg3OFXlg5g5hbujXNkjJL
KAWZx/pLv4kJ6rtmiHRlpa8kY+mjYlgHC2K/hRlefAxDmeyYy3IjvWhQCi7CI8tM
D1BR815g6BYEyk1I05zMhDSHvBjJa/6SBlJZyS1T7KBDvUtmcli9DivQWu0D7cfk
Q5n1lGT6/B5xKCA7fMdo73wvLD6NHv4rCjR9hnJEkEAP/Npb/Xf2SXdKkVz4/EVG
RCnROzoa7mX0WJktSccMRRuwYF+OOsb8TAigCaiuwWtzTvuO+71OxmUDlxbaq3bi
Wvg0UQ/hAI0MZMvCV98qRPVeZD/T2s3+ExwC6kdhTkDSK9yGJdu89gwtVPmjfZ6g
gKNhPbokFW44teiWj5Bcv8PeNE5QmgZxT555H4ntm05KS7a05jS5Pw3CCmUE9t+0
DdVdxzPrDAsbbSHQiET+xmdBMufsxKTmBZhZYSFXPA9yX7BLbL6HewkHh/qfL+m6
3ZuME5atmKXbiPrB5s55T2qMYRhoSjGJYL9fitHz39i0mzNdxCu9tngTqNqMxSbe
lIvKtMB4MyNdsKU9whxymjE+P+sxoPEPQ60dPdhvWwLw03oRTalAI7IOARo3sZgr
/8Q2vEptyPZf4hvjDZMkN2VwfKvTxv93y0mkrtBA+2k0cSgjP8mZJ7vZ1ILxF1Hr
e9tap1xuZc9ix4syYCAAMpIq4MvK2FSXtIdPtmFFrIUmTXMwb3O18lU2WaoA6DRY
pfNMqgR20SjSw90prY+veZ/OFuuyqr65jaRq6EiS4iy5gXlJaPQnjp048x9+EbVg
egTcnYzzTYz114+Fet910KgZD8Fc2VPcLWOCs0hqCjATsjbTUi3BvY0BXWEYsBK9
2mVNyYLx6Aapenut7M2xIjAaFHyeJmY0atYRMps/VL0mMDfbL5fsWWvwMNyzygYN
rcRfemLlquLUFogT0DY/ktL8QCvuIbJsAeRn9nUEhiBSSp4xSeypSSHf7JKqmtFc
SpMzzNjwshqSWTqlSjEfO0tNacaByDa5Y9rF5kvZIZsuAn3U5IyA4IqtqOmisw9T
vY5RwB+HgJuGoZnr9ZBFm6DJ5EPrmTZHzukJAKzEiKDQsVTGQENmDzaDeHjxavhI
nZSWwMPlJrBtFlirA9VdgdguLgVxgvAdoKEIiZspmY18DR6sq/Bs8urWsQ89sQzE
izkbwgzZ1dzq93o5kJXQWgEmtiTyDnoinlYbj654CwNYwul48HrEDUnOlPJbTPaX
cr6tgKb8I6HuT8NHpVQZkzZ3Iy5EaastWVjeXyI5Rqf2+Pf0XD9Pth1ohzI36a4l
NrXnxO0A4ebOO3Cc7Sp5rboDMgaXc/2VuqOXCocxXQKG6SlvziTGjL/KO3nr3K/t
L1rBb6cRSYzGdvfZQvLYWSjEqHbG3BHHz2EGCeNosn8I5LI8JFyJrdgTJEQSxFL1
Fw2DGqzom8fJJInvGO8EnbR8iDvuX5V/KyvT6juEp2PtgDLzF3q1a7fGH6lUVYRn
XFT3AQK0G79aGHX16r/sbqIVJ8sRFDqjX7SX76eViRHoMvCzATokmVrihkJjNsw4
gAKLBvw3gp3NFOzyC0Py7OAPs0GpwQEi6ft8jTHbM5jeShI58gUmasMp7Ejfxgn/
px/EqNnusoIe2Bj1555t+8KCofv4znlW92BjUu+P67KEuxjvPT5L6HWqkrrArpj6
00mNIWEqQ57uaQEK30OwMqDjLEJe68ucfSArsvpC455Y2sr+NzC81Qf7e6yDo8KO
fkjvtjmXqAeSKK1wcbFpd60EoKnsDgFunmj8sqqUShMZDpXLZfPUn14jxFisADUN
+39q2JiJdLlwv46eX/zlVzaStuUKgGDTYdOz+Q6g5EWlvQQ+fQWrg8JoFTEj7iFg
MN+y1aLMZBkXJYqFvgaq74s62Tz5iNOjhplM24oCm0l1w0bGU42bftE2mj31vv3d
WAj8BGxu9byMdwcwI7jnuuwS2yoqlgMgIl2NthPKT/raVRWOmd4QSGpZvDRWPkD4
aAW5MjtyvKwHWDvIPlJP03bAf7Sm3jFd61/NT9sw3SegabfmwfZj2vW1Bp/7zRP3
eE1DubYa0hnRcBsr7jfUEeEJtQw+MCmSLXCSsL1OOuhOdvf3JtzM4hwmed1oDcRq
DlqdDZKD7tqDa5UxL/kU8iVl4OTa/RHt/t3kFyziLTuwZgyqqkl4ddGvtzM+9wqa
8GYq2TLZN/AJWU/tz75eVlCe4ofGCEcFsaPuSG+vFQLjASKg6+ucokcRiKEm/1tl
xO4JWLyhFlSD6dOzGFtu+H+c5nxgmTySEu+anj8NbMeEfvaa7G0LHSlIeWQPMB1A
B0C9bMIjW33taTIfV8Uy1O6rLJcJcBkyDKq2t7QLMCWaV4U5L3eJN0F2MGlqn1Um
yBs83m02a2DLBbZv4XLyZXG4t/m9fvlcjcBHvH3LHvbngLn1E/jy9ZU8EjBi2hZi
NUkpAqLT0eyars4X3uFEIzdUI60GHOjE3kFJH7dt9QwXKMrLZJC6wdPyyjGHKtOg
gE5liHwL80gS4+PrwFoQIOTf4BGX3f11o4KJ8Q87XDu6D8/lINXWWqNyWPq6wgWi
gTW6DJ/6YfqJCa2Ww6rBdaFtfcOOKjAU3NfIBQIMhdx1pNaWxF6jIe8fmqVCafbi
JmCKKIzoNFACzyG6UCB83SnTBu/R4wFhovkLobG/RmLmSJeA9g9v6YZhtnOeLnM+
QxWEYIHrU5XcjLHmgoV3uPR3eODE8NHDvpkocCq4ELzdGqlEf+YhAkGg2PMwW4vm
SwO/QWYzzH90pOeud4UD3erSHAYxgNRht4usSt2f5MdNqCQAmcKAehwGrpZCDCnE
bHYIJoZGPN5H+MdwXaGAs7DUa/Mh/kk1fsqY7stzotFqrmoETIV9lXdyVu0b0Hum
nWOxwKNydYchgEFKi6+cX7AvMRbAc3CROoO0DkM+EJQZ9dZqgfm7UPtnUiss5NH8
/i9ioAH82r1TJNNJB8XDV7IQA+d/ReX9FQgXj8DSQgm9Y7YW0vB1Pjc1sqqTRtSo
RchaTxFnlF64gAwLdghOxt0vKXjiDl4UIt03sMj0MM9by3+ZX+Yc6f/x1gT0VPzo
r/Yp7223T0zsoFFGhBGHNqZovnpDTSEAXDpyuTArwTS/JRWpzAPAGxnFJ59W1I0+
1U1hmQ9jdWMoMwlvk7o7drkYtY0bL62t/J1l5MH7E6HIencH/WPrllZOhNzyEG2l
ECDKkoM/TvW9IwaK+FCQ9Hm+UAnl+jkU89+F+XZbhR4ilwPfjlNF8+oojop3b3ok
Nk8yjiaCME71OhCzulbZM8VS7xmcRJguKci/c6vzvFeJuQAbIpcv7x1LFlG3kpNf
MJf0ojCYkRtz4LVDslWtt7ET/BKRda2ur8EPo0p2DHMbKLAJt6YNwZSZo3p4IvQ4
mAR3uNZArVnHwlHGKqU3l+kycov7vctH4oOnDcG0gIAxwlA8E0EQfJpsQcwLJnVR
266AkZx9t6rqOCUlWKNVhFAe7c+3g26Xegw2LxOUQ4k5gEyChIVD0RcKbp9yDmac
p1QdlDmdITwHsNik5Aa7RG8cCAm04E5lywpF+RAEKgCgxoDj4rLPZ2cWXMjPwCFz
PAbpQ00aYyI02TT49Ovfcgk6fQk40pcAhv30rn6OGVN0L8pq/+UB73zzyuJ5HxBu
b+X2am3uaj6tSBRnxcPsakTw4UobtupsMKzEwP7Sm/SNE7dJ8Iq696k+Ya4T+gZv
5AR+gNXeqaGTyP7m2vohjoEbnEON65/Oi4tfVAHOCXLRWMW2Nsy/ji5yM9bnFaAg
rX6j82Dqz/9Qtp+ObZBR2t+p93CwDV2ljgn8YP/u+6PalnTL76B2gKefRcyG7mr0
9XbXTpdniA6ztEFjTjUkccQxlCURIyCFOjI9OK4iT7IcXoTqTlTFD8+oTHnuF024
VJ3nwQ/j+ycH0f/IayzrrVGby4y1WjcbeuiEWNKNl5SDTdulGtnoukVbO+JPYQs9
fAPCcWmQwpmiZjEYApujOT6sLQWzsXz54vti4re4QZ1w8bNTF8kzkVsQL65GpWzI
VY8PluHjX10ubrPnaqVpemMTH9EZDk33oGz7nOQKlSPMQVgIVuG+vc1ZqMbHLY+L
MiFXFEOqcdHj9AgXCr3oHPvgnI7m0ALihG37xAR8KtSeIqhko9vfxWS4LWzzqIkZ
aw7kRZAiOtxsrPsDokL6DSQjjzItrX/D2EyX4pA45FzNXSDwZ566Ur6ZDAQNvsQK
BexFzz3Yar+wZ3SVFC2JjNEIpFjbOqSgCi4Y1yJQoERWjlg1iXqD/rXlah8MrLj4
skm6ZAFPGiU8V6CfpRUcr9/LjOnvdm14vP1YkVk7zPY2mXm5jxageoeKWQgenX24
507ekricvYK8YM+VJpQj8Hz+bDmAht2wnWWqkgpxWacUifimTe//QBlYA8k93yZS
Hu2gSJjfcLjqS0aHaNh5LscggY0xZENsJgN0Mm09R8bg/xoG+S/oSAgE+HPP6vqA
BmHR3spSVwWZEsRLc3LUJknfCH54VaAibd1f8hlmeewui0ejOrE9URw1YVv/9NFV
8cPBW+hbMIU+0Ii56q/PLGUDZ5CSbIMtSMklIqIxHm+GHLUoePFKkgDvP67jnVc/
LRS4bNIxFODWYwNF/Veg/EM1wmyyfXarUq8pfExWm75aPOGTe9hNdN2PkhxdVL1a
cu0ErtjlftmdodvolanJYhXwWW1GPo2tU+G0G98IEecnuZEnebQ/2rlvu6VZIoCq
T7XtAVntkD0JWKtQvP9yi3/4MF1UgLUaYTY0szef5qo7rKT2zgq5WLWASniDvGec
OIssdczXSfAYfyNVihKSHLXOCB0rsqEgIEIdNUEDHmnXM83FpU/b4Sv2GRNGaLN6
7zj8WMvvh/VRA5YvicQFVGB9/CzMFaFDOlHq6/m600nhRovcJbPTJyIQ9UKNjsgD
EwEKAxG5XQFENc4/OVO2V34dFo6tH3Vv9Lm4ELOvdNRtjW1ZFxgGP5wdxLkyQie9
DdJ//CJYaAjHW3Cy9H2oTqgoxSL4/2ESHsGAXHDBaAfHOwmoumZb0gf8z/n5g2c0
pfC08wVp1zNO/TQXRWWie5v1I4qNKikLXN44lEESkluRo93zB9GQl7FTLU/dwcj+
5uIiMg1bkIeGbvCy5y9D9EJIzmnp2v0Vng538N0T8KfanpJaV0VtnATKOmgdSjoX
1Nc0O4IgZViqxjpTlainyfsyjUCSL93MVySYfbH75z+XnWjMksCziwP8vxKCgxoC
p/VhA0YvpLLDctW/sTrMFLyy3IByfZJjPdkHnBfv8oL+NFX/YULo/2kWqZ35fCj3
18yaEWAySXfLRlkNtggRLaDGXPYzafxcxG2KLOYxL3uq6oF7hLaPyKtyWzESzbTe
0dF1OIOQj5bH50PixslaD8KyfH6wFZpjru8hQG9CP+VM+tf3EKYJBx57DCVO8PQ8
S/QWE4okVMY7b5gQZO5x0FpSK7TpYrNvhjHGnJujoDMNmFe/69X/BIjrV8nBFkvN
vlEu9bSgfwVR0zZf8P1gNDQH1fK8d1wBTHXQooHRg1Rgu87OObzGAWkPilGjWIW3
pX7bc6tyQiD1QlE6C35ees9DQ6TPN3apE2pc4K1QBdaATPff+9E0jZ/PFqmheQVt
dYy8RcmY/+S/r7moH+IFyAuTiWtf5NF/smCA73wPJeVusxsz+Gf2IU2jWLT26weo
gb4QoGzcyAtxa7s3B3nrC6uPy3/Qb7Bq07SNmh3OIz1uNeq/LzyJnM1ASDLgNOL1
SFZ5Hi84fBid63kcvkKw5SgyPcy7VKdEMujQ1bpIfYQ/w/vrcRaTh2KZXA4kAm2k
SJLOy5U9DHw+0vC4EPsXyDt40sFqwrxbuzhjfyVy69PlnDAEdKzW1XSxzXglwQIv
+CUpNK70puG/O/Jv9qKs1h2kPOATViT2Kpf+0O+xHi1MU1QHJTx4ClvFu0R8EGA/
prpAbiJvdpkmo51Bqq6QK4YNuAyATjikf022p7kI/B6sSsEWDXHu1lA9PiRvCem6
am2DjqORIpa+/ODCn0uv25Xxt9qBLPTt5IEiPgyqD47tWccfkA38zcfiXDDDg5V3
JhGxuXVgMKg2yPQwp1lSuWNC+nS3a4z8t09CTdIyQWe1APwlh6uCam4ZCLCSCN4+
MWaH64NPiZKns9ySMHHijJdIihD1rtK3g8/Kk1Xev2ssD6+GNbyJQFkt+2MrZyfp
GTrM6sSNoDHxwV/fi2PSyE824savbZGmpdSMH+f1WvUpcyokk7pFMGR97VuKhENo
nl115am/zwaosYpXocLcdev19OT2POaJHB4KUt1Gbg/n+fz+64VVOhQ6hOGtTpCW
AoELWRiE1FrDLnmnPQPTaBy1dQPIgn3LVd1mpQ0kVdCFCqsQwNu+hu1hwoHO2vdS
dsegQGMLi3mrt3X+rjIxArFmb6Uc8DQEPiJgDogA4MU+8cawJFaDohgSQs0lz8aW
RC7c/nLLBYqBp0APDlPh02Oz8kY1ZTlX84nyAOQpdOlixNTO+wxGSDOIerIZKpcv
KUXznqAKhLy5+l9q+5JicONbCgs2hTe9RNAaWc48ULWAJYeR5rE2tNni/hbOWnH6
floS7q2nhUof2D5g8zXmS0JUr565d5foVPSL7auhuFAtur9LykRZvPf3T6cTGus5
K+RT8HSh5ZFVWWaqEksm1FSiICAT9eBNo6uF1nKmmAHrRtDCqSVTL/S/tL1BB/1p
DqQk8AajNTIMezB7t7HqnGpe/SNU1Fw+D9x3E+sEuS6gXeS99Tum6KoxngtGJeWJ
IyrkyIU7lEqAzkjT/1C3sfWpIT/WTKKqBoV/S3maFBU84SH/ES76bQ4FrrTgiXnK
5PRXcocjHSOE2ONyALLPA8CbLeSJDPGjpplAlx1UWbyPO/9dsAY8uapdIiX8BlvX
FodFtlpzrynEpOJjTEWa+HCJip5etBPC8a91OmfUJxzgUHzJj7Vu2FxJiFcOLxKj
CZ3mzzbGowJUMd+rm4BwKJPQGFIam2+clbON4EYUjjYWU541Xx69mibTpSIgHezi
/w9O4NyhK3HgdEQnBQgYgBUnjD1aku/zEIfVD61nju1VDJ+7pHlmw4aOmQfA3xRs
ZFmm45mkb0/pZSA9T/RELTDAkq7NwPW6npiEQO9KvX+CQsxSnRZxv0T5yaMNwd4a
NxO2Iyawl946x0FGSmnYSiJn8Kz0W13T/satanlY6oQwWzh+pKTnj9ThFUD789Hm
hxyxfatfGcCrlOhUffM2JQg4b5S3RDvZlsKXC8bgh4JmAAbel8wFK2x27gOfd+zy
ajQJOXyVz5MIrEacfXuDaSova2upsEcCHBYC1lh+on88bb2BDvV6tgoy7Ot6clqP
KjBuRj0r+ovYgW7gWJsPnFlSeD0ZUSOI5zsIjoRhWur0C8lS23mxjcPX6Vp42swm
QnnOBXQacu9mVBnri8EBCwjwq5Dajdi3gjMnXYzO9ma+fnckyFbqS9T+BgEGyAiU
NeXkJ3ZVIeHm82d5Dap2xssFkCphmlR0sDbdVV1t8sNY2EoJxWt3YHNBVY69YEHs
1kc76Us5rwzLvu+1rrr0+eSg3KMz+6xgdaCvX4kB4uBpQggAdVFSVtvpEyMZ+xhv
gKIe1+sdDZ0sISFnwVCEHN1723eGzTHL98k8UZEm8ZYHq8JOC0JwVPhg8QUGeADJ
MPD9zhfIqFVQnJ30LxyAEg6IhENpLh2sMWKbONVowBuefC1KpgeQ8uYV5UV9nzsQ
/p9qnu99bh9Sti9h8Y/RzN5KNZ8BMAdUjl1Qs/5txjPXqC9MictiyyTdgXTo+ThT
/JAtd+jTcW6nZRW8NKfqQxWE9aAD03KHssPNu+TUZfGDBWG9XmcXTq+jEhIuFw0q
xxK5z3KPvTtGr+KuO8XP7COKTRZiyM9UO7ztUP2NJho2aHb5VPyLtcsgG4Gd0n5h
J0kNo5gxijl6W3du2sUYHbhb7Q723W6Zyx9VxNE+0BSfSe1dR4S8sgCXEUq/xflS
BZLt3VBleTOFz3QSHS+FKi0n0XPEq3OqWne5/n3Ivh2VAiKpl4QPibnttbm6cJFX
d+ZAPfhyfSLc2XJtQeHpG3Ipceg3hbeJl4AFW3Ai5rz3mqXugy3hrMJxr01MVFLp
wZ+sbDpJH3aGpJHBKLnMDtE3Y5NreS2kAQQVGrmQVWoCzl4GwGAjkXjsVt5oRepp
sVT4JDrMId9LaJYfkOBu6agSc9DJct1jokX2yPqcuCTnhT5sPBRWzAHnCBaV8qEK
K+ndCiS2CPLfuE2MfTl5QoggxhZi5zqEnl6HB/KLEJR8uhDHYCqxaI5n95uYdy4m
1h8le52Ie/nYhwQ4CWl0YufbZbBb8xO0iIjfJ5arFq64+m03qDUyZL0hYqYZRRZQ
/5S5vD1kTN8UfJ2Bxr6WBTQ0WsOuSgWIWn2EIHjWH4Z3IkAiuv+WAxBMzJLufMQM
aQfp441KLq3VL2Hr02i5MhH8MRMqR0Dd9kF0m+OuTkTHbOCca3PTbmJOrjHPFMRu
YpBbjTA0SreKXSpx3TeJVwbfn9g2L8te+05TXTHwSWzENZ+MAzVt8yfYmgMRuSHh
CGPapoXDptiUJZuhzOhKwfVsEPJkTWVb5THTLWrl9Q2J+FCTWOWlpVeW3B7sBJgW
j01C1ASluVWohqqnXmR2TfDLRDvwTacijQB3Lot59JLr5LkOmwwtwRUtUEr42uys
5p8JZ4dRTvagzJGoPOBJJS7ESArZBRdfzlxAytfmm1dCVtVdgjwbVUGbffZ3pWRF
RNwXeIdSgqck6NQYLGsfJLVNjL1KS6X9v/+tJCQpxdNcO/uUAf7wcfsr3maDg6PW
xYDELjg+gB6rQX/VnfeLwOl1pdHCTTuWHcIxLrB7qWlOKwYETtDbX0nc+Pz418bR
WvvgLuQYKd34NRSwM7BvU5Yf5O3UFI4onsFY3fU2V8vfjz8yOqwBguxnrmUvYBYU
Czjz/W8oT3vs2wfByuGcfFMsbcxFRtXDx25PAuYFGAK8MTBhupsX0HTmeNZQSON/
aQ7P1K5XNza7zMMUYLa2evFdTwCTYgeTDMjTXIQpqTFs/DaikeAtZtSJ66tcvabW
Rb3DhiIfK7GaZ+2NfZ1vRhvdX5yKKvQwO3EZ7Iz/wREDHhhDqVw6Zdd69H4/Q9TX
brMdNXSKkBE3bH1Gj9HV4S1jKq8qmYRxq5PmwR0jgyBbdONZct490Z3NbN17CcFS
3M0bJOB6uFeT/YWmDVL2vEL5lwqE6Xlj6OQIwKTVp5WZYxIN03OiXy2hIotGK8j5
dNqsZNa1+DCySq703L+wML9yk8PxMKoFv/c1P+w9XwT3HDNe8CAp0B/3LwbXKvEt
qmxeoreyJBJQssRJD0MzrnOQy9o5wxLdaMkcdWX9/OMl3k23ZtJc3v2mYCJI+MwH
7Xgz8/JXSv7QZ99st1aRVi1bx78AkzcJZ8arTyqLgb7NWCzr+ANMd8UMWSLix7h1
ZFCtuCsCYkWtkGNrZxidMC2ixwDUcvJ6GH6IHuEbg8enHTcMWtjyHE9N0+7/C9qo
W80Qkzp+CfU31c+22lsdvURPddpbD/BRj6y/3bvo7fKzgtMb6RM5ete7lW8QaDTR
lVbbViLck6QvBWQnjWFi3Y3EIDjWU5oVCOHbgKR4RPF1ho5AvRWwuXlxZ6ZJugD1
6gTp6E+7JmTXkjEUpGacrZIAKvjxep4iQeFGJCyWonDM7mOLWCwAqsp/1BDvhHfy
0ptgS/A6rF/aqftwikyPOPf/lXYyrMduAMKurNN8fkS3B1T48DscyALV7SvW3UVs
hWcFBpa2V92KQfNExEj4uTlmYC4K/NP8ZrOHMP5azX8oL7NVl9HLu3TNPKGHiNr4
dK/KBR7EqJyFaW5k+oeiU0eq3SCKCiiMW3xnAWoriElokAc2iyNJUtlXnNFL6ynh
gFuMYo5MHUJ7UJwiKkcOeAv9jOSpKDXiiFNJINbGTtYVhjUvC/daEtcOBrnfoQFv
2FEEYmKLWUyYncDPBs7Gg47yXIRMqpl3bMAxwQSBlBexJFAVDEGR+q+oT4f77OUX
L7F59mK3bXu2yaioy7yH8/yHme0+bHoSLjjIVVsxZVUrptL3ZfGIgKuRhzASAzRJ
U5nu0SVchHAc00Cr8Xz6bNwiYBLZ6RforGzpnBhQ/VnWVd2bzGG1AnRr16OIAZxV
b7X/qXxZqC5KV0dOIj+DwEBpH5rbmt3h0b6mVNypUdxVFJFMFyw7IC2g8Wo6I+Fd
1KTGxLakWMktMARVwofU4xCBp8qRJz1T78ZCJSPSs7OW7wiMQSIyKcz9OmNBkDEn
9yVG+JI8oxK0WgN/LqoEjNWFcmQewSlijjyw9qWcuz9Szu1g8w2gr2Qy4Km2nfxF
2rVCmizduy0jf62pJOumamJyr9qwFMwllcM0kUyUMtvudy+QyW/ZYD6lgG+8ERQV
iHzebOlQjkCIcUo5ReXF0CzKBY1ZudqmomBHgDhWUGPmeP/7NZ68g77y7kZj1DzR
ezE0zWljWF21/omRIxHGvX7gE+4Ymi0aVpruaj4jbd4SxbPjSGeEc4JvttHYMmE3
yXCW+4zxUSM/8TryvN01Ny76bOXSP0KmXnlm2Ts5Cv8OWTW1lIEEheyA9QR4ugVL
dfG+XuPBo/b6UtVYeWpZyo2yD/zncf/xqvPoWuzihg4N0NoTH2z/nqg7V5y/PYkk
7TEyDcKc97LAHd1JBBha6n9mxvfZmHb+nHnrti80FnrIXedDFymi0XOczU+9px0F
Q5Gh2L7JQZ3PISHkaVosKMpdmNI7eA6cxU+fBv/+V/TEB67HESs5wwnY4qZqmTS5
zgzovBYXSjb+wgXE5IueNqFm36bbDkRzq+tm6RGn6579ZIOn8MfYJQJk1I5b5jn/
YBIcczCXGLYNdeE7dVx+mDbrCoAXLOEFaFnXbUxU7HBUos5OiPPq45RjpUy/+ixZ
wQzhCwXQTNo/vTOkEYcf1kUllZ0WO/Ej2JAU1ql382dc+05GHhBmQcdso5XuUfof
+KYU7mQsgyQOa2SUUxOs6jbxcWBlocE+ESWIysDbOwmmnhpO0VY37SOXcgO+eVnB
NUs7RZXD04ooCHtHQvPESZ4Cgajrb9liUGsDUZf3vct07ngf12mKXt6Z5Wlo3naA
ojDPMnDE6Nkwdcj5pfarHN3J5ggfULX5cB8USK1KB+r2N/ckYjihZd1pxbmBdd4g
nC8+Abtd2FgB+LOvTPkxcZXGATI2rkl+17RYLlkie4w5ve94CK9kLj5F+/hLIDRD
E0sZBlKXC5aNpMtoWthPF0rzsN6799DS6e7rsXOCfIqplZlBKH+HzoOm43B7+tlF
gsVbDaRAdKUtaynzhX0osIXVkVr+/5eI/X4pdl7qsg5HQGV3l6dxbr3Ef/1huktk
lAXUfQUJUrlI0HIr8wYI/eaJfK70gfdusKAaMMQODKAlU/swBmNhR0oJmSiLUEZl
QgY9zcN+J01KPO51lsWDYbqzfaqHVOYORVdze4sQ3L2hzUsokhvuldmPFgVm0Z9P
XTLsuQujWxDERySvIoZxcTVMNXzDrjLZGK6Zn65kI6yi+WYN9oThMXvU4S4tTHc/
Xnfzl2DgGl39RGgcHRq574cschOUExfwj1X0yVk92gw2OrEMAGkfuQgroCm4G8DG
jHiwmMchDU47Df7Kx8ZXHpTiNuhE49PlMjK9J6boIJWm0/v/mwcmUUIgG7MqKYt5
jW0XgY9XbHMVjRvaVERRiMKC1AD7VoMQxDNlB9gN6l6mYaR90joagWvMYcjGlZnf
Cude+kjgWKMhsB+EiQ6VFWGXd9h4SkgKNZJRi4PnFIHi4+y0XHxu5u6CMeKps5To
NaTKJ8MyJDGpnVFWW+QV2geZ+r9i2970f9Q5VWc2KqzRbcFyQoChDkCxm++XemW/
wVx176RArJHU3wpGPqEAzTGhK4J735x+7f/1EorObifxFX6McAmWF3GSOWNRuHJG
TFru16gA5pFAkXfNKDCrS/J6gDlfosT6hH0IhObU2ZVPP1y/bIBUprBcofeoFrUn
VavZBuRYNwoyHDzuHwhiuwyHnyHsCbmufIpimaQbks5YEHcJfY9l4hp2S5+bIAdw
hDhIrhNGsq6xWw3WWUzYR4Pjps3B8eCZ5a8BHKGgokjdX00JmYZnOm7bn22/mui5
erPayg2CbEObbP0ihTdMkJfxOYvCNy07SnpK85GYLJhFs4zYfvpsIh+7VMDnLALf
SSF916wLRgChGgPpI5LwVpGBdYVyTYVYdLTYlEWVXqQpvzS62C7fn8X0hBOaM2gX
jWx0XN442xHFe3Kciq/daLeY7v7bOsUrvFBIKdfJ07kBOIPWXVjXXKez1UmmnYGP
p5KSRED+wgAizkXUU56xVQLPKOyARCrH42Y90SeDTz+v/yQGbm98IAPBX/zw4jvX
zTaQ+bT2br/X3jYnXev3KTypXCveieEm4on3/zeqWmnEph2s+hHHEc2TZEcj/dLU
q2mp8vNH25QhjGdb6hjOn+6UWqIVCy8CwsEfNuXihe+En9wnVMQMsyIF54DsDSGS
4o2LLuLbmzC0eb2qoDSblrIp7Xi4HcNn6RDlKpL1WfOfnXhURRcic8mFUJcoRfCg
pWac59NYXMFsI3jglXG2HVBpWb4l6Mu9oZ7rhtMIuHh+UyhmDNX6XIIn+XYa5J8F
ENKU3gGUFU9eg4tfN8+CB7/AxWeiC3k6mqQDufala+Z7dvgNN2oUiiM36VEdR0sb
oHXSvUE1BwymNsXTtTewng9+GLV/exEks57cGn8jJ6nJpqNthar2lPj9UHrQgZu5
tK0LwMNTzIZNKFplnwx6G4tGiVauCNr6V5MXNyYAShkZIRha5wXPZGZrHfciuXij
vAxRfMBgOJSXFSgLNJN1CaxCzqicjtnyiX+WuRARQmLPdznIwSQKE/gfW1xhvAbH
E3bvmtBVpo5qzx40NlDfd1CYhLzHbM8CJ3JCO6GfRQq2+FZ5c5nl2DI/vIid4sgJ
ltssnpjt7aaGF7fZYvMX2S+HmW1kZvGqYDTiW8/NVns5ksoYtanBf11UBef8M42j
Lkg1j47UcAGkK2H2Cx7i6EJP5TRpiIVTihoEZtO2Heh1INYbc8yNNnJ6nIf8jBIS
zB+kQbzdTn5VKvFbndhhmqqaBIFz9Qe3dcdO70NE7hhczVlT6bie/X7q5QrX6vbJ
onMWPC4w5H/mEi6I9CiLjeUpc0d33Ld4WuZKFonXfjNZoFxt7FuFgEgQ93bTiLh3
EATdH5KuVq7wUxouBiyymS+jR7MtAMgSzRwFonxVHDNySDFnMI5RhtAby0HrlLNO
3xycsb9PMh8fgc610PdWexcUGJHFPX90DTRuY42DkQW5H7528l27G6bjJwc7QEkG
PZ3xZ5yYo9V2TaLRKi113Dp9MnWj00VZwBi3mo58+FgaukAxIVlaNzQSyZwyqsh9
LCH0rRjsaBV0oGALmX0P7tg8zOmPtZJClUT4bUTjL2ldeUUs+c7L2bwnOe19hT7P
NyCIw+7bLqwoTl5B/oEmWIsTnzLghFGHMmKpft4JgWtvG/oXtZcJtE7s5zFkes8j
a49wZjmGSmJ+dH2DIeeJNJYT9ygRDEbodz9UjtasMptYeV7ej/nCqUWVyguOkM8l
weSRklU0KV9Eat+7agrHGa7LzAh+DhClUlX4cEnxJm/kMZS4ocImgafE81h9YjHU
VxBo1pIgslfZ2dc3Oer7HP3g4wfK0w7JGXR/dsLcwakX83IejGLGyUDZ55i4YRUb
Kzs7oh5A6y1zWVrnYP4vQP+7Vs/m11yi0voBo2Fk+qttIlNyZCq92KM+maGu5tHl
lOFYTveGiLq2mZTnUadnZq6IDdrTnWOPmu1/29BBKdmSPqm2HZPA4eW3KVfmnKnt
G3/4WExC8YS/pM6DljHB+EwD7UNr8EsbGEKO2IWPUxN5D3VHl5j5RS+PHtEuRap/
ZcriH2JXbI9sRLweMwhUK5TsdOvVeovfH4amiAfxW0l75zZzdzi2ltq4KO2jrpC1
GNXngQnV17YdnUOevPun2kZgiVb84zLUDy9ku/h9P5nKu8hn2s1SDehe6j2f46/N
vr5y8oQ9u8HueBRTMrpNbcuhcUDR25O8MAgEL4QiXIK9Qjr6nw6lQJ9Xf0AvS1bw
ThMGZij+pPkwbHHrLAZ7YqA5drjgU09EtQhBHF/EXglSJ3W+UuAG+CTApPsOcZvW
RA0dnbQsbz1gQ/j8+1Z9pzvgReXPPDMa/KkXXtdXmNQfBtdNfDOTHuKtMeDzfYcC
r4Lz816IrZMqisCs1CzhPDCALGGlg0lXhe62laslMlPD1tCZZSq0QGy2f4YzuvNX
WGt+mtmksVgfIDzI5u80IeyOzEFmC1lBHDm3e0GS7rjbD0Sj4iekJ8rJTsYZ0zm4
oQFbLLcpN41cIVUN9Ahkh3MPAPEKByRHLvNMCEOhHllfJ3UjFofJ78IkrzoBLN4n
iowYH8jQCiiy3ThGH5qcogJ/1Z2VlwRc66TOAp6mGqmVFOJkUksmGpDxGf2JOJjf
9yQWCBkMpmz0G7oagyjxLVThTtrq36btQesCOtr70zss+IF2AXddGxeGNFXiPXyG
jemVZIJnHy/MsgVzHB6uynMapLoPKu5hfuYX/EZp7F3TyRvj4P8aVhdEawmXTpPK
i/Gzn5hp7tyau45SdOmvU6Y9AlIhq7bI2DxAZVsHvj+oWbevja4k7JMYmlHrJNuH
K2qR7enuswVKAI111idCibPCfgbq6qwHDlF2HRgAmK4Tw10FB5IzTeXcsnd8rQFj
Afdw6u4/EXW1skM6FsF154k6s9EF06GzYoxzavwDCCuzCQ+2EsByL3J7qZgN4XKK
iS0/HDBRBJEsZZoFIhNMGCIVQKstIdxj3vjinfZvdwVzQ/ThLlMoORlSy8XM59lL
eKxyNVo/O9Tuh68L6MgHGEHBDFVWixGrzFcXp/5O6v6rlW8qmMNEYSBx1bx5Mp1x
dPr/Xz/G/PeHby+JRnnKkDnGRgbEcYbyFucMXgoespWmgwCXe/gO9MLNud7K/03a
R/zT1XkOtjmeSBM4fu+AR6DSM8IUm3onlAaB9Xkli2xlWcrT+FXvoS7o0364NL3t
05Qm2FX9mdC6NVr266bLE22wl8S6u6dohp3wilLpJnFdR6S3DYsP8AnFBqg3umFf
Q0pW+Vks4ktXFaTcQ4NKph7fwqup8hplzzAkwyU6iwUNMyKjdSXGlCb3JMytTexU
4rj4tyHGl/Z2cPRS2gWhdMPWq/fbDlxkLA26rxZ7/CmVtmHC1uoAvKBEurh3dP/P
IjkKdgvW0owjAhqhbwFXXLFfK1Bk5SkecKSH905bAVCL9p8CjUfP/mFU2biAAKkS
Rx00lWizBI1hIzEMac00rFxjlR7cAFHp43S1vKQ4zk7cUGcwqQKBoSnpNWEyrizp
nRNE+4spq4cp34zWhPlCJa8KsG+keDKP3wjZ4Aj3hY8FGGgo5/eb9ZlIDgBhQ2+l
a7XjdzjjxhPn5odeok0dOPnKy385qSA4qM+pa3LHflHskpRGAMSUhM93F6RAu3uc
qS4OmXbmvyMMKnWpJO1OL8CmnobdffA6EEeEThBqizggL9vq11YDqsDoi3vTjcmV
lB4bbfWrscuwb4Je0DJ/rPE0NjoBpDJX5zKiNgU5N2wHF4hN3n0+0b1FFLu7koFw
76QqcAiN6VCDUUzTc3v8SgD6y/YgW13CVId2bBE/OFHU8jqKwyDWX3H1f1eh7HxZ
+qyAuOG1IdOM3u9ixj0ukK7jn2j70lXtycsu7cdO7c0Mf4ALJLyoiTQQGU9sd0oC
RexWuTCKGBYnyLuZsWT9OGghWrg6I+Lzb3rBa5eBfhegHQgiAOYFB9/I4eSMmUto
+S7NcfgxVEsLFbmE9HernGQYQw7ZI6rmAmDpZJW2+8ECV6v5vlxFEY6/whGRIlfJ
ofWwY6Mg5p+7PMFxD7PdnpjceuQtfkfKmvo0bII6MSG5ivlWqqUZLZ9vdkU87A4t
g8N/enw6tc/NuqfWjPRoKzjV3A91Rr/enpmDz8RSqrFw9pCPbtAzgQToB5F33FAH
Jc3ue7hf3QDSUVfsMpuqT4qeTFhWKOefKlV2IAA+U2FejnaKsc/XTw6O3LrlKRg4
sQhV3ukRJmvFRK3vkyvJOQy5mZmBNta/srHxzJgGLvUa3ZJpaf/IdJgtch6WNJWj
rrJ3xWPBYormo80QUvlMCsaAwYJQ/6HhaNFyCC1AY456Fs8ZGavYGWtvWa+57dW/
nPlzX1e8TjZfpqos8jodSF2w6u623C5UWS76W5VOJiPPibVnKADgs1tf7KCHbUyM
gpDCLvt1SjJh4kZnaMWlrTxnr1zxzlcaLM+muMXCHh/fAZvy0vunHUe6EHcQ1aTh
A6+LduTa9bHCTmSuDud/q883JPUxfrIyzxmFE95gD31IHNTAQcQ5+bBmXNrsc1Ab
EkBOwj8MhpXc6CE29r1lNzvDNC5JzukWjJyHfe2udQ3RrCfOIXurIFeTcLKKHJvH
fILVN5+T/PLkXBHF80xpneFN768ma6ylu+WP7QEOkKab4uxEIElXfP0te2pcnqXO
t68apcSuF3v0VOjdxeSBoO/m+jsZBeTe9SsYOxVoCLY6WaeiYsT1+I6KCh0hF1pW
tM4EBaE6FXbbezIax2p0o2VKH02/aH0AgvhdgGaL1uGzVZjM3jE2yckk3s4xkIzj
Wi2nAbrP/19MEQXlVKNm7IiVVwMOhENXxCaH5wfkeq2O7Dafx7TVSsCr+mpxTmEf
KOTyilA/zE1F6Pdoilj9g+n3EUuvSNCB95IPYi2QtMkmMIUdprsW2cL7lUwo5mkT
fVrTzi/Zm3alXpFJLLJPUTVp0Q376vY9QxQg3tVRdL0DntDkAdJ+vRfputQNHq1r
pI4BVJLTv2mXJWhlyALuYTFCM8YPEH0ce3QC6cGo+I63RnnE5nieIDmH1QdpXX6b
sDKzItcMhf6LpBgZlyR/hNxVARh7BXKnHZdml5UQr/BnxOy9exrF01nJ7E0aQEKL
u6TUcZo3jJVvxB4gTUqbSkuMyM1yW96vtoCGICJH15wruGVf4WOHtHAWDgyD/29N
k8kUBPX+iTRFIJDJo9gry+HtFlGWC6Z2LmH13UgWRmnI/YB8LBITHYTcDmgk7PjU
URIU7SLrhofYv0Y0kbEQadywTMdT0tozZ4DptBwTKD1Iw6/KvJ5Co2IBptJRBj0K
xQhryKIlb3CWfOxY9X3Qfa20AGTyR8DR0lKs6h5U7dUEMaQKwT748BH++xkcLPJf
sQ0bb78cXybGRW4aqxocLOp7881Y9clD/1WctU0kahYprgQaxX9YTnJWdnBOjtA9
DGj2xppHhYHMyxAbsIZE7M6yKXQyg5JMwiIEoh3gQVIBOQdZKEOOyIkIN0gFWvJp
amNRkvASG+VdkDHq25yrqBdsHyHNh8IRlPh0Qs3nN7XtdywCXojCOb6avsw2Fm/W
C0b769N3gHkJFmV9GeUTwbnl3iTXJlCjF6Irp/oOtXb0u4of197UFEhWv0Gz10DR
ePWoaD24Ec6tU3aLmFrRqtgIQWnfh2iln7g0zgejP/HYPAwIGLUJwFZnxq8fu3gZ
PqYxL11nFm1zbxmx64Iimv7F3AYwVZ+xadNyL5H4V+G/b73y93NgvH+XcjQUpsJB
k+AWl9jD8FqbK2ii6cBpfKE7a2Xfh6YQwSmswGL617Sa6XCw5UXlK6GUX78BqVLf
aLHK1ysyol+OVT1LOLwg55pamMhxsnxSOQkGF9Cjk7qY6mJPnKUcv6dQCje2DOn+
GdJs93gMQn6bBKZY/UzpvASifiuWeCWRLzzk1hjHO7djrqp0UTK2t9PA3axWGNvM
TATkvHn0sRHJ48WV93AgbG7x1SCb1m6Omf2mVVDbkHkwJoMGru6bnF6AFdIvO4Jq
Wu4UZIYkkmx/jQLzzxjZHhXNK1ErLJpUjGxuw2C9Ujz9Tk+HKpz3smT9vDlfFiFO
imoCVK5S/rompR3qphTqoul28mojWwk2ppHskflbH3SAp8R+ovMCZFMhrev1GhRh
fwprICPL6ltuC6etSYRinPyOdB5cH9Q0oHlakT+V3G+OZ67HbFGvNF14jIySJLHS
0LJWzlOs8CZwYJg9u3pNLQGuI92EY8x8gDdsgZPCWsgq2rQlkw7xWjknVoZ6Rl6l
Get3KwlRMbBqITtY6r7Cy5uImpMTwB4id9FuaYIJXMdmikDIJm+QDj1mg65K4uBG
FZgZ5jdFxXf+O9yXP4qKKK5a7S0O433RaEgNDjVRYVjjI+eSmBIpL1aD3Urh1YEy
z8Ujn2DDb8al5QhHa9agE0EZ8RA4HW91q0pxSmV2zKXQNDtuauskxx9TxbQsiTwr
yLx9bx2GQnf9KYs1Pmuz9yWnjH3Hy7wSjAsT3NfM1mId2GGJ5mqm2yWtk9Ty4IHF
8IFaWulsArEBvHVneZD+Uir6s7uot70CEsH4C601MD6JbVVdo1MwtH9d+bdDj0x6
KlFf331BOI1aZukDsFpwW/uBhThWXmMnsq/QoaphmlqvaT0D/fwxncRCyV5+Q+CT
y01u6KZeeM1LJZBHXnO34Ag5OCWckP5mkUu7k4LTh8Jc1NRbK4E08UN250ghTwyU
rv0kBe0yGXenAh1D/aMqdWU5i8FOB5pC2SA1GQfLAE9gfDW/UF2E7W7OEIB3iDsx
35qdc0qJwpZ6Gf/l04NmDKJSesjvqlKS5jvPRhBY1Nh7vYuGwJG/veFOMphLpOeb
jz7fk7KFYJ6VxntUTWcMdj+HU6rl71qiB/2iblkGBE/ZH3IEgif77nBQHdOwqaR3
vUhaUIFbBm+PkWdyiyjBQxb9fIQQb9FuHmq28xIhIwJpD6QEjsCKhVt3ntD2ZJYW
QSQDQIxpFnj7LYjvLIeqxAXM3A2+Z6i94Iw7TAyrOYV5J8pbmCJucUfmFwh2hD9Z
ux2h+wczxmObU5Ss2pFDhDXjpLjo8s5BsoD5TZbApNzQXnQJJ6mBi4WS9rYYYzj4
DvKEFmAG9Mhdsc7ggMjhfW6HKLUPGZpixhRFuCZjn0fvvpUFJn/JfTe0Ms13dbEB
AObvt29ov4BISKg5GKfV3iB8N6/WRrxuPzgAh5FuNtN7BOC/mGOPGQi0Pmay5YzV
uR7VFuvfwaZOeLXn359zDC+OQa8d0eMVJ8Qv0735uLMpZmCEDhQDitjjjqSYg74W
aPzCTI6hzTyKs265uc0v4QhgVspdpqRYx3f1aEyM3KEuKJsCtpTEVLi5QEJz7Bul
gSaMxY+dJv21Z+5jPZeQihJLLnhcvbOKxSyrmkkSRjXTMvz43mC+5kwM1Ck+i8DM
GL8Nyi5wYb3Bweedi8O+qv0CBrtqLq9I+TjiM4cPE2Ol97oqosmSq6E0lhEXbr4/
pBoNOyfIlWLz3hCO8jNd2NPLJN3bD2xjAsLBfs4/lfhnl72qC7C0jkCNzQjSq3oq
gTvlOOqeD8JiqeZRo2EsCr06X8k/va8NaFC6YL/7dmEsYJrp0NbqpO/0mzg6SW5f
opi6wE1guICww+0x5L3witEaUA2CoHJST9KQuDFOePUUtxc0UilMWCnALXgh1X8d
Vgzzz/tgSG7Jm5bK0EFP35iBN8SRFwol/5E7UpEEHKcCQxL44cBd5RpfHS8pOV81
Wd+3hmClMPzM49SsqAzkG7I4lVhZTJWOgR+d0GlwiWzFu8c6Zt+a29rx0fTudLfj
gxosXVTwpMoqrZTSledDhXE4+h7kqcqDmHfsPucasJg8eN5MACN/jTm0C5hV3rdx
Pgd33fUXsaN7rUclSZ/H0NCx8lIP2uCMnoepS0Hw0tYM4bizCzONo/Yt1s0mhsSr
nlZN/GeE73l2j3fyf6mo+ZJ4RFMxzSoZObOIBwsVsJ63oal1q6Lv/qME24T84E2b
biyu67piatAc57XmctqCQ1wJl6ePD1xFOQsTba9sqb6e1N1726HO50YC9ws1Si7x
O5OTP4k2rDLnx+yysJA+Fp3s8aryzR62q5S6Wro0uSJRyoBpPiPlnZTlmmfLaUYh
dD76djaQ5mSKlY4urQ7/ODGOlz9n/urBdk9LX4jLFdPIwqUicEP2R8KBto67Lhum
HtYQN3JeGn0E9876Z/mDMXUi4YUvpuFZGk+dpGHZ+wQlaepOIxJSR7kbLTDojcd5
KsFj+zFuhwEGoamsgggQMwi7onM8FhgB42cL2BXvfOPQxGPc5zqqruWdWj/g/aNb
i8McTswvzI8s9GyIcFRU2uq0e098Wk5f/ZyHqp6MLMLX8g+12mrPtaYKCO7u3wPf
UqsFznWVZL+ogeRmXlPkSGgqqMUBCL7057CeffCuLJycD+QkdtXDTVFoYBwUhjSi
e9HsgidBvkpVHw5UB4xR+diRMrCZg1qu1TrieqWgxuAhJgriID8Tje52TuOI2c1Q
BPNTjm4dV/lEVqimg1fAMhbhy3q5dL03guf4ad6J4mP46qxXTbtBhO7VYkXc8LYy
WVmeiJh7vBAFwTy+XN/2/N3AtKvRHULHgGmbwY3RMWdW97MsKhXf76W8eI1uDZOg
9wBdOAgjwOhp3C3a5rfN8OQbV7md+5zKweXYaz2dD+Uf+vZEOxpEKeQAOj0DVs8g
OWhWi/IvoSJSZdfqbACOAqLZxCObbKZ7gF+4WldS4wEvGAW1PU2lwRtzbwqcQvEr
fBNNu5zGq4thYokWSs2epxj9nIw4k1SRYA5vgxItS952z9+yacamlBm+Bx5/H7NB
tEhEoUPXEb6xhOrplk8HeomEvpTKAMHTf1ivikj8HB94XywgqT7BsE4QI0UcABcv
r3S6m0kN5cwDBKsYnI06pjYlvco/VqOL0cfIgb79LyOnTFipM9cW3bO6mqnRZEW2
5mC2TszZhye5MkhP8uBbW0SL5KI9xiNTgzUMhWwD5q3ESQX1aqvs0Az2hTdT5zs6
t5LuLEXhoZDjDacZsnMctLrHZlvOJ1Jkpfm5bCiWchXfwPH4kKPlskTd4e0c92CB
N2nj/cvzhx3v9ZhtyKsVlfGgwzHPW8MwrjQ3PqxcyVI2SqWt5cm1pNCv9S4kO/Dy
kfzpwHoe5UHi6VzrR25NU9/3KlpNITRmFPkxQZ1iqq56RsUNpHFbXIbgiL2VxGUj
qKHzmORtVz0ccO8ub2Xk93g5Y4owOTARVdAlW4/jTJlF0WevrBA2YcojI4zWFrzm
/wrr3kb4UN20+KRFiUraK/ehgiO5QLpdoOHmMjWyNFZu5/TwvWXtu/8MCiPB/mdP
nysUU1MZmTZj03x+57sLBOuM0v86Yzd854TyD+1s71dv60aBpEqIzWbkRoPBl2RN
6sUtah3UYy+WNseh9B6VDJgqMTjX/748RlpgndXPnr6PNE7sv8m+oApwUVdTm/SJ
jKlxqzNsoWBNAed+0gmNLCVhR6jSi0k9OIHhfBUGxhvUX+9Js+Ff+8xy7G4KNXkn
6+fSVwbau/YAbY12XbU4gqyOFldXGXOf/WzwRjdsn5k2JMRcJ05lBfk02YZ5kEF9
/BJ8eMZoMi3ACuET5SZzDJw48TejIjWZGsedXDfZdak8uNBp/5Rah7skN863lp26
lfj9/lYDPT6RH4JEJoVpXW+FPs9Nka7/pN4X0xSNCT4tN4VmfgjM/hLuaEFjM9Ky
w263ioQkotTK5/RsNGyTUIyC6QWtCeAs5fhbLiRus/nm3vjWLbWaUkViiotJJBpS
/HWlaWJPvEoC67eJBZtcEo14Z57hYSj6nI/dBvqOJ2gQvk6nX9/uWlXfp1yaPiCM
acBQiYQcFUjuRPU+f/UQGIMccY8Y2lNNEYoB8nMhcoPfoWt5z1XzcMQ1YIdEvOTf
iTTmyNa2IL+ik3gTr7kaJFcNuvI88hxyvXtcyaBAXOxfLG1kCo3fDh8gLLG+LeZy
cEsmMBiE3JkS+/3eNgK9uBR7hBnT6+QLbzxU3uxKg13oP846brnxK8ZXIf5MWSoo
xa9HZp6Flg0aNAUraSY9pY3Uw4CeQJ1rIBQcZXxNYZxTtlRehxae5iLDIKFHX5Wo
yolUdCBRF3kPuHKR0urMnNmGALw65j6UJiHoH4si4Z6pd0JgBjHYyuzTnSGlsFrK
F/Vkbr1/2OC/rB/LXU4qc8sdH3KPvz+H6m/hXMPXGV6AhZzMvHBPWVH8Sjhl69ST
1qLdDp478f7/pHMduMQBuLt/ZOhHo3g5/GTp3gpl9HsxIrWHUs+VCJw7isUPRiNx
765LyC7OIDzHisI2InRieZu87dyL1U8EPHUw2/2rn71NI4piPFzxfHdqxVJEtDRW
N3CpRmx+HiN9EN1ppiyJY+AefkFvZu9cY1z7ejQDHG6Lku0XbtE+O/sHTGNVm42c
t2fDpLjqumtrTA+7mfkP0xlFt4W3OUA9O/K7zax7ocglT++sXjs7WFC449zWBjW3
R5KSk7boAQhliOfMrIWtzmCd0Fn8yYenBQIakyoxU6/PEYYyY3hw9Ary3g2YFj7L
o9J5Vqg8+x9HrHM/pkbJHt4ljUG8fkZXNcY/xyG1ridnDRyG3t69rOTrBhx1YRAJ
1fH1oHvNIGzxhIGO8YS5JoDJYTvRogAiCkMUvh4CaZHaz1SwrJSQ2QOPJ6huPHqq
Tq2Xq14IfFy5SUx1kmI29cQRkZGCRI60Lej5pN1kLlzasYVeiqaB9E3yt18+CPnB
Rzx09ZYbs9hSPlZ7X1lUV2BVTSb/8JB6isZRhP/hhHxnNVGvKzFzs+iacQY1wYvA
B0F2IkpaNZabfMOkJI4ay9S9jDbOUwJxNHSluN4vp1ii4K77So0G1GwnsUULzx53
6A+z4Hba8yKSLc1emGu+FFwx1zPTEMi9J+GgpElr3CDHuF7aHZ9zV938qFfQoGMg
njBxLekedrBHkE+NCcNvxPT/gzD8Z+C4Dv8IjpUkx9uoCeTMqysFhDlD6Ee5YN5I
K7NNJ6aK6MxERSFMcPG7FVNe8FmMyqRAVrUDc7IcU8lmnxFAmNbKcG+UG4EpFAwj
armmtCAXVdG40J2D9/oDG04VKbPgJ0xII4u5Da7CytRVHrmbkNh5Q/4qW6FsXSLy
8cbcWeORj0eW66ScJIGHrO1xdCmrq6yr0InbO+Ygq2hYFCZydpsqkMfELKjUtAWx
4RzeCulFc3LICBvwe7PFOq08ygsGZKlZGfLF64TOodBXV24sjNxL3vxBvfBwVw+U
NUaAEHh18ioj8v35oft72LT2EzWTu3OtQ+xgZnBnH+jxjNRyMW1FHmp1fexr8ZX3
daredyE/7PxljuH5r5t0gqR/0UNvqkYsZwe2bhxtLOPtI1bz/GMpLH0EC0my7GQe
9nIsuOCcqtO+o6HGZsC/tz2UR3z6/jz5dcvd1fvPUuwqNElHVPY1gZpbp3Ms0eX4
Dhdb9ZgDU1lo16pkRkg7o/jo5erixAxX8fvzNe0EJ4DXm3UrnAiwUmwrEPEUV2GG
0ydGLklrOKSodpAprR0LeOM+5R/2P2CMYGjdyFuKjX3KnYmfMrSEuBqYKPdr5EEL
VB3MvHKHb6Ftem1knNVn3P2gdV/ehXKW/mW3cSaVn65bnvzzC/QjK+weMCsXub2/
ab4kuo8ffcYhBeczgfLPyCtRVJcpVGxnN45h4eQRFli473I9VIHFBFEgKEpNUjVY
bgSupCRvyxJDMZdgYmayDmPvVZ4Hi+fbzQXIM8mad6KTE4hOk1fnoRmSUulizUvi
NHbaIDlwRQT/RLR4UKtcWDJaB/CIQnP8Ygc6wB8csSgmV5vOlG7mbgzJJrAsv1mH
Rs3344P8hmzcH4UlW9FAPny3Wxb844zT37VYflXypKn2rg7YFD6wqo9RF7YBICiA
vd4Dmpk+4U+e8vIa2/VASrUBTUI0Xt0uRCtrjYmWsH/lbgSTKKNDFDqMjHFjeoDy
dMUEEGzqY9MuJqTXmBPnKO2eRJqo3LtIps56iwkij7UXhOaEF6wc97OipU9qDJoC
jq3UcPffl2NiBkQb9gakmBx0VLlgey7+1udBiJb63+OFE/1T6fHfoZ1IIKG0TnHD
u0qEEDoGNk9t+Vcw50lYKvfNeb4MLQ85pcWYta5z+EQdwtLAX2tRMNnNeV4xdI2C
iX/g97uRVcVl0JEjTOVIZifbpW28HY5s9bhOpJtt0pPNcUwuLhMfw0/mW4cuGEE1
UtOibsSsJK83HGhv2owCK2NEw8l5RpgGd41Eg30cIpZogRWLqLjCsAs1B6FjlC5L
X3wFN9qx3BdW7+6pX8xxTyYQ7ThgBKIuFln7DiNacd0pN4avlTgQx80AI9JeKJnl
1bVXAZNklzhWTOwIq8rrfzsGQaXU9jKHz8YGS6HmQY1DVXbx7hqAZkOcf8FcsPpf
cvppMNC2CBttibH7bmsbStrpMMYu8SE/OeclnDDNwV2kRRufkNQXitk5rmI2WZB2
FE79WZr2CPQnuSkBjVCuoWFj7d8qjfLzx27kkloapavoJ3DYu9BTEpAQQc8B0H7B
oHMugJA4zbawfXUW4ItsZw2tBq3ETUMjpQ7az4YC0JPirZ362scSL4zkPMvTPPGQ
XyIFj1kX1Ke6DoovCaSwDYqYKXOfAkjZTutDNWik/gbSx+ltGmkAlnAFekIq1OrY
pzxZv3ZLMIivR08vCbWUdVmCQeQQBescRmPq2hdlFXuEMimOcTI6vNGX4mhrj21K
T7jZ95gM0oU7k2+sSfMzjaOyn5em84nJ08IV0Aj6V4NT+q4H4CAELuyzU75YYXUr
dkqZP6O+81RD4TAbZ2hGJ2ZZS6/bZyPbIhcUGmyvnGm5Nm6iqNJc/qlAfiZ+gLuv
jfujYIZdphMUcvkHuQdq6LVBZphlYzCyp1Vxn/PVRHfRpVh1Bd8kPOcutPeziGmC
Z0QA1wm9q1GuQsVszzjUU0or+6wc2RklDAR4+BZUctDsAQJUyvqZI7gnnGFRxy/1
Xoto5O8NfQn9RmSew2Grtn3J/TTrwjQvDtz2hF1fNI9PIrKzB2B3ZJAQEEyWLnzT
vUdZMG7T7jKsa+GjOJwrkoFRs+gvSl3xQXUOUWjZwuerNlHI1sd1Ouj7nk0A2JwL
OtvtygzxogJb6AwKEIb5yDWon1LF7pIe0ObCpAhmQA9y5f/U2zyqMUg29ldiZf88
s1r5fXDIa8umR2e0huM5OBfpiaT4Bq7buQDq/tdNZVcSaPotxR05OUIzG+SY/X/r
RGn7SIb5TK1pjwgtz0BNSRD/QVOauvbizAjChqPHQTQ/sQ+V+sPToInyIVH156/X
KqiwWDWLayZukE4Lh5UEWOpNBMwbfgJoVLshE7tit3WcBY22YPrGXKi2raIxbMGx
xbNeuuaZSTO9XHbtHaU22p/npWsuJelS8KSJRIgAMyzeTzLCHk2U3nJgoVV7NR4n
Paf0ilPJ820N1x2/gwxgvZ98/R+wE3td+/BIrjX+ib6NRmLCzPkSjJWVKtcRwyXz
Mm5QMmNoJ5VM1pEoVlVdEWAJwf0ntOA0TN0u5QMqrppAjW/ovATrtJD0VUSOWWJD
RzIyhlXpIivSgxQ3ENqRbEKPYJnqrtNIy2N8P4cqbN4fpOYucqpmM6xQcZZX8iUU
62JqMvy3BG6q9ZY/zdLmJfU70vmv6qy6kDfBClFp8scVzta5kabG62J5ONWVppPG
TL2VX1XLAT8hMD15OMrkkFQSV57l6IPEHj73G1x2H9iJswP7XTxKxQet10+n0PiJ
qNIUgs3v5+TjxXsazwnGlLa+FPHhsobOSNWtmNhHuIXhIbda0k2GRIJ8Af9YlWsS
fLGWH8DKUSYZtWW8h0b4f5wFvlJr1bFHCVv5MeYzXwlF5YhOZnVcptUT9Ez9qL/v
6Ch/scfO34TGVbTgmCwGufEPtT3E1yLe25Xy8SWQNhsAI015U5LmIVUhQWa9XykS
8bDJ3L5slIe3ndsOBBydOHpFzqkCtjMRGNK0xjTD8HYY0Ifjt0LACUVEzJwQwSGr
Lgc1QEc6iNtIzIiCMw3tYSyIIWhtuBP+5RozsjtpRV/mJ19hIgoBxyJKF0mlU2Oz
4/mG3hI/zqXaedlPV5H9ZzUnO8kWI5R0bHh3/fW9YYgSqeHQq5RsTn/JPCbSZQO8
mIYHpVzFvilQLDwLbuMv6eICOkqAtxGJvIUgaYIYhUGcBnTHALRRA7j7FmSzgiYs
Yc7UAchUXOMYQll03IUbZPZlriJiDeDjq2zW40zAGdbD7maywpiznhYYvUKx9ds2
Y4m6pB14NSfp4siDPvIX1sPpcmIbF+Rs72Sj16SPiaSS7FkZ0H9YnUKs+USmXobe
Xf7hl72fuwSlU1MC9uRD5IdhhDdeX+yiZpoq0xbcIy+cjv/MGaA1/c3ej0YtKSlE
5flbMKOzTWWjIsJ86Cda3SHZIJK5T3HeGLR/S9n/RDiFH/FXMokxabR2i3nUKozE
NVhV9bE2dDQsa1EKcXZCF7RoYzIzArolF41aJofp7b8ZtAZlxHsK8jAHK6WkAMqf
sa7OiACSJJVYAZikvuH4pdQgClSaIJa5kW9uqGktUepjRgCAY4QZun/USCTLH1cg
3MDlbVEgYVCwjiJN0Z1zOzZyhp/IXGSn8QPnJEeKFeYTySuIVbETVJNl8H00X7vL
ms0ty//+Ev/j0FUfibX9tY2dcB27v4VCRWlr5GMXEpTFvuuNtUwMGR+63UuZL/NM
YcIKgxie1aMVbgVk8zaBD1YucrNtd/JZ5S6Qk+NhxRUXIKhqSRC9eMYuRjY1MX70
cp1wejevdW8t8bIgh9DmwfHxagvB1aKe3+gd/O9oWTaiXGjqvQQZuxiITWSpXxsx
C0q3aneUmXeo7TTYMaLkv8fAswa3qPGXNgmIN0C1JaL3CFjlllC0h6aJxl+bsVvD
M4RxE5pZKmH3+xYvctixESmQ/L1CKOVCx+v8GrA3O7q0l5QdxLQceo+b0imlfW4g
Qyp8wsH7tdcTwsGXVLvmDuhRMOWmKc+ggdWRJD7gwjQXIqK2YciKKod+ko+9Q7qy
aoyR5AEzD36Yl82CtL3XbjXVnpAzWDXvh7RzYI4A3stxDCAKBzLIdDn6gyDb6/2V
8tknIak1lEq7GKncovggbELvc8SLbWIx7ow2O1fQdDA2vkuuQ4tNduYjGpuB2s0H
Acs56YiTKXQTeMM+gPJuqVx9JNR2zyj1f1woEKOjIG6OyAvq7NIhOTJtd3EsMRHn
CY4FI05w+qodESzRk9BWB5eHy7/TFuvl+6jXApFYtmRfIG5X6d+cbt97fqMpobm/
8RVG3UA6LxIr89lR2OiIlt5jcAenAtHH3ogfJfL236i7MwZjKuJLCZPOiPAKMNWz
wnPiZo6sfQ+rS86CRRT9prpJ6P9RSeWovmocIzbEH+NrnNkfyG5Iu9SPwHeCZ52Q
RlbTJWmITenQ/77pBkSGC39YHoWJ8SrATAkbRoh2PixmoYHGeZNaeZn7VmHhQnvQ
KQ2rUwjjy5ugyeTZbA7IWkDoJnCJ7tNDWQtRl21yJHH/6COVXDJe2tSYdRoVKTzW
xwLfW8FBZBqfN6dHwzQLMro/cC0jhIPQ7eUpLtPvDOuEWwrx1qd/u7BE9FdY+omU
K+htGv1HUBXuo9nf8IzYTYzHPWAP0vhNw2sc92JeRCEtVPbat0ry4Id1lesgC97e
A4QTnd9BktXvsVB72095ienFY+0rImoCCr/nVu37cGZoxaEX6NiqXv2Q/MWuiz3h
fjaDIPLWf48IJ1K31LlXsyYFJ3gpTDHFncIXMVcwmoyllfJYfSlw9woxf1Kv4StO
JLqTJ7pCKLxQXzZ4/2H5CVkm1iwgR375J3NDB5vi6i6AAWE5Z9iCZVI3dkEYNqPH
a5cxGUTx2FX/2te/e+5Dd5Ke/O/JF5qUirvd4jANzvjZ5CSml+1FQjaflQ9BZVzD
qqUVd4Fw//kLTjSeQ3MvbDdEAIgCYtMBV6JUdhTqkKiQxzugNMjhE/GQBoLdfUS+
oVJFU2fyN3pgfKLFe7GCSSooqf6xbtZLDBqyx7c8+yQmU/qGoC4pvWUClmm0rku+
pthPl10sPVvo4rKTRZL/hgBRnvikf3E15GqywQtg9vxsl66CWUd69JWMzYsKu0we
3utnzFUAn/IihW1crll4DHqQnNUCHhCn42zZa2XQuMkzuXUgwcxMo83cj+8nJ3PY
rjpSnUbxAk9SE41BEBsU9Q4R97LB3PtEvaG+v2drrbu0ZTXMwYfSlICOt/TPg/3z
mzSj1WWGLDAzAJNRjp1tc01sFYV4iBDUELx+5ZH6KN4Ku/eXkMWuyAtH/sEJgS6k
ZJGNCz8fXD+TuGUxjvWiyarmaBeC7W3OaEWXj5K8i5mUFwVYYsezwv6WeCbjKB69
14qNGmNbx45rH5aB8FnQhj5mfqoeOtRGV5AOtaHK6aWa9gmYI/YcBsrMYOTOTMie
FpS85Zf9670LAI12bje6RUjzjPSdSbO6Bm0Us46XBs/fKN9QQdegoc2Um5lkG9Vc
NRiLjL20LqysAuNLL0sTaH8sJay5cPQhSKzYgBjMyvgKOjf8eViqQnSX6XzRdJsg
2XSYpCaBhKJKXKv8MtVi7xmBnNn2OmQHqbgIodve5zR5WZeRwTo6id4nIKyMLmTe
sfhlL/cRtdzFqzlxykZdZMDA1yhfybC+UbZumRy2oEVoEuL8uBcVxfbwj6Zr7Ssv
0NldKwNweiPlPWXwx33jrO5LbGRCKM308zXSN1MLn5DadgdkYJrFGZs2Ry03fvOo
ovyHqto45eWRxvC9cOgoOWjjUNQnvxnie/nSSG7a7wVnN08/1+JnHSXkuKOaViUc
navJMAaBBqB4DjZoorqipZbfc/BVstXSVdHqkTyRQmPScnTH/8QgQbX41nbPY6OO
vIkqEBtCAGb0b4zkiNGZU1DEZa5MtAQ6I2BdkDaJrNFMC9GCngy9+SQJr6c9lP2P
44JwAGswYkTPsslvnj94oiIAlLTYECCDLhUw1v/kBcqZM09DSsnsRkWO2XG6mHQd
MEoRe69T5KXT+peV2DFGS/3BKVEHQJl3bD+XmL7ciS2z2c4zUR97KfBcqxJxGfM7
k59+bLAsZUmqbzn39CDFOvvoXOCg01jKotdnnxeSQsrqUsN0sBcEMPkTmi6FSUE0
QHZjMEjyYMhyvOmCZ4MjWAqs/FEnq/Ub2jZdGG22J23yBjp/oJLeAIhb6UxmuLQw
mPLSqtC+XwOwpEQdTXiTzrZheQRkcGLFZ0eENqF8fIi15wa7defng9SIPS8YH4we
A9dtJpHhqSK+TOWssy2fDyS+y7zYqX4jWv2AIPZZvKnpcKn8b5CuC+MEdC9lQGCP
fyP6wKvVD+PgytIJu28G5d4mu2oucq/u2+1DpPNJhZlPzFOhIbsY04cb9D1Q18c7
Wlv1LFhINFBX8rV7tP0PktlqB2+xNmfMEbsqenQp/27cAph7LhEPYcwsMrAcBCCZ
gHoTW7g9UaSg48CPDnIWieD8qY5CZWUpfn4XPfXsmQnrLATpOxGvwADR3GhpWha2
3YsI5+dG5/Z9QREGpx/TwGUuInhjtpv5BkOWNL8vbGP0+aPMlCaJ+QLzJLGH2apX
LUdP8RkIFZuVJ3Oy+Mh08aX7VkrCRmNTJ1AQW6K5slkhwK1/Aou2lD5CuPKwhp/p
bwwU1bp8jbfRcFbFFRRun9MIHzzhbdw6CcnJiYBJ31gksWYhk7Y0mH/49EW4dr4v
FbHuVG4slfQsi03xePefy9slubuyJkQNZfC8VAQ6VFqh7Nma7WazQo/mJFAUYvbN
dT3dFmt4IBB9eCOjhAwZ4j9H7cS0mvBUSRoBayWED9ps9wuThkjQ89OIgnCeEa3c
LNQE4QfiGa9BtgEqwn3PtC6Q8i7PGHdQP5zfO60rt6O0Yd21vmJlxHLw9K2WsNk/
I2jSx+zGxMx/r2nFvFvKfZc61IZ3PeKBn9T1vIsBiPgw4JkNYWEzFA/UHewij/5p
xL6viRjiD9WUXtAmnpf+BA2hVFcP3kGEI00wtk1TI2w0n5VDhK+OYDzhAqZ6SuBu
WQnJ6iBTFh78VKKLbsv44Lc7JsKEcbCNuf5bf4DABxaa866fuw70ahSz5XbdkdfX
XseCF7tRd/NeDPsgCo9felDnRn03UC4twyxZ65pLAwHg0FDgDF81frGKwyNxNIYw
GfW35LwjYJk9NFjfN0QayHwRtkIV+Rpz3yoqyBkGLNUBDegouBmGIlt4694ztUNC
BgdvAwS5y8cAwVwfR6APBY5OJnu4xfTJJx72VGvUm+S2vD9rUnwnnfYDU/M2fu7K
7AYnfpK5pA4dVKNhfOfZ76cebpXzEqk52/5cpGGiBFIbtymLs60hZHiI2n5Geizb
mt19dqlGsg4R2ridrJx9P1Xpl6gXxx08AOATS4rgE4h/E0iFgt+pU2U9PtxqwgDo
8uk7GF1eVJ/uaiZijCZcVzjgFsktl+83/GvbstB598Zjo29NDnZ0h8L67ZuTCACE
cscgvbk1+sCwgP4V3SN8C/IX2PdgWSQNrGeaberRv3+D853sODmQva2D0TH2JoHK
Zu8lbwRV8+O9kwAV7An9HIisSVeWzDBfNblm0C2zSS2ttzspxtG5KZceqA8HSggW
IS5HiCUJMnwdgHGPEjj9EqMNPe733u0nueD95uTHgiczihhOQTFxYlIk3IH/xmZf
tLvlxI4Zk9l83LOBKuMORawsJyINbQKdQ64TFvakAWR0kMU7KMyHSeQAKqAkJu8e
Ps59gUgHYSivSyX6831079RztDjvigFWkctIKpTM+2OYW9sjTZyt/1a2BTfkTqbl
yrCTUxaW+ig1F1XUUwobeTVPQGaJ1TiFbnqj9Jr1IhQFscYL8kDpSBRka8JUmhJA
KufPPo2xoFBDuHo9ZFjEor1nnCrpjoKu5TiEu7IGZG1DKIEUuqoLGfX1SDC9ECJj
8BHYVNBuW4hFzavqBDuzePNjcUfvpAxWaiVa+bfiNOV1BFtjhst/REXb4PsjeK7w
ohH1XMcgKcEZkgpZP2m3dH7917BBo6QkbtEAPQzm4DLsrxNGOipXRa/vdd1y3E+D
WjrmrEEh2jThR3WWYkoLy3S3L3KAJlWYbSlPos1Bqz/NqibNa/n6kUf5IrkA8aN8
iF9iNFyB8rFY7cyDDEvyDBzfFtKQn6zJb/TT6NexKhSu/hDFVAaSaLT4V8lHHqta
5x4j3O9pVaSxqAFGMyoHxAkkj/THqB8D2KQt6jUFaX9f2LLkfwe50kDIEoNNXpbh
7lDjiFyRPPd/TCEnWxfem+qMypo032pE9ufNaZbhLUTLXW/ZA4I9xY+pwut2i/AQ
Hq/9KzGobkQgf0tbPK118rtBPpgwl3CRn+Asa6xCCdyES6RaRqUCTRKT2WCfyrJB
wEXSkRflhkwqvoc8NCYDNbLCA23KOP8cnVIsrQMZyAgIJSCXQE/mVvleXE+Jg8a6
O+UZuHCi77SKWpM4qxiVxwXCtGJJyAQrcy15lN9zk2T1I5ALbTYcCWRCsYkDjNY4
H3HdMgz+9tc8ZSkksHc+zw1hkYfKNfGvU+jWI9jMWtlaT0oM+ALSepUD9n+xIFHG
bF8vgHYBcLMapc38xSWCYnb0kSVyqBiyiWeMa+JiqZsb5W9Vbr+y6o93tN2Egpjb
FB+r9h/ZiXh8E0681Qy6D1yMSx1uuA+V/WzMd72dfd/20tCDLVQXuPizinVp1xLV
dgj9ee+jGheouF5v0RV32pkVVRb9VpQ5xVNek4YmmmcZp96g8bwA83K4jXkgGW7G
lqV77ffDPSqpBKDlYBWX42qdxlsbf4wKiOzMRAO2r5mFyhLw/UGdY43rQuCreXSe
DK3Pzom10Lsage+13ikqLL5UKNf/m38C8yUXXIhj7YwhJuNrfT8JOV0tbU3g74Sv
rkQnGBBJjg819XaIeTkz1Qo4/PuMvLPDkoXp/UiZ/wktRYmnrodKNM3vCDdIwl9p
6b7XwxKFu32xbjO0k4v/NE86diu383Ka+1XpG2uoNrM8Kbd4B50i4rJecLVQkLvH
o3nj8Ovsc0A3+vDyZ2NopZTB28wX34zFFExk7BWbQzgnxjCrmW4OjN8SiLJMFVIc
VrUQkpJBtsXFCKxOAGYuM88oBq52YgXfiIke+Vm25miP26aG5sHm12so6KP0lICe
GXb2EeuIzUzQGXDnS/TEXvv0n6uwz/9MMT4GJynVGRM377PecQc+zimhg/bopt+Q
+aSnlGKF+gs4BGGvlYdU9DncZl/FkS24Kv788rObmUyQ+YBoWmNOGWmTAJGxy1Id
p3M9leKFaaEn/uaYu3z5W/3Qsea2XyhEDsgPYhwTR3UA15YSKQyXu1pCcDZDGrGA
A9SzkfheE/nRwTb0kij5vOFFWG0pYQ709AkWVn2bZA1NwK68KslqJfDAsq/kgnyP
COr4cUMFecvgG9B/BtSceYAzKh6qiYrJTfXHhQ/R0KsWShWYHGHBjUdS10PkKl0o
g9qcgetCnst1WTAY8wie4aDt291lKgy4S9ooI8+dUKELnbp0WgBBiRtX/q8x27mW
oX0+L6Jn5jIcdt00GqyzLig81m+kfjKGulMHJcgkkJYjPX2QAb4f9JfrYMT5n7H3
tkeAzE22YjoJJGviS2b95Y9eOWx80RaJAp/dbmldfWRrglkCnhPjHPEpUE+h7elj
10AiDqKsWShR2nTShU0hl3TlCl78AM+LQIgiopzcZbi2pgiVrTNoWNnyiUbqEVg6
bOC8wXwCi3jaoO8tD6sCtZu5e95vTztAbVcFjjb74BxQ2vd6paAEAGBQ7CRzyaLm
KW8DsO8eANjK9bDBjFc5kWpwZiUOqBbx8RJerWEGdYpRkCZQm81YcNeTYVBrmxp1
BVrWGwnaS0K0GTw0SrBx5w+lJXG+XpMXnzFctM++PWjIx6rAfNkmdnLjf0WD9hL/
XaoIPsZk2DQP6Qk6hYGhPPVMoZ3L0N0eevy9fGGNuiEGcybXLjznFFh+BbkkA/Zv
muPQqwR8ln/LugNf0iQwvZO4TB5lxDHBKiMQ5Rl0U0QFpc/fiv16GcUILwgPwC2e
QPVA5VuvJ1LKHXvghGXM7hscWxUaNlsH82l7VQxNfySlKaO8hLLtmfsWdtjGi00/
hFJ3EglKd7k+XjKJHuCeP2idRqvvfNARgb28NuL8kDTkz2UFaizpsSbRunPZ9tPY
+Sjc0NVr4hmclTRFZNtzHE8vEntWWZM4TKqVJjd+XQtZwmfp07ETDuXQuYz72sG2
TAQga7LLZ4MHWgzrMY1xyq1WDN5a3hXkf42Kn4nrk6YxR3luayBE9EZ4eRmjfrfB
e35kGd54IiLkiIYNJ8PecZj96NiyP/j7sUNK4Q2jpt5MkadCZjaunkKufvwBa1ug
ALpGk1V7rVK0F/uoDj3MwQGMvuWP8G6t7dGu71H4dkWSorYRwD4KQlvHrk8Cn2Ln
axsmXwqWWaBDABaz4Qo0KvhdVVjbAezGV01RDKU2LTBOy79NguuCpTySQ5r59WDf
McSCKM14ccHeytrfmpeOQmeLbk2bQgOgpfljO9nQZnXofS9dpC/Rqk/fm+/m1v3V
tFHCpIubEV28B3lotCYkRgDVSaHbrVS36tSPCMYAU6fQHn62g2QwCGfXe6XTeDPF
VZPkEHPMIkJ3Q/TCucgwlp7ke3i+QXBvhu3+sOFJrtXX6wuTQ8V10lEm1YfPylvZ
kUwMw8WqM2KINjGUlaVEaAqB+CM86JnyQUedaDdvW7gKz2+hKGcgkdwelfsHaB0J
+5WLnuwvEXHa85fGKHApU2F2ngSECtQJBAWh9kw2jnTMGPm0lsx18XsjSXb1iMCh
HYCY7SFdITHP+g/2IvJfzdapoSVakI2m97ntXhvXKz9h4bciM12SWGma/I3UG1TO
Fsl60DFOXoEqdD7HpnVXBH3kCYEdPjz/37Ht4g0kum8vK89DvXJsb9D1dyHAAYXe
7j6eEAqtWQFVIEYJ2IGCuoijT4XhziSwzo2i1e5x89Qp4T4ZT99XsKYtSREHZGvF
bPjNXTBLF7gxB6eQavk/tNDT4wSQTnSC7LqxqvFF8ZzjRw+TUBom1sA26zyBqEmk
qNQG+1DeTAmAEKFCcmokeSOiMcKlhSbKRHEAhOLQGci4Sy+pD7wv5k3GEInmMwU4
je9S1TZKSQceJgz01AZEwnOrpvyw7zX/Tbb0tki5xRuxfE4ToaC/pq/6Rms7s9bg
TuvEovOfVg7IRH709z+7sg1aCi9fMtFVaF+Mqj51zjeqseXC/cv65W/yjAZ/CzNd
PQC2GIpg4NEAf0PTIWiI1N9n19DXfNYMnJbY69Al80vQCgvxNLePWTyhcvukYMST
CYIQsaaDfFyjiN7y6EOD+andY7GRwhnS7V4/8UtCU53b3Lotaq1b7cDH8wK26Vka
M0si/eX7vyEEwIFTpuNKDNCq12OGWyh+IOUpgPW6XT8kIuJDxrjdUxQVOf2fOwJU
Jp0aiJyCfrYvL4YjXH7Yc5flmHys74dp44VL+j2dDuo2rqmwoOmgAhs2qg4flQNM
91yEVeS8TEJ8ZDWUWBIKNWaUjgrINcnd08r94bM2Jw/3uU+FMKw/+OeaKNMTWX25
7U0vz/6vHpNRqevE5sPSbgAWosmEA5q0b3yYHh9L1/JKwhQ7gcITHrtISG48mOYQ
YWSi+acIBqlQkNlnGJlXy6J8nz11+kh6/9AbhGCoGVmmtHWdnyxx2XuwXn24N3zU
/61p9yX1te3RNduq9bx17r9o6aqyRlre/6JrvmC2ZLoXZQ1QpbZPVsIUkaO5oFv6
31MG8v5iqkR4EVYIdjy12nE/R4ycFE6+67ZQygJ92qrYnZtFh339IhEtFmdpTHFo
mUguU3LSaZUBy3EYjWR9AZFzqmI/T/v35tw4GWswPz7r2dgh7R+U3vWT/I/jtm2+
4BXJx/r4j8Y5ABWpeWFsJIYDozAGSj3OxBTkH9D4zujVI9rkzZn+Z4v4QRasN7rW
JN3AvUk5NNc6NJbmglwOCL2OeiSq2czVgVDCZ0EL4is0ToVcqroNseRkYyCftVWs
cLeVg5RcjZW5kLn43kzB7bhgyry/k/C4OmnrnBj+CCx/Qv1HJSytThkkcpLSRe1V
zuqCxeP7WoyAS7wdUoNgc0hLQyKjAd21snJkMosO+NB92GYWHd4vHYu6Uqgz1WjE
N14/hbJSnx9LTmLJLDfZP9GCyB8KwZXZY8MmKpdwMIfoVo6JJc4/cQrjX0KHvRvp
8r5xjGFsa4EHU8p3g+XBm1bSYbAd5mhbipxrrytNNXhEd4OXpITpCiq/J9JpzB+J
J/lYE/FzYJB9qiduHY2MNfevtZZUUUs3Sf9e86ZuD4x0TEsEM6TxKE4LaqMXRB29
bRqrlRtjLXFsDGxtLMG/PTc8AUsbAd2oxm5ZaK8iOBDK9WypGu/HCvef4TxAm9kC
syOJ2s0FnWBuhX6coUpQ8Ccog1CbuyhYgta9J4ZLh5ffl9vh46A/JDCx9SXCC+Cx
NOUDp27G3HpPRjmM+Dw4s8wXRUFhj7XJkdWllWPTnerIrDwVVGOQct8xGvjsgWCU
Xk38la3ApqIkh1eWRHU1YYYfV+/h7CMGmTBuE3O9LFs1qYRk7SleqhKB/wtwxdZE
yjygnB/xJK0t+2oBbCScj+UTACIdAycjS2yuNRaoKaIjasjyfV2gshd95lZgspeU
b5lMs9qom8AqtfbmCI440WpbfPdfWktt8KI0qpysQ1hhdsebxlbagMSgWCpIgbQ0
Ig55LptwkLCazJI9HVYL7PbqsgX+vGXOChQ3sueb5P6d8PLcVa7WpfAdmwC59vmo
FTVn8XA2qLYX5ZGxlN86uJpGCzlOj2i9Qxd60P6d5LocRsJfjzhSXYotZIgL1u49
1Lwu79ZEy+2lFh6lAa9j3UU4Iz+AnT2UKF0GkvuS/cxLqCJ1xP35kTEnDcxz3nkZ
YNDLegCI92O+1rZyG6kBfX+6UfGiw6Wt4CWHHcZpLTP5EXL048IBpgU3i0OxS1BX
5RUw3aUo3N/9rtl1nMWAMvXGFaQNWXeT6uQXjFh46s1GsRhPidRcC+y8g4fffTMI
QKF4MqqS4ZeEpe2vLML8juZVrTHrgtFQj2LhNjBSdkWH9ET832Y2jY7LRg1L3oVT
14FXT+0IdyeMJ6zl9lIduQ1yVQ9WmCQ32Wz9qOCGo0cwNibMwDygx50xaA1GNbUN
DR8sAzLWjvrnpCKHtVr6qu5SVYE4QgFKqco6B61+AL4HNNXagvIUw94DEUM2SZMV
THHXqXCetb9OKjyNktCqEICTOX+34Weg9EPBIOHlhxDDWR+8pMI0QPFVJyaOU1a9
Zc6aw8YT13Rq/Ozhy3Q4wKXiZAtw7vpTU8rlqmPuWFsrb+4pNpAEIQPqyufkCaup
6ZEJse2wsGjuMwagIaF8P4ecb2IHWaSaDNsRYj9Vsahbh0eto54pqyAD2Jm1QIIK
tvW4oFKthx84RN/SpQqEboTf/AZ4Q3wR1io4hfqKiTvM6e7+pk3ixJzzuQm/7f3c
J15Ab67igi2ydRRIqkaVZyQxxLMsdxBLb2YwTCzo8H6w0LY0vyxxMAGahfapYMDn
HazL5hp7SRPG2X3QrM4JEqzudZ45kUcVn7SXQxZgbEa7V8igqUviOo0kGvg2TOpY
IGK1YRSeqIFwF6uWeBv7yB1UAcpUpPH4HrUwbgSCA2kLZgK9BcCBvOE0wvV4ISXs
MqQVPPCfqf+Wjp2uatFx3VXP7q76xLWoJBwfQY9t8KVFQA8TVzdO/GhOGFcDHa1m
V+UDZ1CwUz1VRPGXRRgtXvJvaf43lXgqhjj+pn/zJ+d6XDx0H2Y3DH/LHjRpWGKL
SSyONKEUpIJ2zSG0VoIe4yMTjl1+wHbIB7JMS1y4Jh8XZXS68zessjIQU9pnqwz1
5yNA15UIxN58GMwfiObhq4+TsPEGgR5BamQBD+f705V/QUbasXmXuOoy2arCUBtF
qjweePzdo1BmWEQ/HuZ/KoNjRYlq6k8tTGurRvOOCLmG6PoHBkxn0P18VyLl7CVO
NGGsi1kDm4IPoQ3YQZa8bW07w/geVPex7HsZKuwnSL+BL2bONAWuZxdvT/vTST5Q
xZ/QA6YifCkVfPN9wLLvhKZxhPazci1Kj1NViGWpE8RO4vMlDyPu8pZh0saCp7oO
O3AFKLX41hw9QDbrIkkgDPsAeloAbeD/j+QG6A5Yx2keV9pwESXaxrwTEKF2F0gH
w0bbKsUc5nosuTOLbmvwDIlzQHzIjAUz8X+ZaG9irw/iPj7s4gjZslfqj7JLae6P
DNNGKMiRZn/ZjVz2mfARq2OquTcW5LJPFJ7ZeBpOrzgnvr5yWFKrDq04DZu5foLy
A0bcTEZViWfEg8midN1BZdkS2Sz+58vYfOXleerXoPibF3L482MGtgR9dzJyuzKm
Ak5QOMMjXtDlIRZdBKb6QzW3Vahc3M9j6lzRAo04EyqN6X4mPgdG4vPEg0XSub18
fV1UkW5BanCgzVeAIsDBjYEgQ474RGldTlAt5pCU9N1vraZwwOlv11cDl9D03A3Y
GIwSYg8w+rd4A808+gmVUhn1rUjteuz8t/c9Kv2j7w3ZWnjOum1o2LKwFPVEo3to
H/O2z8PB80LvMlgv+UMm7xkFKAsuibgsiJtav/GD/4coKn2Dd7M9bgM7IK6+yzNK
/9BX4pMLXxCJNG9YYKrBpPq4t38mLE8VFjsFOXJ7W28OSNJrr56A9iT7efsx/xvL
J88ChX5MBxdqM7MhrgMG3lH07x48SrQokJnaAlSCYJ2TAmYazjsEzQX/TGhgJNlZ
Dtno1Wo/y75LCrzWUXUJ6lwg4nukI4suohQv3+ESC0ZhN5ibdhCIMF19xb+zoi1l
NIy1wMXAX3uss5bLWphAY+Wfq21VTDx0CNrGhDQAFapYDSGz/7DUcQgHv+EitIWt
lYjYJkwaylQ1ilGPCdt4KW5FX19NXnqX1NSKU1vZtFmgsTy3JJl53/BdQnI+QFdF
wBKVxsuCpO9eq490NyYepE2rhJ/QP+anQ/rY/J46hOkjaMNUGxge5aTzJZL/f8Q+
p0FYi1PsMCK/qT9qzNKPRXnwW9+d0BNuh5MQI9ZwA89z3FdIxMVweTBGdA5JvyIN
qtaIuWgsIu9FLEgZa3z8h5gyZD+4Bp3doKV4+DnjuYOJG+d3D8anN90Gg21oC/19
B1wxC5Lr0IeQeGPDYaWmAm02J+dEmA3TbnXQgLdUtnXYKd6aDCzJkxsKkPQo1aya
fWRzF589PuIyhmDBuKEcmffqT+mrmXix/kohWy2FmrHeunRx0nZCtIIsI/rmfUlc
F0htOkXqJURAkcdmO1j3osJxhVbmi7f3yVpdsh6bMmrfwOjMCAPDjKBwHx+OiOgd
+06GEYRv/kzxO7OATiQX5L/GWC0mN0YYYowQW6Yo3CO3IExJjlrQbgIFUEjACq8Z
stMwwI/8vkk7eTtOvdu7rsdW3cZf12ljnH631yeORWJ9SfMqEoJFxeC0BQu+jANN
fLyKUJfN8ZrtA+oYJQ4BLN+jkHQhV9oCHyluH3IXN35XXZ3ChlUPqvD2B9d/pOEW
LbtaECTKtwHZFxxzqKpYjwXKDuaPyIf2459+Mmh2B2CHIlIk7oiAoIhP7tnOmGis
v4El66sdyEr5K4M1uQEVA0AS5I6kqzO9u9Uhi9IC0Au1nQ2i04UIXq5L+RouFcgp
zH7YTMdJyrIwCN8cgECyE4Qb7bdtnZ0Q9FqQCWPmc50PYMHiyOj9RTrl90Ekysi7
oZjafXmDscFAjYBYAtgtnQoLDsWKQsLrhd3KKmAn2+0Dr2FOyoghH3DXyW6pWeih
M5Ta+bNd5rS3IY5wyqDbOSDH72B4lj3eRZJpK+ynjLy7Vpcj1Zfet4KrShmzx1Hm
RC3Rl3V1M1nrQiJepvKFTDx7QBOwEgXb3uefqz11bdxzQVie+20uHLctLvxa/+en
rK33cfQI96/OA55MXPG6Fv5Pvj3Eo/syFCRt82co1gJqdgAJoq8cyt1oaC+KqROA
6gfuQeWKNG78LHb5p6BaZwh8Ipzq9BLd9SGFXxPNXPIJsHVkHbjGJetqLWYeh4y9
uosgAWATAWKNbJc/iQdlVccRiUSzZcYnF3fWPc4r8ZAaiDgFc+WKlJD/sPH6/xZF
lQ9Ebar0m6Iv1o0MI6oLaEKOr1c219svIkykk9rzSRHNyPv+TmOhZXzQ5MgDkdVP
yR+ZmnK7oKtQKiPx2gy+jzI/IiKn7AE8a+4yi3r5smm1qLQW57cm3Wfr1uWe8SG7
biiD6cjamymMop/BcyExVY0PeXQUkiVk0rM06Z4voqQBKFOBuPwn1uiCr8o6o/eR
jHvUjgH9HhR9ehztLYF/Mhhd4jwzkZVe84h+397Oqug1Sjbac0PhU4pDgtJdBQAc
2RbqghggM3Ed4HpMa9Kr1VtTf4PP9Je+AxEKgLn0kv/wZq0VAwxTGQAbQe2j1iWC
g7Qtt2GO2UNjsdzt7yXeNEl0LK0nmn7JIOu+cPxRFm6R7Y1rJGzjJ4mi1GZFd1dB
2+Ny8hOoEaJo8Dv92ZTkEzpcrxTqPN8IhjLvprlrffWrT8A1PqWUIZ/88TFYDcG7
ZCWghnjY3hHy8+boLRZQW3TW6+BahP7WHbtuoyvOc6UnvGqFlBDhmOWKv3/iPn7c
IOGO7DAbgdn3KWGUyext2ukra6nHqyTxTxvwtQUsP91PTe1MEvM8iwU8JO5Y/dSD
ORpvL3G6KnTIWKbzZu7yIdWdln0TT5iarCplcu+6T6Qy4x+SIaR7yqPHCtJ7graM
GAhEFzFJNEQOGQv5kGULas/c8osPARjuhq7yZAugduO12ZLgVvdnMP4XXCFT/60x
6P7DPe4NRKEqxID2/IAk0c1+N4Db4Mj3kWSpCLUGj3VXK1MeJkQ9tn+wmHm5XF4I
TEMNI+wIvoKIF3m5SF20N9AMPk5UNEgfVVM9vwsJq/hJZdYOht1oy6I3dbqi2sZJ
yIn0MVcHM88ShSc2O24UaTpTTgYSVPy14w3l/FsCLS2z9Ix9+Gj/09YwEq16uVBb
a9c+C7PR/T4JuXAObgW3SDZysodURIEjdmfDKyYVE5TNf20E8Xu5YlV/ZM/iT7df
k9tab+qlJKI32TrYk+5L3QvJA+YNLtvVZwZIG1I60u1Q2fROHG+XYiGmGA8uBwfk
m70TxtIfexbeOTmA7QEfMjJNjEi6RR2K62NLthiVVwCRKNE57rwiEhqXJ2JAhPM7
KrLwMnClx9cZTAHuh5W18yFDVjdnSMpBOLZrNh8ofb6RYfGM4Z7KLtPOZZXz37TY
ke2dNc55yLDROKTskS71L2epifoabYWooxkmniTyUCqzXAnD2Nl9a0pr8HgLjKv2
JM0ESFKkqrTH+1sIDNsZFqUSdMNiiyJvzI0fjX1ezd4OlqRGAlplgA0b9xKbVcWA
ax2cFurTjaolTiuazrDQiWI1hEy1FFSVq5EEVUWHvWoyub+IiW+ndfaRZQv56YGB
8T2cQLjJomimI1KwnX5bOAV9GWnt8Lb2zIcwzUrOybWtK4i6UH1DH9BVlFTmhLKK
vT1b5nt/EXjtxKEM1GFv3ELZHQ1mi2G2kiSHgIDbI8BvNs6cl0u2DlLS5AzvFtKL
Ts6nRI1/n12iUmx49b66b8OrEhRKVV5/DQdi110mBV8PaSrcQUEozRE25vzGB1IF
ql+VRNQUqyw4jg4637pFkNjPtuffvAxHKBsrxUUVxesChfF+PziqS/Yghgwhfssx
KiFRWzWZdDEI0TMrN4ZDZIR91ipMRoXOQujAQ5aBuwm2H+iuuKsVBsXGCJGcYYcx
msdmI6sGhgePJUzafjTmDqqe1kSU5rz8Vgzn9gQPigp7BUj2mbCRY5XyRavifLr3
osz6bPXCYklDPlV4fETRx57bGrpLxQV4B7rK3Wn5HV80/+rtwpKSuhuuCZwjF9Ez
TwTZ+78TOsdRn/HL0rSON695jWCb6jyMuV/R+WFVHfp93adJJrRcGy/hePhczINx
RouDG/rz1QhQrV4FOjrgfkzjayUgnjNIWw9r1ngdrWm1xwl/4Bi1ew91Vk2M4PLh
5steD4kM5FLhH8fJD/2NdSgyiuKsFGOAnrIDnEeiSoDdCiG4ENw1vcynPsVaQ9CY
kBSyTcBZuSQjQZP4K33WxBJk5djzMgmDC/zOWKACU0Mal4eUta7zcQm6k0bd68oM
nTImtk4tA1BCSqHmzxtWhdmSRTn3Jjs0ap5Lvp94TVk+czAB/Sr3g7wEJDNjstj/
1Qc32L91+BfTvrYnYaZgIa10vXa7B+sovrv/dispAkhs5ijHZ1GlinZmuQnxr+/c
4g/PNr97UEYC59soXzEe2jHyoE7r7w0Ly4iWNYbA4CuhUkC07HUSpKug0SJw2ych
kZbHEjyxmZ/6q7PDrgLMCmXr/TACLwYxm5QKh2kz3dDyEr3HaX+GoQcNzozbG4au
19yrUKiWO3zXyQITCyCOJyZqnrio+cfZFgM5wx+iCMp1n/B52iDOwj6bU7ckCirY
ltyY1LVNgyusLft3WMfBCfS+328l5hC4MTP15aZy+83qpXzPi1g7Hos0n5pl1Nmd
wdLdjtnvt0EVOMft2xIMos68sLPYdIkqzCvHwKSy/q0CmDUOdYvE8iyUVWXBK8WY
SPixl3HKQaxLP9FcufGesaKLo1sZLs4WPIiNbLrydjB1YIN5dA+LglkryBtUTlPH
/alN9J8CU+z/SEBtgoICGxbbA9jxfaqP0zfqbMGEvA3VQvb9grNv78TSNH6Eetp5
+bNdr2/oVgGLCf/nedUnYykOlB2oRloR4BmUpzJa1vzF7WzlE13Os67H/BejJIG1
Cgnx1iLSiH7xjHZfkBZaFYltEq1LiqQmjw2dFxOAbLfoM1OaUCUG2jcdK7yQIuEB
Jdyz9eFF60qzF6jL2t3IEEy2pNww1qWrx+/ZSN56LQKAAX00xrFGWHe3YcZNdGr5
Z0Daig1j2BqAUXsWW1Epc+r/1jAwQv1nr2LZTm2m8jN4GC+jZ6IzZfpT7Ho+Mkf/
Q45TGi7l7il6qTrBhFYF3g8hjtK0qu8QY8WHm6dMaYYNc2e0qgTlS5ncFkLYU+qv
9lc0CgsV1yXAwYFE/0h0c52Av6r11+i/ZJnca8Z6xw6MIDVe8KbNVBxgWD6sBCt0
byEOz6y1EStOMpsoRLQpSe/7pO8wGjm/n77rtofHaK9dTwZ09bLFxcXJ4uB40+Qj
b6eWQ+di0MTG7lwGN3bAx6irf60FEvUUT/HLgEbWlRzrIrbflESGnoq49JTJ4Pux
1oEjMPDr15ltuC8Bnt121fs+qJyLaN5/46+GfCFm57ocWFqVQF387I7zO4uqVPb/
kZvSbi2zjTckKbOCkQNfuCXvrK2sgS/yoyqCm62blgQwR1kunJl5N+KUbYbG52S2
1bI7yaKD1UDWzXGveNxbTr3o5Qa6QSQG2kwO2r9SNnhLVsmZV3ic57p4UgI35bz7
6312l5ueUHNOx7bjbTRLY+i8iyj3FjNAmdmzskaS4i4Q+x4J2+1dGa3gehV1PGFS
wA2z+jwzrg3vfLqEXCbgm/ddD7aSWrmFqVzb2/XiCmxoBOV8VFD0tDeXZmFtVK5v
SoTxi4HWATMDRp1D1vbTBwz/eiTksXNPpPMOBoc7s79watxefoHFMhr71mFuCEtn
Nj3qi76kdJPl5wE9O4tj9eE276mozP3gZYIaW4aJxZ8pC6q8V8o2BvR4EExsirLB
m+Ee1KqAdXLc/euvO+68CSAx3aPW/FgOfnExMo582uUn6srnM8RJVUXScuyPxsUR
vqg5S+eIA4SCRs44OREUYQ46to4V8NDywTdQqzDGrCN9G/Zp+v9NMiQbYkI9iLka
YPRIWdK0gFH7jLJFl1yj2b/fisth4QMlKa+2G4UHfpS645p1yxUwxuR3cCA9netu
Ff2CsrmzpXOu+FFUhlDJJLLwDiVKbnrICycOTReKtzqtWyQO5F4BZoiCWfEbRacW
DC2PauGa41NgAIj9FTjHtOlyd6a7TplLNt2PLmsplvuSR1XzBEu7EYmKSzFKCTs8
Qsv0Sm2LPeXyZhJ0iwI8DjTzwNpjQ93hSd4vftfT7kT75nfE27QeVClBTzcp5NsF
3cZ3JP5s22MFOnlS9l1Rk/5wlc0Ws7sENO/TUgSHPSsjN4/VMK3ipTas46ACb+w5
u2620vUwmTJSYQNGHUJ9IcVE45XRKoXIARKvlGI1++KMUiVH2e7lVTaEmhbP65Ts
IdddfUelkk5wTSO0/39B/aU7/YbBBqY73dE4rNqYKN5wAAY/DE4aGH21GxSPuBJq
yqA0RumP+9OkPEXkRRRv19k5Rpe3lcfzsjZAMeW/skw2m+iiVzurvDDJEpZrCQu5
4mQuitzQcrtPPEBEAuzgTlwVrrpH6KrkxCUhW2/FfRpVjT0IA8NiHByn9aQSATlQ
fQwG8EbkyjnM63D03oRm1IvWCEt07wQjl6pyDruQ6hjRgfqI4nshZntVzmH0qkO4
G19YsLptVcXZcNccI3RQFC4JlZqUTI9HxoRMePE1i6qQ2xweh/CarcoJT2B3wSaN
mCI+EXHxoCkLY3uNda3M6mq9cIIkO5MPI+Ay/Ns548O4OH1wc7Xk3LjaOZNcujpT
Q4hbXsZROSb6vzoG0V1gRwkWutnaldCtaUqQ4BsipKPIqJkLEl4RJXEDFkkKXal1
flDtYrQacc64rr+/gDGr8M5qaH/YEorcDxq9QTNfrxyAE1BNbZPxeKcYo2EEHHLw
t9gZ/RcC8RKyV8EQLiORl7OjuQi2zHXiIFzWfUjtXYmBaizQZ2Jytau7iJ0KipX/
OhFVEGRzaK6OOguHUIrz/RruJXXzTY0hiev9Ba6IvdZGlDG4ShlyJ+cxbIThQIuT
SmrV9POUFLSkaRabBaAfkN+nq+1SDeO83KULMJuH5L4tnR7Vv6FemCJJYLlhXiez
UgrGnAPoPJOz00YRjqUAALHEhuAfnNJ01mPxTccTjWCKRaOuN0F8AsX1Ga/8RcSp
Qdykos23I1OITT9X5HHCT0MPgVBXZm6N3yrshKNJxqBMbDdps8dhUku0UxL9dTZy
iB5sBw3pOTmqm9RNS6+M90W7Gy6IqqD4vN2/lfSUrkjG1QxDVCi0+ikw6HFIOWbI
swzFx73ghKmRWeVx1fx0f8jIbYRI3Xikx/Xp0KlwzyUK9/HraCV9hAoobVPgmoMm
SqrSJSHYsos6GctYEEIpeLAssuCmEDGgL9V0ZeKO2xoTkmQtpaFNwR84ctfdcgqR
GOY6wJ0XnU0SOoXsKQvvYxS6wGo+JiMAM1rc9PGuqbT0yZqfH1PAcsaREYBhHbaV
TP15UFaWGHKlAYgTP4c/JcIwKEnFC3Kz3ZoWuRWybHiMcBWJrpCgvi/w+GQ9NQqd
nWKmU2ALa/w1aVM5EwWpqs7xuj3GsmYm9x8836XpMzgp3HIQ4GSRRpxCuuiijbSG
0DA5h2nQjoUPX5Upononged3Au5gMabmh4TABD0aIRdxifD5++RKTO32hUtBGxSU
uJdsWoX0fVFIjxNElg/Shprap9MLLQFwztUbWaDqBX5G0D9T+p950EapipnpgFAz
B5oVp7ZPWCmGvq0yd4DEoVLc6+gIdP8nkVHgmrc84JpgF1Len6Af6Ubc5zvWSiDW
lry0VZUJindV1HyUN/KK3m0IfmdWTXootm/9HN2aq66VYG4rFIw66hF8e0qKwdTL
1gAw50dCFvz2joF0MJL7gMCbxPSwtFLzRI8PqwdupQdKO9fY4w+NGh2Qtcyi1Oe1
jBdFC+MLiiU9pMZ6hVm9urDQy80faItFkv2yOh6a+OjpcD+MQ/8Z/9J5GpJjh+qF
sjzxR7j0shijp8Hjb+MSn3VPE/+In07FC/86Wg4bPS16T72GATI0DxUHI/v73ccO
J1oyp0QTLEXSI4/ZG+GIo7H+ZOlOSO2t8IznQhCNVpBOShaY1hhP3dDxu2CDTkbP
LG9QTq76r2DAvNbe0/pA/ayjn3PH1UxCwh6HrUQaYFZLViBcI7bY17zk397262NM
7+jB2uJqOAXQs5ZVLrH8r97aFCySjnGihEnihGb5gnbUG4RpstRzC9Rn5uMEtymJ
XCoNNWHrCXqXtFoFjKiNc4fBjMrVxbRgXuQeHSoy1gzzYFm76HMXd7WwbzU5ns1O
mQqjRB4xSYl+WVFFvkmqCbBgKOPqZT4wCgj1rCU+7/5H+YgoaaG+sdqtn0iyy0dN
OnTpnlPq/nmQr7fpO0Q+PV5LaE21zPMoIo+4a2aR9J0RQ7+v1xy2sEmK1vaUx2iT
ynAxu/618UQNzoF1p079deb438m+Y932ZhJHtRoBHxTf8DyxAwIPyfd2xq0a2Zfb
qX17F/qGHwj6CZyDGm7rLR7r9L+SOzU5RcaWkY+GOjYjliuxV7ymt+W2yRMQS9rN
9wl8MQncE74zpaArk3nlWfF2Jj4jLftNVVfohbyq+8yv9ynw7T2Jaeo5ksEMZFzJ
qcBIjvCLs7QU+gciOzivBtJcvML1pHFtTSWNHIfS6OF8wchKFJcJitZJS8u16M6B
/yxfFJV8I39gtGcJngS76cKY5bGPRpuYW4CbBIqTEEmILtrMFp/5rtZj9ImCDg81
nCqBO0mgg3cdNbzMs+ozb01CwEJJRcak2WOI2aZyp+f13LwXqDU/miMai7Js4ann
qJxz63BIEiFu3ft4uHD9C9FRq/7y7UaUT/uWmA/rVxsnNjzFaUdk1RE8tX+wX0PY
DL1n1ag6yGaBm45LCAmqALYl4S1BUznVdqTDXulnG9GuVOI8nw+Zlm3/+BW5oWRC
r4EMlkVXLIHlKvVVFXorVZfUUglwLqU1Kd9gXi62ihqdzqrV3AYYZOcR2Q7HZcne
AW9LRzhrUa5lCtc4okQIUmnip2cXPko0XkVL/wmOPxBG8sgac2yWljiusWqYcY2d
5GmMl6RJFLyFslW5MgUCCwzW1BXTnzDOe0aGze7KzLKCoEnYSE4da+EBJudhlTc/
uXFdzqXsk2MDdviUWmOYIlHdNym+4FX4NOG6R4roQfxv2VZ0TKThlHWy8GFM5JuJ
EU9v22f8xuWyXzLA6fiod/CvXlEQIMd9KQoG2h6oYGPTu09kt/pNCb5IBexD/GBD
5xUjVixSd7bD+gE/FftHIofe0viJvQHyD6uyMABbdsYbo64js+RRSuBomKctehRF
4fpatvE+0/DQx6yE3YuTrMJYnen5dRd9Cf0rkP/srXch0TXVBqYvfQe+uJX/SogE
jJoLsxWEd+wld6nLueKVEZP50A9jT0c8FZGfZcjTlPspr+QP2qvZ+o3oHaWEwJ+X
BpnTHiya6Rz+4HW/+cm6sTF9lhgY03I6IUze8RDzod+eDi5+nhL6ZiDVLLvzOVC+
zriN8uOfIKxJS4BpNMUO/Px1MCtc1Imx4kEte0e/6QDOpMk95FUuzn7P202Rt25a
lhrDPqmUH5cRklSGn/UKW1uoOT5et4+y9QEG+P/0TGWpv/WDgdXLPlOlPkaiakJJ
iK5HEh9oe86af3ekFpOkAAFSkcz7JDYxK+Tixe+6gKC6o+n2KrPyfFwYIYOSuDh7
UjiHe8rcLZ03JrDR92C/ar0iH2pvTRMZdG7rDGX2C5gx03Ac0uSYZNvWIu5hdmEE
ke6MssJpz/avDDHvd/PNhF5lvH16G/feFUkHNI9eqUb/Tr+Nd4YuxwEC9LKtMIH7
8j6OM+zwMaO3iAanycZbM9jRB0A9mti4fP4UbvTOMRQ3Ez5E0sEW0lN4mbTKYDfw
/BTf7FAvARTu61M5gwiH1l1Cq8SYrc2N7uvbLj7SOCf4dMwXmQ6zTkgMbrsl4h9z
lmDZnFFkWF0d027O7aFoqddaEYTZNWc+WOX73OhARQYuMJP1qUvqB9VeC4rk4gxK
BNWjlaqlJYgab3iMgMgUvM1c8JSJO8z9Uq/FbLq5xsq4fOMQ/RDFCtfETJRSpZGV
AMLpzj++oeIAWqN4/wJYhuB6rwIsOOjjI3La3czOL0iVizqXFZrTsDg8O3pwQDNp
+hoJM8WZ8JA1FJp3Xr7nfdajFok/w08Rm/Qma+wNzYOu6epwOTibvyJfU/+MGxk5
nmE28Vnk0s7Z6K98u9gGgxHL1baCOMiwd8y8CSjn90Vueie49rxrLO2SXwYL6I64
CcuLCU2B2Mwyrmh1nuOmna+kt5gbYzkTmARbHJih0X83Gu5EV9gdosYx+CogbXFR
bp/rCRb5oZ4em4XLT0EEOn1x7DVG7RwMhbaZxI6YNFQzvU235cQbgK2UHhHaFdiQ
lmYDQuEPmabw1d7Q1UDUm1LEbjuhOY5f4+dpe83gMCeO3ofY04aJxrWOLWlS5NHS
6f5x8vwnMheDpYPGbtdx5DbIVoD1z6Ik0Le8zlS1jjXZgYUGur/qSYrRRhRDkPvu
NjnbFvItPSiCEghApIromLTqqoNe9fFw+juS6vGuzxkJzP+WJLOV3Rb3fBKH3AwE
+uTIvScGXmCgSiLH4xQ9x2fgFxmgOPhhMrkjEcKq7/Bt/Hnv7QGazhHbzMIiZ8/U
hy2OMiBQtnXK+Ozfk7tEaEJidtSL2ZAae+sWBX7VqW2sdkVkNgf5PagiS7ZOo0cG
rQyDdxtKfe0/n2+Woswc1dyPAHsvkqk+xXDhIfoiZpTXuKWXQlRD8jChV+NYBrqY
Lzl/WqQ8WjZPgr5LQzl0Do3aT61ENyXuv8LfEF3ZbnYJhoglM1vGyGRw0fLVDf7S
0j7S9mhNHiIzuCLSAhm0kgbs7uK3cc5lJ6R/6ZfXH1SlegXCFTk0jYTDSeOgg0Rg
mv/pPiX/HiuH8etddZh34aQ/0e49Jqq0s22VEfuh5WlwX4rpOthrvmcRlJnHh33q
5DPQ//Rna4zH/gq2PtA0exBx1aGYPsyuCAjP+TECBkfTkSk4yI0UI2l1uc3njvtJ
XhDbDk9grJPLW3cQpcEnWSw1fk7ST9KWiP4ru8QgArmxOlEk4kNMhKaVbKmbH8Ri
WYiXqt/ypYKOPbuXYsWkMlqHQ5JR9Z+jZ40pXxCz89MhaP/LIWkwZwwVTSHv5LZx
59V4YTslTVPuRvfcCNPRqAkKJJYHxLAszMRwsMLbXHHz0w4JVCBxCL34efLmLO+o
FAQ4y997j7j4zkcTDb4y6ViYlnjRBd6sf+1jxmJfnA2eDvL/ZHbGoLLIp8qKb8Pq
W0v1V50uyv353W5DeQUQdXeH2QTY98LUQ3KqJWfEp+ZjfWTP8slkrXK4zhwLs3f8
pPxmcqnkM693uOfEauhTXXHK5jPbrUsy+g0MtRefNfJ+wPIBpBhuyuRnWQhUPcEP
TVx4youh5TqA4lBGxegUJnH/XomPfJ0rTwtPE+yLtqqWDvdbcKdyodArBzIvIVoL
CnbxcGukZ00fBxcMCq4b0IO+9+4SFbtc4H1f+/6z7tGpnbflr1yOQoQKEz0vvCeT
mbaxU2mqY/L44DyeAtaRXIPdbHjmGP0HVxltVDZ/u2CHmq/VuAlBQG5EVe71jt94
hN8HZYlVB49fbN68y0bF/PlGfN/tEWhrCFO9JpjA742m3v5U3y5X4wEbdcmyHzKN
f8zRGnLntXlrpSo4JHgmk0pRZGqDYoKmZWmVlj+UUCBPzYEkAik+XZxz5/Y59XCK
c0d7P3u8GDnDbo3d77qJgBmXwl1Q2jmU/HWzP3HkHB7ufih0FOS7mYuGoUgvkxe8
vjfUji7gq+9H3DXYEarP5fcQmZZcdAGeiuFdAirukPqwx3KhKL/gmCxNZ4eHqfZ2
w/O9BT8hMEpLNtUtQWuIDLD+KctyCeQcWw6RktqOWk8rkbiDb8UDX/Gf97IGVJAt
UvBA2XTuSjUruhcpG0bBoEThcpge2MBjMAcQuGBg4ePcdTSYwsEzS+TCrbINVOU4
AJJsaTtgtLuHGBc7y6jz7B9b1BWGXVuW7c2fjC1LAtdeHhmGa6oepMkBDr4xYrmR
oXvsMx1bwbhrovq38AHWK2lxB3uA7JvQLW1KAWHADrKUZ39xzKTKZFw9hFMNpnnn
wIdDsrx70xNubP2KgSN6nHSekURfshlnFV2MQlzPoLmjLUCv16Gr/YZROxs3UBdh
6itHMq3BKQik/xo65iXcdJDpD6GtAlwz6pwUtzsIxEhPnLxsT1xQ2y9IoGUaNCvF
zwn55t0jG7aVkb2l3TzGf39fqj8E37uXbbGcUmIkhBOuinl9N4TPjhHwuwMnb4u8
IMlbN9+vXxz0+DsFgCqOIJeJirFU9zuE2OIKDZ6EZPlLlXXO/+ZXqbSOi6jzdm0U
s18X/KoyazyLOaJXpARM3ctYQ+KEiGZ7XkeqFNVsOx+ut4BP/zt2Dx67f8P2NDYB
QCEZu+/iyQgcXpzv/5wcxsoFWYJluYSFDb7beDz9jPsuCUH50WPhZva5qLUuyuep
X1lD+s/JskjZZitQ4dA0OxrbjAiELnk1nGOWL9LE6iKBRLSnvo+9Q5e3s0SwkW5R
GP6+452Y+jwfmWUZlmwpbVKa4P7jgGFq/kDdol9k1NPDCON3h5Oy9vQxqDs2mL1V
/w34fjIkVRIUYmfFLp2iDX/yKHxEvmYA+lxHkBZZQsXrRSamqiEjHfGqRlS2iHvi
vp2y2sKg7mOMygi+Dfq8uQNqX6MlX4JXqiug49IAx/oHBQmGJ6QPu67rEQ4vwFDq
LJYzOpkFZkGvzFFf6UHnrh79dJUR5cB4NvnpmtlBlvpAgu8huhd8p4WBHiA2yY0f
GF5OnSAZr07DP0xsaECGvvdzQvKZ72LYC15tLbqXAj3elNOktCkS+zi0qWJy8GJx
dNh+q6jCztHMouJdQCnsXopCfm53jXul/rMenfUsUuT7sFrgo4CquBfYFDcITHgN
9cIDfsn3K7Ht6r0NhnWDEw0UQYnAFYKdWfNrMJzTCvYd2x6f6m/9GCb27hQRYzG8
HGbzOmc8ezbtLF+bKisZyhhppM+MdFBEoLKvGEQuXz9/rMBi/cwGAeNfqBI2Z4Qg
/9gg2QZqHYsVMXcU7r7uiD6gjiC6Vw+Rmljmr0iXXav+MC8guubXT1FOvdKOOWIp
BtDmxNnJrdIufURtWjJa53TA3/d1LBrcfueCneEjYTGsk+FcC5v/33RnBMJWXC7f
Qmwv4ikUE8HhrWGWLBHh7uxUn4ZHRkeieWt1B6nbKY5wWGBSaoRXIar1p98SsXIz
P98PkLKfoqOpWBzahGqjw8VAdBNTM8wEnwrOCnyflrTWjVSq1YsF303Gmg3GDpwD
xwZG+/VcZeVOlK1lBAAB34wRnv+iAOJBfYFfs1rxYu3gOU0wgkdJShGihPB3lq4y
igNStxJ9w4FNJZOKziFoGXHSQd4JTueQI5fjE9TOUW5fioYU84oBkzuA9ST74cvI
OMZ8MmEaC604ifPZIiEWZUyTUv7+BmanBJLsThzYJp9cHcXVmT1oro3v6lttxUjk
FCIWWQdCxta9lZtfCQBxRTO52lTNMGEKB/Zm0FfERH6YmahnzyWpOkJE04r8dEoG
oyc2YFYZX52T+5viPirhsOcIaj6ag80/+6tuVgbwRiVZ4bkRCc9gSZfyU5BUyaq7
z+L++eJbgMO/hyDzock9pMttOeeJFTEKZMQSgZiMYgoxYgbO5G+8K+iWN3WMNG6A
jAkyPfBKa3EPpQMTh6orlOO7gyUR457YrkoHEwgEmqii0SRrGUzPaRHY/YxXQEeJ
2fuEVbaIWMXIPBeHDk3KsYdCl9xuXfmsPm7FXssovpvmCzJCWBdnoVgzk+gRVrtA
wmFnyuHbcRJ9mlOCmmtGwaVD/4FWaRU7ekYhRzVAvdC7oOLrE7VNepq0Rt6j8kDk
qbETBPIIjfqhTRat+8XGSGpHGWqikTTzzH5ZsRRzrGveUyIWta/L9rD6CLOLvgAv
VncoBuLKweYccZmiZc4mvDStX2NgpzcKpIPCUrz5wgLl9/HqGDABGfFvJn7bY9Wd
pWFFncukNg5wVOH6ma5Xi87opHsnTjP4VTlHlEaaNvtQgkssWwuyZ21bz0e356oS
HmqM/+HGNSyqeIKFAf2jKDtnsQnTMjBg30gPc8WiV3SvAI1GjuovkluuXWkhaxjx
QXfQTYMa+ITzaHe5nmXsB3L7BFgbEoB4bMYYtr2Yl91pQAYrEOftKDEdVlpZWiKB
JTWtp/aiXFaHVsLHbp2Ls28groMvPI7qsfd5QUroOGrRug8kZ50aVBaa15B7EQmy
WpWjt/iIEEW3Yq8xs7eUSywJfe11J/HqqhgydfyssX2fKLBO/PITyIUBY230aqpM
1pOM8F8xOHNaky+CzahUQEdwZHwu9OXmBrj98N+01Yd8kuIxGKnNmHAwf7HBaFS5
wxwai1s+Qk36m1+MFdTTfKKyACdT5lQV/73etji4Q8Aetg4gubw30rKnORWdXaPe
INxsVmiQQSRSODMvaDn6MkQH3g3gJv0F3j3UPKlSrSs1WMqLjN0qY3kXbxo6BCik
DofAT4BIECkrNCSKvM1WCEUtpGGV7KobYoN1cwV4apzkGORWGILo32arJh3hioRv
9ZOb9iAra5N9/kuE6ScrrGSOupM/yLkYgtG3Omap8Jza9Jvm1Jd+yO771zGKtY+X
eU5xcp7QHWOZOkSgvB11YiXGb7uFGABgNwsq+gnBqu74iwLBtcgwwR7ieBIanp7t
LjorbAvcaqiMV42GdAlDZBztsdTSrGy6oS0XSKYjeMqgpLf7OI4sO6rJV9y61QZk
IqygkWct31sAV7Zg5JYFT31s97v83m6iD02sGEFxWIXFxFbZjaMKH9vCn1WTncY6
eJ1azC8MOdGu+kcBnBjmEgnW8zkY2LNsQAnmthFYPsfadJQx45LxeuU9s9f3UGIX
lHxm33pqAtMIwyAm3QvlKMPCEEnyQqPS2kC81kic3hjfKiAjTr1sDtwg15G/soLR
XNPGSygu63GVLdAYfC2rrcfzxLLAEmPCek/ihLFalUkRLOphwN8pyjQspaKxoMB2
kFAqmI15vq4iFAkq6FUNdc433zQKGlisgLpzakGdBwltsZeyjnB1UOlzT8dLJ1o4
nHpZpgMWD8kyVANbyqkF1ow+m4hObuVH9lbx86Hs08l+qtEMwG9WqT12MTwWSCaC
wwPgWBSeaL7SmsScFuWB/IoF3BE3QYgNohbvTmQbBbGjbYavEajbQIEJF41qDZMc
hiaDKVzN8Y2QCjykmEQSfYzVwQDNBV6+zxxQ/wAKY0cnbz6x0yaLF2UtxGT4tuUo
jxCfsl87pjYBTcdYqeeQWGCaGPh2taC8FDkhz8+rsV5Z7yiNwLhk9BwWZg03tc62
WfL8T3DEJr+WWuGvFFckDmCW8QEgSeT+vT7naotNydjSO7LNhJYiXVT7aQlSj2zr
oCgEyT2/V5EvFQSp2LUg80NmYc/oPa9gyzpV7cbQMxRJV7Tx+jwCmA2ZP17UrRj3
TCsW/bF20VWZXqqjKu3kht6HPgZxi+2f9vDz5iKuBOz48S2GPG4AkzomWBfERywQ
xX45qOu0WX4A9FuKRtbg8rEiWAvAFo4GXWBB/6hX0owCqVXVm2R8mPIzy9V6tlwf
G4NXybCEeYGB3gaU7OxDv9MH1H3YCZy9bL8rn1TD5ZQeuS7M32T3J6Riy72kMT10
9OeWlmWws1evGQFakiy1EEv2iEboeinNjwwuYgVjB48IVQchMRO+a7ag0ACqQ+fk
bypyOOlBg+O3Hu/ASUDHwMTDhAF+9nhEmkUxE5JLGQTCI7RgQXgT1b/GlqZ1AXuI
8xaK2BCLpfWREXRSfl+LG2NJ8w7ZmTn9yDIu0TNlYBgozgJ1jkWUXhTXUBdxLy1k
9Y6h1P4CHvN8vNiKaJeFAuzivG0DtnkJovcojmWovkLnhrFTlYS3KVac8t8MxnKy
4EQQ8m+vBfRHlJjSoh+XxeX2i3kVx6HuOW98/mLvJc5Rv0WZJn38by++kNzT9pVB
HhdXuVTjRsGgMkn6/VVm/qqmjuhqJ2fEjL3zbESjwbP8dmuSCkDHgCzg80GnqmfA
HeD9/pvNso0ZuNIYTta18Eko1UZ2MoyKahEX05v/7hw1AUOzJ9tYKr6D+esDVJzs
wuwa0BGMAuknrX4pEK0PLVl8uFR2vRp+LOuYx52y6enoWQK34N9JzmG9njrIcsBv
vBsSF1gg7SYvgWe8q2BSH5fRwsiMmOUptEFwPpvjcLcgf0crSMCV2jo3q0L8oYy3
DuYqA29gAdWuXCCv+oXVnNzn0+5fQLqYH1pqfXQ7zZgS5Hbyu0+nsoMbuM0yLM2J
BCQuw424k9wH0wQ3hqcqFLD8zO+vJ1MI5SmEf9nJGWdgjohrRz71myFu6+maa859
OUwOIyhfUJIEWdc0S4fUhev+SL9uOInH46MSdYYxpLFbyXR4sl/33NFzbrHPIFjN
H0Zl06dEMGAcpa7DpyyXPlkTSOnuB8Yj5wAqqO1x5osRqDQzYXfhL44GHqrZUQ+C
v5JYUzwGp0GXuHnQXCWycLSvWoPxBl0l3Icywpq93SHAOLMjS8XxklQTlLsFSmeT
kyKy3zzN8O3dSQusOFYbtowYUWlbMeU9qNx+ycmMDK3P1XGSLSUXTRD+E+BR547T
cWv0MWA6LXIS+0osmBDgh+nX32YCNwjQFHCB9OXV1bGhF+RPiKm5QfhPuTz1U0I1
EBRAadrnwmdqx1mTv8p99zdY+ujdWn+lNrw76NM0Kvb0F0EBN2etQqnA7fi/MrFa
1czLRy1UhXHvRugISQT+ROkwC/GjYUrr3COAMuu0GNRRFHuTFQNcZBQPimN7NLTd
z5vsdaLbI8KUafKp3Ss8+AOc6z/S/Siu3Ck6Xr5JRdgSmdT3gRNMCCBr1qerlbMv
YS1OhbFlCFZy2li6A8uZD+LqY4KnUdnGj4o8GHq4r2f2ZmgRYPMjYhQCQvBl9upF
ODRxn72wWLJA9CsW8kySDJmHyNP4TqKFHP5XMkTchug/TSXx9Bbbdw7iKxfYlkSa
LBuZyYJZZx0Mc1Qv+FaOJph9huPgy9B8q3PGQNHRmAjH5mOZdu+vVoVtWZwakVuW
y3VMqLu/kRKoEvZEsh1IVR8fFetGLOIPJ2Cf67inDX4kZn8uPwWajCeUYj+qp3ow
OlTQmos6yOE212gXWp39LC9li+VPW7zZ3fYQ0xkq4Z3Ts/QLrf6Wvr7QhWtw2A07
2BnWQ7+ZEAvE1E4H9E/PtUkcQPtszeSyn8H12otg+tg54qSkdq7KuyQRYaGz9vJ4
BT0RDz0cZcTtMBGDu16LowjmD5/yGWW12+j00oAXuhPMi1yK6HC5O40A+WGhOfct
gBd1jbQv/YfOEPlDOgCQD3u92/Wk6Js5YuI3BhFCI2C7nCBH0pPVGBqqeRBxMRKU
+7714ySf/MHzDpSDKMkb/9kyonxsI7wyrfRH1MBoO86Oti9jdUfUOAP7GICWICyb
CXqoh1X+mHjnvA7kZO17PFDBSgTQNrRUy/njrjKKeJSgo4JGUFEedonzRswV18/o
F0TGEoVxIhQhG1DE1nU+u3uu74TFkwi81+ncBQ1Vworm5594fnoUV+2cTipH1l7L
U3ZEXgLUErrKL6PA/UsLwAqTrqD7PDpZEZy5S2xGFh9B4RTrMJ70436tz6VSHgJR
vFC17645q2BnuShYsFNArrDI5mfwyNei3wltoyctFWYoBBslmNCmsUEvdEmTPtpe
pm1FDTkaYbqksCt2U5/G0qAeyWRWdY6Jam6xa0xgTIQstnHt14lloh0mIWlOLarE
hLMdelvEqcCZZS4hSLFviIXdeHUB+jXYiXJGCKSDOZAY6A2sikxwwrGIXnmUnKp2
/cxpTDn44hRlVw4TuuPPi811vqlRAfInBcs/3HWxqDWPWJcTKQVRMipCSBinzL66
ho2ofaBm2JKc45YMAxjsrxuX7kofPPN8z6h0C+lx+iSrxUE0R+gw+Jv/zD8G/uxb
gA3BAQojdvZ570fyCQn8+gifhI/ZMVoQmGB1q/90ZL2E9qauNm2OKVFkUDwm1hS4
2rzRxVn9GDoNgzrEtSbcOPEW98DekRXQQ7i+j7+HS5taoPXWtBFkqd8WxQebS4OI
Vh3CmsUf4LX0kNkXYvrZ3x2G+ROONZhWDiU0vICSST4Lj5mrAOn7O0ei2qgFe3kq
58AB/dYodEUTFm6QIHvXL1WsB21LeIQCFkGw6cCqrzhleZQJ0kgzPknBiLuL2V/u
1sD5VU6tI7f3thIRrJkTBldNCkLnMMFhKLRI40GoguzHwYlz5cRnw3cw0NZlrva9
JSqt0DHUal2MAv83lZLJZAh3YfRAqJ68QZxTDW7PEzrvlJhKfWqTkgpTB4Pkl4tt
WXxtulhmyh0QxRsrR0caqS5R2I/pVHWdUSh7+BX0aYiJ0tcQ3uP8JwZvaEnpKEPN
Z4O92IhfvNVB71vo8F7m1zO/hRZyLMrDRKbUtOtjyLY738zXAXr9OiuWja0ODX3D
tQPEIlZ1PVhn+mCncLYwvG3tULYSHM/Bj+LS+nPWm6yzLMPgazVCXPYw8yOpWmXT
1tD07uDNNJG7oEJy/L9B81gMel2TMI7nXTuQR/2sOr3qcvpGohAh/g4f06uvha67
sZCn4vz1e5wWzPKP1hZUc7PzltH3aVGd4pxx4y5vpQ+9lyeLm8kHwj2JMbKwSKNC
ofugM1KEOIpFIavionIP4EJZj10EaCebHi5/5rzHmgXoNoxXg6JD/vJR7OxBbBV0
zcBJc1CfGc50J7g5nVH3L/mLuOjfBG8obEE0xOy9NWyvJT9wDUj2t/8U5QcIXq2L
snex6qQ2kEsO+c0cq3cKZYG5eHQ7GMqsfd2Z0i19N/v5YucN/tDK2CFNHGai77ov
I59iIl6QJZb2a91bvlzW/BmC3QvLYw4X0tScjRevOOgE9e5S+Xaw1DHAJDVP4Iph
DTl4PgFqZUBlhb+Cp+Oor7JVyvRdswhUdJtsUsnVRnvts7VpxpBq8u/RTGy1EdKZ
LYshN+Avl3zp1nN2QVXzJ0+0FtcVNfz+CEjZESUUOJ2PDfjipkGX6+abmNe+az0f
+GLOXi2M9k3m7/HaVGGfEGSUKrdp6YoL4G4aLjldvCBCcee1tzXOPOesSIXWLF8C
o4MD+aaZfkBHBO91nJrTWZl6Lo7QbFgglmq3hLcB+iWvBRo9fYxsZ4NdQ6qta00X
0W96ldh7ZSVxHYOlAHGGRdD80sSlfzXnuMtJILAvILp0w0wNxC3wzypFuAx79wkc
L2RxCMuekMGYRA+f/Jlu1wlurAxs+tFAap/DM98njIBNddJbPeaXkLFP+vzcZm11
AxbnXVqW2TMQ3TQXO8lbInrcpGryojhbzHKZ+98/9IfGbOyLI4OU09otDcnb8wIb
5hAUY6WBf7ge6iGpIDol4BxYeyfFeXg2N3//IADEuO/Av1mz5FaTjcVB36qEDrzP
LqUeePTCc6+eUS7Y55qW7pl5sblrAABIFOSPTtzzwtEak0abJoECujTrhBS9Vrg8
grhCTXdctw8DtOo5KcOFHBK7y3HZwXgZfR2mZAsW7gqS1MJZQlXrN9lURdFLAaVx
DATDy11kydZHXZ84Ok4J6vGamT3D5fqRTn8DBWHA4LGRM+EAiASsujIZ18lhw47M
F0ai72yAUZb7yp7d+HtRJ3scMye/rT4VELLtf+Mdb7k8sZ1eNFK7L2x5u/yam4PE
GHWWbYSdBsi1jVBsLWoyYHLskllZt0xtgsFb+qjT3xxJndol0gOlai+egTlFg65O
dmJfe6tKXTFnM6c4/psL1QcDP68JAKDyZTOyt/UyTDTG5653g3o+QmrdzWViat2B
R+39Hcg1EVTFC05Z1HhSCOAwxt5pCZIZ7Xg+MFXXWn6B8Ik8TtmOyOtrXSge10v1
Qd4OPSzT8vBQwjuB2HW9XwgybKLNFg/LBci5kndEGBkrh3leKldjRgAjXBtxPSJ3
RYl9v+ONUemEE/EISO2F3TVRa+0fPuvjLlyzV1PA33b37PdWmiYvXZKtn6+LQ0Hw
f9BesBnB0W/8DfVT5or0DuiQyRmDAs22DZBYJ56D6sXeOaSh6Owh36ad5zEue9xo
gT8L1XF9ngu0d+4JkT+yD2Igxn59WrH6XCd0uQ78SL6UM512a0mqd4Ztictai0Tu
IVl4Rjdl2dg2gg1JnkFQ+OcW3ciYBsNXHWp17i9NTh9I92hl4DMnBtAykKRsR0me
DQDsdfuH2KN1TeXlXEPi6zlCLj/+y0h1/owB3pd2ybUsz0FPdjF6ATtYArRgR94R
WYQBukvWl0KTI7rKZP1LBbeNvOuYu3RZW0erYHkMUjQI30oBEOuDtlbmxDCBQiy8
dc5bafVIfYH+lRkhXtBtqsN1MY2UOsxGTQh5crrTIoZf7N6J3qk8vBofcKbqP1cf
snDhf0eut+q2vU2pptaTnMIiu2vBcDtwTkFH6YHVCzqI5QdQH8jOXLJDwXLZ7gou
k9fFEvJ8jCkltoG9rt/RiTKTGy76Joy6/dDklonJt/DNi9g5Ys4oCtrDtZMCgDzF
hdL+7x33Gv9gSjJflSsff+O629xEkKsQVYSOJMH7F2FAEh6CMvs3pJfxoVqb7gIH
jIpFldS48bJ5Bj2d9ehInfZHZUJyDVE4xaEWdOlzwEL/dNMRGDkwtkmBb/r18S6A
v88JlO+y/AFPDG79piR9GJT96/l2IcN93MFLUsOOB+Hq+Xcon8FcKWWugKt5jt6t
c8tCSO7qvVamYJ3RB1KbaZ4ZvLnHkQ8H138McAGLUHJZbBf7cd9PIos9QpSY4x+M
RGrQKYydiiBQ1MTCdQ5FY1aE7S2tPy4dTAKVo4ihbCDiYmM0MGSJ4vqs4/5K4wHw
/G5H1gmJq+hY8YAzWKABv17Oyoh/wkUk16ENGKvdFOxWkwPJVVP382wWJ9zdefeF
zw0fD42i2/CnjDrn/DQ8TEfP1VUaRw4fxdD4xL28l+C39VghhTalklf+ZIEJxFDN
NrMjSgjGUajRolr1q6G4sp8WmvX3wVu9vlC/AEV+0KA2Ry20QlOhaQ/etRcCIQYf
jaKkFfq4efzjkZkP/Un8TPC3FYS1ymWqW61NUyOTLLTV2Do65Ta8rn3dN3pS+5HH
D1CqZm/7Lat7DSLHwFvKz/Z9GM5XsgXnNejHBZPsOiXIglOC4itZRQQNyQCZ+CM0
79JP1aw0QGGWGzHoVWzX96ijh7uXN0Tfl0VMElkqMPCpRfXL9o0jLje2BvIwOfsT
jvJUDqtTTsWh3bKkIFvfsT83yNLET0wTC/QEVhKU39p1VWQUPgUG/Cn8rnOmHXG9
Css3rc2GSmshsuuZL7N0FU2ft0hIunckybDkyxg2mnjuVyJNmJ0HgK/hml+PZTKy
EbGpbBzTypQt2pxr4aM5h2gLeSqNurIRWkMNog1UpOB37nn3BrBgjTY3egvV1uVA
Ia1peAr0P897vawOx3EXHePuiRZvVr2kgKC1uLpwZfgGwf+VH4DtGwuJ/V+KymDR
teEfFyyfi6HUSaSaDMo+5lq6WixammMl1ZG5o6pbTTsz4NcpeEjlT/k7lPeUAGWr
mnTQq0U2GvwGNQ7wuzYKE45JxznTGc7LpjvnF/BP/CtqSYAnLKwX4Ba9H8AxpmR1
dDx5WvQBxoM4Ob/RMcc3x5qxWUgERlNtRPeP1GWNpRKm7xSJoq0hWWFKAB+PA2Ii
LK/8Npvw8PyTtgz0O2+laFYlKnT6c04e/pbzxcs0UPygl/DCkBJs2VzLdyL5iVTK
Eg0PSKYCIzrEN5gNNYNoQrSw2ej5dcqBrj2ihVW/VUK+/+jRn2Zj++USbI1fOWGs
BZUC+LPf0wDgSSAAfjuSJbe0Aj4CvL3ot8ga6sTJ77C2x/xetg/NiyTD5EsU3DjS
H19SkK+Z3L8In4fLbEnVDDVI3x9S+AM9GAwcIESxZeZtswQnbQjIgZIWjGfjZT0A
5ejPe6M7VphnK/AlPpitosCWguC0N4t2I/qKN6ascItfIMT0r6VPFafuLWtNfnPP
tEuFaxYfBZf5sGruiSqDqfOcovEb3HbMCOe7F9VrczHSwP29UB1ymeEPDiv8Eyk0
kWUDU32jWCAd8V7hk8ylLpWZCEKgV4yh+nZB905VlmU863JNW9a8OZWZsaA95PfQ
zJyfQobiFUcOw217sv7ijTPxHe5/nAh7o1RNM5OITOwWQ+ln9jrQ8Cu0U1WBWbXz
85bgGcKuJQIGjMzSL0VuSWdhjcx7MiR5tbsgmjnMNJANWMQo9XDXyU8dYbHnjV9c
x5gzImZi/vXAMaR0nGrkuvFJTsK6R4wvIhIQ2vlR+e7cCYSl9LxhHcSpq//okDXT
WfurN4oBryWggdKPe1qADJorVlc5RC1AS8uBP6wcWYL1BnwA3uyEFBX7J4BKOZ/t
EYcY+9Cq7QmLkhHgHJkywHF6xvhO7T7wGAAi0fpynCEGj2El0dT1qbzYETNnKHqh
TSQ59TghdCmR42d0cvz+YGnzN2bIqiC665pOMlo4rMgIK7lnlSr/C+R9e3RqbjU+
iHfLR9MloezpgCGBOSlrZnPnWYgeKNmmql42VZf6gzb3dIIpmS55sje04YV2h4dE
sr6PDedAd6thv4LLAp/jqeEqDrTDkJJkt1ry5Vgu24qbN/OAlQcnjOozWtXTkhM7
gDTvQvg303PtJ+3TM8EiaPo7sChhzYm4kV7CQE/e6qcpsKLKABvB0JlQ10REozC+
3vh7UHahandL9qzzLtLRUt0LK2VfnnioxvjuyrRlM45aO3YN02hZ5gy5VC5Fqns8
28FzbOdH4PJEzgV7PBoQe8wRwgNxoULikBVURRTxrkt4mtmyl8Hb/GVKgkj6he57
H0uj4v7OqL0NzRsl3UDfstxBViOPrgh5KwFLGhNWe5nrtkLJ2tYDbi0GxGhRvPUD
ToXlL3DAYrb4SGiSbnAl5IUEJj6HKjGwPgqvI46qAg0vTXx5t3+JcUvy+wHYK1Oj
+WPUSki3EsUHpxHiPtbjswUMEr2Mr2QTkVzMFt7VeUbhQM8s1znRfJdOxp/QIi81
Gfme/2axyM/1hJOuWReKF1ct5UIOLUEdEsuTiu6OuNZw/nbWJCI9Yjmvm3yhuS7p
yrAHlcHYk5ExEQvTwnPDoAhaxCfcqpbB+M8Rj5LWQxwHwasPpqbJDC8uUahx0x0R
joLEP+oG6j2BOHvVxquBX2U60WdCPNv/4O1SXf9SSSlxaUCRh14vcrwCan20yFbl
d8/4vzYxM82Mgc5bMoCk6KA4Y+zZt+GD0CF4EtwYbMgXmzvgfCcavqgOMPJup6RC
rOQyx7I40de7lwSbNrquRJUszF0i1mJ97JiraipH2KZCxBF24ZkXMfjAh8OMXAcj
g7yYqyvWJcYsYLpuTDCbuOUcl3cuMT1SdARuU4/okmyY8Oo6dTrEhutJCKdDQe7J
ZiWMJzz8VyuPWtPCi7lOIC62HrDxQogwAL0s/ASmZOWTQtCoadfepddZYP9pGr57
s7GMHBq1Dre6u1Lufxoplt/dl9DqoWDuUfgsZ3LaDJrVldp9IT+yqNpK6emfTL8p
BIKRR4wLYLJYDcA1ehuOeZAiGQ629OkTdcuV80mgVm5zYBNnu6Kt2j3RVFllHSIT
Fhn0hWsmUuDR0QixV1uXAAh4wPkuuOuBWMc4wT+xcFyFgYXRLPqHiMA0gSNwzyQ4
5V/adnDbEFsKaIMRI9e9vbHMyN/i9IABsUAgE8eDavKoIaNJAUtatvSty5UEsh6q
aGPIGQGIy0tomgUmzD5CZzoEpsRxnVc0iLCy4UXUQoAij28ZeKjmzB2zTPd2wiBo
Z/h9BS/fZZKY1zJSgYnWZZwm3kLm3o9qC61wOY4RYHgS9zNv8WQza37jLDP6Hn5c
8seYI8gh+Ml95fx6ngcjccD0hyN2SevGufGe3wYASH7e7maIBuszN+sIL97XLXbR
xSNZvMbBCsWRZyiE9WcHVI3Ml9gp2783o1EndG/hvA+8j3AcTw5kRHXmx0XtS4zl
QhKvUr16pbRVVn/vU2geAD0ddsi4w3iwC8FwhHCQzfEIUwhEMon3VubLjq1a7gyy
QEO/NiDbwPzLo5/7NXEoGXZ8cd9kewF+CVwO/PTwjuG5MbDFja9+d11Y+gPOFNoT
gbDXKsodqEm3RH5XiuW27ZFUDxis7XXeJjtW9iBq5qpH8eC8zE3lwYx6ftbPbIXw
eM6QHZpd2MT/7YJhHVPg+lyJTMOpBA6OdvvBWF5Cv+gt83z5v+QLMr/cKqdiqFrj
eIPKoOTGnqT2QLOMhq+ZoJ60E6OiLjIucJSFxlqgcvPl30aK6JEQRawuL4XBSHxK
fK7mF5D4GyMSXImt0dcUjiUWVjvRoaalsMPHg5Q4e3Xjl4WR4fAN83ofBQpMGwvl
t5OZbw/jVwoK5OX1aETKJrCpuAImDW/JThLcoi+c1gJybe2QTjzyiGeu/U7M18hm
QyfmMy6nLhQHk9tX+ZTycDVHtsXKgsamOFSMnaj/edQ/YTgRVGdosn1XkcO9dl/v
Raod+TLL1/tjCc6KTnvDbYY2NHwMItLKt7Wsd7eWEZm/WtzJGfN5b09DdMc5z4Ur
zzvbdnA85q3ORuu1ZtfVeEe6UiBwK4r+2Ypki4QMSC/HobkTTivuE8kYFYbqkBRT
qQVX2ZCNpQwR5gpYWbxSr8cY+gUTrnJFvo1bkO9myPRB6PlEf97LzhtjrtG16rqA
EatyeTaRAF19UtMqyEfp887mUxaAbVTL3W6HvcefkfLxnzrKZJBd0xK/cjzR1CCj
tauIaMi6SD0TTWvXXBeyEyyoPPly4CxOFok6qERuE2jrVUmldtzULEepxV7GF/tO
gxwcrh29U7RsuOZLicbwGyLlmxmjrQUO9yX9+pOw/PqAyJrNC1qds9ip3/cl0QDH
HOXaHEx4kPFvAfu/klV+5XItTM6pxG5kzibF4vLmBwohQr8VB/h/3zXq8MY2/Mcp
A6peQXZfKi2tabNmlLqjZGON0T1EMfYM3WlXrIuxQVEeS7vR/cVtw96uKiMqvUHU
N+1sL9yeMxwR0x7QUXkn4J2Fbvzqy+tD6mbAdiSaGzMsCzQPxp/0wffngwQwOEPt
an5Yg+1etz6lkIKCAOTw6fKh7acfBhsMPaZPbL/mGG3hmGBhmmgqhcGfZVRil/ee
/yZn07QqeeM7+P5q4ERyfJc80sailUdjz5skSAIbjD35tP3/aIu4itCY3wyYcWHm
UK4Q9d2HvIhZRxbnEeY6ZaWOM8yF55aFgN5DK6R6BPmNJcWNmB0jieTIS8zfqoDz
vK5ZOClPbQnop9zi3iA5LuPL2WFsehMf5nsLIsFOPQLZPgACTjtfQ5fCn4KzQmCD
+Pq3mveZG5YwQ2z2KDgXCkaSPqv3r55DrOjohurYSZiN0XHFLG+2tyncZzWpf19i
TsShPe7yJRBcbLdBN6T64/16xlKz1Xs0fc1CsTFC4rNUShdvXHA1bD8cuxtHZpCv
U52EmNrkARvPPYPytt1ysoGSFrK4eihB+ib8lnYjvz0wDXUCl7rcegGN+kiUIggz
TN2sXMDPfyT962QOEFntJe8ub7mPry+5HWwAZfomdhhtevGGhOy9u7CVSx0ikcmx
JqLpBo7e/QwH/rA8uvlAyvnv06RVrVLluVmVwKPQ/mJpv4BAyZHt3FVIJVselcj3
gtB0QW1elTbzSIrggbFbnifurpm1HZiPvX1gfcPzgd6bjpqTeZEUdUmT2ioxy5Yb
91Txjt6GRN/Lgt3EEnLhzrkT3x8Rc5Uwc9W7msEpvdi4zJhzdXh+hCLXgx76VyqV
Ob0bIRuMhbTIoaP7GRa+Z+K8mds61dBuuWja3jDQK/mIX5mOhYOwb3J/MDsdlI3C
y/Ky+6P5OeBqTizIpwqbzqKD1edm9XBhYaqXmvw4QudoayELhmw0uEhHnYP5gHHD
zihOto8oOXP1Pmz10rRaGuN+o3fOBdUlxFl7TqtFjS9OBVD5Hl2P3PVBUpHNa7XW
FtGCEvdamNYeTEnFbPbRg+qDJOhpH3u+GbBrN6ZJG1hvn8FZ0Ft2cIp7Xk5WIR9G
5gPxScSLTzoPXkH4eDAG69XMn5ESrHUa4VI2QWr4qSHWh9BDrMvuYIAOOZ4eWrns
kcnzwjYzE7BpXZsWOTnDWm8MV84Hy/hNKVRTyJz8kh0TZiyGXSpzfsEgjTe2K6j5
8myXLpGhQviA541NuDevtVXewyMWZvghKGhLwxajLlTuRySIrlEqX9TNEZuW/agI
JvK3QGozMWxQlRkNDy5YZaOndeNj2tji4CcNDYSMhnlMOigY4vEk1tdRfVo7Vfje
Dj86SE8uZaLEB3OyhBbmUvdkDzk+oGh4BbNUZVsVw35fTRb6z547LbSg4a4nUj2p
ujmdMv73ZKkHpZZlZ9eYWsQMD9ACGXkS5yd09ii2Sd+TzmhGGc7QI7BnUIuX0oXa
5pGG1v0GbsnMfXzmYO4tSO8wWaGU5zCgHKkHoQH86TcUwYL5dU8dynWN8ZqA0tga
67PHm90ZQFpx1pk9yE8Zzot5LQj+gWXDS9vxKIH0y5eQ0rB0tVbvZcRTNie/4GT1
EegRqZmPnGFKJiu6FrD+BbKXGwi/h9iRJ/VjOXgK8IM3zW2TedRUOBwhJ/1BZcGk
c0hMuLp0SGpjI4irsGMITPb09DVjPzeOm5mhDdBAtTtfrxa+zOX6DQqauEejv05x
1TaMhr9qXk03YpRc55Zzv2ypPI92Zpu2pAIHp9fBrxqqFlN89S7UGiOORSO94KAD
l0pENBiNJP0wz8VCormpeO/vBPWDsahi/8GAqYuOi3VP1BvbJLtpU2WB7UfjVYWr
5JnPTsPfHWEtj0YX2/3kT409cmxtgLM6SuCfRew0bX53Ww4xebMQT0QwkcEK/+6k
iPL+unqps0X/Sbm7xFlN+TKZaHklyVOtM0SRr7k/6r/LMegLZvL5lcNU78ibSoRK
GihTKMUGbhvmvSMWzKI8075EUh1/+378uxs4vlgnMGpD1XRv0sp9FvF5EzbnwBrx
64r/B1A+t1ucEyDhCAvZhFijiSnecIhqIQHVc0uSZQpF+GOBuI1jIExBr32jl8Xv
DUA3aiScXEu3+BnXJJnxLxIGFPT1mQcO2cwrPSKGONpcpj9ufwvOx4cfbOsHRXus
tcAkkin7Uf2s7Od2Tdm16ns2/XTY78pRjpPh1z1IZZIied2zThmxTPP7GRrZvBnD
vfxC/jE1GRw7sNVYMbxyvfWDtzvExwnRe53QtpYaw7ohD0aqlneQGo7UANxLIniX
Ce1NbWHhofiHb8cKmLyrHqOUySvT3TzI5mwH/Fz9du3IpAeJlOj3HDxGJKr1FiBi
ERJSEYMDsifHoT0rVbhPERoMxlp8w27vLQRxmLGTfN3fev0QpVe2l6W/TT1YDbOW
FgVqDQc1BnoF5nqkc+QLsyMRMOQA6EPAi3DnvJ0iLv7hPBf4hC3Jya7azJsSEtji
CADWte2TWE1zBm4sMuuzZhdaQw2azasSD9zuE+e8R50J0tV+slFKCAFpnkuOJhsq
HC0fefp8UDFut1A8TdlowbNqmg9622dz2zOIIRJc6w3sOFwoGIUdWMc8AfBblHzr
Eyhn152PIvSQgLxvj7upmLtC56JcQv4QMRHoTtzJjPY3yg2k1MiFTng4UYBqzVSR
99CjMCswHMoYMcNil5snXYzElMNwSRnkhPgpC9/mkEblH5O4ENefMaXpv7jFIl3y
Et+p8jAIO2xmau4jqHbb1Qa+tNKzdR2jpoH5mk7y7y7T3ZMkyjQupKbYEw1FuiA5
p5otCpoyYPHUo1H0FaC0SwAPuynOGrRWXOSq57rC4H0M/JQz5/bfr4UYTL6FuGK+
2Tp+IxytiGzpQm7ZLPn3lKLqx+o0301mW2Zjq02aorw7MCljtvU1UpXSxkaqOJMi
XhZY+WPLYQfIiwvewN2O/+LusYx2/XXzRxfHHM6EH1SfZve13n43sNxfBj7GJrj+
nR6H+xGw0zaM6N/rQCYF+DTj8OinEm/DI3uDuLqXBjLACnid8SuITDk4Fo/xefvR
5RQj7xk+DReS37jrpBm3Het+oveXtIaq67K+qUnTmdR2rzVyKD4eZqPxZ7uCKSfW
KQZUzQ+1pp4kZbp//uV8DhhzPAlWgEoc2bXl8giwYrtC4mn2g9a9Y1nWXnTQXRG2
47j0YSM7X/Ik3dSzEOLGY7dsklUbmdx2KvtNrG9CFgzdOrEpCjiRvD0uc0BwrUdH
J+Cr5aMaAtdXIzQHigOWKPH9GCxW/rU5I+UEnDb790994JCpCDGSKMSyYL6CC3Wv
o2q+0o8AT2DeD5W+cyMoM3wWY7BBQLG651eUGVx6HGe3NohVIlKvccicY6RLFiKd
3QSDPkGOYQ5fRulUgScC1DkLgxN4Ah0x+SbbNJFHQvs1wg1zHYeTttJJeT3FgvhA
EV+G1AwbZC1xgHn60ttPPDSgXNKFWyik09RzGSeDVjrBG9ZubNwVAwDYwnnMWheR
a/r44fdgS8wbwwc7ymGm6BFxEl8tmsVJL9XgPm10h2KOd4hWqIZMf98jVxCU8wzr
V9NZlLm3Y0uevWjzrb5kyrw+rkiv+7+ABhDYlASWhk8pdxnJcaorVxtmErhHtV9e
RDS9BnIcWXPJt11y8qlTrTT9fu95FyEN1hu1DIw+3vOERdYwAgs+Tye7ZZdLUP88
nzyuqYVtVd4xQseOEOdN9y5qdVyJqyKuUY6uTvjfXdQpX0sC4ETz+SNc7gwGnNDZ
Kvg8dqUbV6AeUq7wY1KxdeQ2wD7TkQ7MuMNFDL8fszCgrAtod1oLXM52pR9THOPs
Kxgmny3yV4mfrYnq3UzroEplJHUAECg2u3mnedTixpUSpVRe/L95WTqyohWaG+Ii
7ujxdxpoUZtoZDl8kmXJXrdua44HEqA9soZLf8TPKxtZK/OFlx2ER3Gm4mapRtr7
7irFGu80lT0L1JwqOVg+I8TjjdHUlkkKU17H8wEa7MUpY7sgxl+l3JVKxARGvwtj
UCPG4oF8WHqhbFPwFgKPeq5ahd8J4gX7VDQbAfyNhG2kujv2NpYZ4biH1cz02n9c
UUvrGM3Cze4rkNP4AollHwHpuoLgtP6JLB0Et/QXarMXQZQYyqfahUES9BObmN0G
LCDU9R73Bpo9qZhgpqpcmVjzusi017tbkdYyMeDZ/nCppqKUPOjdHHCHpyDP5I/v
ksqbgTAt0mfet0xvTYvnqpuEhrgAG3F3ZHbsxtmYHcVGiEckNxEwGrPP2sih8yLF
hVNoTdl81EeiGJlbLaeA5uQzwSWMkw1h88KrCiVL+lrcXgVIRTlqGZLVlFdDQpRY
/abJ+FKaysLFit91LWT5Km5fZHJYr2IrCsuqgBXKTNYxM154eY3nRci1BqafWDs0
oEn/Epd3p6MzTN/SMxO18vArbQGxCIR0KRn4qou7TtMgwMJX9FFP05TQOtpUMhA9
7V8h4eleHzLhAK21cChn9T0LJHS12m9ya0dliHGG2gk+j/u4jOHCtJbI8Sv/bnhS
WVZLiUEgINeRW09nBJf/q9RIH9Y5p93RFBIJIJe5nSZYH24BKtLkZZ6DiIcDVbSH
QTd8fbJPMC5BBCnVSsOdgLLGzl16tIFMyrChOC28wUgVTQFSElzt/jkZ9HtkzRr0
/tGu2QwDqjR+8Fm/aHhn+d26lTxMMRfpyHmotU9uzbGXsdKtiu/350Is+NaCgz27
fC6MXmgON96y38bu7KI7I0ECwYkoBTL/qu+0cLOnKxrXT4WmuaeBjMxmWRHpZJhZ
d8fkNnUSipMehWEH3D4SP8pm4SJuiLZXNgSuf1bKxlK1QhjXLqrEf4ZOxc33spJH
m3jZ4HwmUpuzOwvgpNVjUpMb8FgT3XZi8cRQwhnjLPRYBe46JDVbTrDdQ/oiCW5S
via03OVTkPuaTiazn7Jtf/n9kg4nGlaw+Scdp8cL/mnk1nCktQ3BaFAJ3GvB9n+i
kJjkYaHj7wcz2lpiyycLJyafA9gdCKnHZZxsRbsioYPQz2HtVf321dLBnO2FbRy4
PUct1XXY976rak6i0WtaI1EsNffJcvdks5uG5PI6j/jiIFuuXl8tKtI7ZxsbRQtr
TqYbaEQKEl2QP8xQ3h3MDdKzfOEW+zd7IWSPZzTtNajdPEUh5o+0biVCNYSqQHYW
xbWVcT30/TpT4s4HXsockGaXyiOVwKabxQEE0mqAG9TFKjZkm9dexRqu/gx097ki
c57/BfnfbRWZDBctpLJRR2teAE3nC1zuV8zQZmhW3r6WbIR0Z7vGZTqAt8zgHaqq
fXmuTviCeFYwIhdHzCDYqfti2VYuaNl0yCILxxvrRM1WyhcMSGy5HQorlL7kwx60
W7CvhRlcQCd0z0C8TNc4HflrXWydkhDWZ3ubiuqMOYAEWNqIAX2LNbUs3ul/O9Xs
//AL31LFDCAiqKPJvJ/6+7vZGPcnrFq1628AMhf08dmQBoQdKptme5CAJFmH0NiX
NAY984X5FNAXR5/8OLx9Oj8wyhNLhT5rRRPpn5Q0XfqGo6TDSGKipo06Avk/gmFg
ndU/bpanzK4K14L3fX2eYA18wzaLTndj8hyWy6HbKZlJnvgqUg1CdBxM16BB3t07
TOpvqCEQDIn4+wSMMeevxD0XnmCb2YWaNduy30TnhZIw+iyay00JwOfG+VfxTD6C
W4AqCWsDf0/GuDWrJFOe8kMK/Fm15+hJSaZ2M343krTS1deqh439PQR0goaxzcpe
aXaqsQD7gzMvLubKaEeEiL088u7C866+5NgsjzITjrTWf0KCFGJiaG75pBHGmqKU
4H9e8EkPvugjhEp6+tD8zz+BpKFBAYxFzxh8joXN8kQKVnNYZ7T7XTSbWYulGr1j
HTIEHProeG8qNt7GNFY0aaa8pfO1yPT308Uv1ly3X6zsGoh/vk4UarXFf6YXZt+T
2AUZNHXQWynGYxNlbJ31iRRnQ0PwMOxPX347QuJLWDCquXsAJgOeimG3/zOQko8e
wcQ0BGY3HSxh0uS9qYxhHLV1ImFf31urPQYnRo5T4PXMp1LherlhUV7hGmnfSNmQ
7SXXm++jJ5eDDxmsLXvkLOelgh7Zcz8Pawf0N/GHDH8ZIIxA3Dq+sN585s6gIKfA
GcnDHw9kZCQ1sip6PCdqyiGRe9851/8zIga8TPjhkAJS0BAmQkP0d6R/YuX/OrpJ
VMXX92CbIssR+5KhYgnB3VgRV3LGF4nYSuqagY7Rk3soWKHtPlYrzx+mWdRIYHns
eLFOS/Pm+7gVrX4Yh2qNLBsmwIlBIQBsh+5g1KwAtKhqQo8LbQfaHWotlucw5bjZ
k9biJ1B7ZT87WZ9l78Uy930yMOxh0Wo4208WoOiipILbWgYci+ycPPKotxwkJ2Lt
II//wPIShMacnx6/EwWzD38yCzlTzx2hbgQv5woYtmxjQNDQgz1mAw80tVXMrUlZ
B33KThNi6PkFrCHQBwQxe64sa+8w/8g/EeM54NPor810g8SfnV9bLeu0VwFd3f5Y
Zo82Re1nt+Rba6le0y4WhBb7h7b+eHpaHB5VqaRvEuotOBtptF1oCUvq3HRnoKEA
C8GtRiUaIS9lZh9Teql/ilyZuYn8rmibnI3/JTLXNdKld66zz1PX9izlrT38sK+c
jGKAPBt23X5xDNK/a+IyDuuEXthw4JWgNlk3ZXryHcZOT89FjqDCUDZfrORBAwQZ
QOxleMKZeXRHzm+oD3Ur6t7/fE3BGdQ15ESglVoUhSxZRSFBHZ9Z+LnjBiXQ1wh5
rGjtJ9RH+0XE1XZfy1vEIJyyBnk+UXpeindkAL5SldwhLNm6ZDXYHInI4uwH33lR
w+XWRhLSmZ58lj2UG9YhWvOpOjA0BPonioB6EmhtDDCqalToi4I11cXcYF6jue66
+OgEVQbPKWDcBjWPPVxBrOOIZ7kWhky+bxnDPwtAII/OyFmj9hEZip2iYyXizYPw
jy0K+mIlRDB8kCP7bsigOPAo0Ija8gBScg9i5tooaGq1LHlJtReM3HKbRPOkFwa3
3UKEqie5GxH9Fj82hL/bcyxlOLLnvIfFwtVWg6CGOy2s1Frjvqm2HSSudynviHFu
W/TPB0mkKWcqfP7hC244DMvAj+Kq7Mels2Gxfub4ha0xv1oB/CYDONtak1KAhm7D
IU62g7dbUqdbf4rBXc2iWyUcPuyH1n6649T8tQjm1WXTgd6WZMgwiKM+slfindz2
F0Gdy7hTIiEdE1AkkLlVVPv6mTxvnVW5r8WEyb3Yi8UmtOzKPg2kLrBZsIHIk/mI
aFFX/1XvUAOx0WQnEXykFWBBnBcg57CxsDGbDGuxGcZAVz4m3dlMXUxhoJV0TC4a
qBZqrW3Y9sd7pZCu7Tegh3l7J198l33d6QQIjVTC6NyZRuWbxqr06wPveYgzOiL8
OSQrotLb/cJb/D6rX14cvkVhA+wdO7kxO069RgYuQgyx9+lGWTYuYbiEUWlH73yl
ocUBTTrCK1dmzZDLSd5Odqzml6WVVzlUMQzh8CFNtcV39+Y0D8tAMvRlby/tD5/4
eNOAOyXMiEMdCmUoyoyVe5eLa1kObjRpxaWVgRT+CPCnlRc/wUkxxr9mvKOzWSBB
4JjsknjY2YFOIEY8AyluNUH+C6uehzcid/9bTgjFGPc1wa5DfHy+IMZWdye2XozS
m6pTiTDePcfpJP//DmkODhOx+Ljn1r/W12vBz9wKC0LfdkpuX0ajiG9GM3WzTc4G
INdKg8SlS5VWKjPnZEvW2NtCyGRG4Nz8OV8Eaml3lpoxgjZzBDK+unNveQ1dly7K
+jVCO5vNpC7cOwALQBycqLCSCrrygv6YFspToHAoV8ODHv47d+dmzuD4vS5NPQXY
oSGaJ7dvA7xI9jyabKelDWSc54CEyWoQAVqb64Kh6MOKwJjR8tYWs+vAkQifoLu8
vqxvb2s8MUhmt8ZSdBN4BqueJ9HyKaDCZ9Eacs6wvNawzceKjcoQAYHCAVxRfLGO
yXF0dwaiakmh7DyHwImUqD1p+XeEEfmjQ2bgiratQbcaabnfYXMYn0O8LYpYjcOl
FMgAVU5CA/wFRBVlmWj52v3W6iq4jT5Gq8Q23yCh3lNKQZlKzn0Kyx/lWtXOxDxN
9c7C4fdlChwXZqD0JNScK1udZXSlekaX2EaZhcWiKf98rWWqDjd2c8Km+wQV98Xf
LQ3G+j5gBoL1NIPxYqlpZz7S7kcCr6qb4X32cFEQ4fSoW1axF1SQwTLS+GWkUGNC
wJ7491JqUefZqmOETJtIcjsrL+Trh4UMPTlvYLUMJx2tZ8ty8EHBkhRbgwSp++Lt
JRW/zMpyT59xSO8hMQNOinVbWuUzZXGRKYB/yobOz6dyAnjYGzCasWxDL576vmpW
pNPCJ3bDtBJfDnXWEBAS4Z+9MgZuLGYBn2vQQw06vlU3hYs6betk2X1Ti4enyIdm
0Avec+jslsQjTPOPbHyb2/2J5ynhQhxTN18nb9hoWSrI5og2gHjMV/0YGLCcBiqI
ffdSTovFL7pPwICz+V2jwqZnjBCF2JYMSecyWGqP5cGb4YLNgsOiScP58RT2ZKuK
XVyDTcsbHvnlzoUFEOfjpx0UWl53leR7Qz2ZYHNDUYLQSy9ZN1IQDLtkB/SrQrXl
0oh7jgRCm1yTn+Iqvy7ecK6yoYfNlb2Du6Yqqprj6rrfviMi8livbTbqpjHmuyku
yhREgwM0+KkEwCJOx/cSZ1dAj/ewbr0PdGk4b+HN9aTRmsNrRWGquzZT4rRgr8iW
RA4LPHIeDnBozM99hxlCUtqOAT/xHfJ0+0xw+sX3/CVAY+yIv2qjhOfSgTEnNGFo
gpa0apyNY5P1z+1YgR2ltIoHckriYgDphUusS6hD7j1P7rmPlxcKHet9wbl9qKu1
ZPUspcZBtbWpN+5tRZImui5j0ATfkqEeI4IlvKuHnnuEmqzkVnxSnbJ+YxKIpPQP
AOJF/O94tGEJpXZtl31sN5pg+mCUo9DC6u5EBc/HGY4g5qOgGF5RYXoJsQVy7kpH
u+pD9Kk7/1s9XG6YHXeZempKVPut9dTvE0rIT4+Fqrrv2zFebYDfXejW11kApg0V
ejhmciBRzrdqvPnioJCltKoc37ggR6nrI+oLBaaHprlXoqczOYStiz8kLEsaLMd1
2ARRAA4kPv7evvGCxTA/WMjKhjACK5qnCMSMXIQFqkL26i5AMNxQbxtEdqA2NmuY
Qml2FWhS8r12uvSYvR5i8S523443QukYgKp5eqEMAu1QF/ccoLX33+Vprs/lQ5Cd
gdUw1MUHP48ykZeMghYnFH4ZIh8ieTx09WeKGBp95e1qtLhZjngl/9OBSoq4ztyn
58DxuHm7RqSPEGHkZL6QucNaOjpsoSnoIm523tYkn/Og8yJCYjb36pjCNI0ZJqDC
UwFhe+RMicSlhxkVO/clJOqUXs6L0EYQF1Pftdx6uDM770P2K4/0gpq+4RWscPwf
a/v2Hvaz7tF68A247TT/ofXFhrEn3L3UhrCMgnGHn4HsJ4GZLuMnKofRkYA6ocaD
+X+4bG1vnjhHXoApKfkn+0bFVaOD1WEaZhW6BrDnWUug2F8AGBZklx2tJ5m1JtYL
zWSVwM6E6VE/BKCvqjoBXbrpZ0BhKc5cLh0AMJc4mQRvJ+A/5CHJUn21sGXxu27s
Y78LRsAygXnssXyQppcYbD5+v9fATOAXVglqUWzi/VYSq9Uhj/VcpfCuIgOEz8i/
+Ko9lY2GrYPgFadwd4Jsx5FneFVIQVKeRCrEaMulqv5CUu03eD5A3RDm3uuROobX
KkWmohAIzIRZnFNB3ZE9eA0tYBP82PmT6Oqnw5lA4IPnxcFHfdkgXWjg/pgeoGEl
s7u9uEUvs41lFYVaqTeWzCVKUTBGmDCVBk+UFzcEY98l/fU0hp8qHjm/e6pcnOEE
/y3AGS6kK+FEYoTVpAwltN+t4tYpY/fQ8EyvCtbkzV1n3eLvekncWnJNFDBXhA6S
EqLMg3nMx4foAiakVKv5dAkfnyYq+7jZ6MmnYoEHY8f8kCA7s6EG5/HANU0DEj2B
EfEjzXWQIrijWm+yZ9ST27HegDcMae0aszFkovo/tIYCEzGj4docYWmRGB+GVB4I
fjuwhfybMdIdIIL/vNMkG5dW+YjLil1J4VSVFJsJhms7YYzIV2rEsXXkaYbACzW5
aJh61Kobl7+w7wp63Buhv5vb7sGy7DFujzsrPCYy9E5Yq6CjB6SrBtimePnFvpgT
9/uvj+9iT+O9uk0jO0uNPWN7PzrY3xLqS4zFrmIn7zFN/P99JzfKC0G04nhTofWH
J2m5FeCuXa/2g43iBR5VK4Usweq4QZokxYwWHDI4bF7WjoA71gBKUzqFvm7txIEF
u0gnTV/4YKgsTz8venzFBT5WN4dJxeQ/trW2wyizHP3NpkKLhtDUAiZOY9rcKTSz
PELOIyZQlMSLvXRhSGSyjLRV3vNtKkB1LWjEHpBe3nxM7eTtU+MsuNfBIIoWgANx
l4uRmGsgFtpjmQcm6rQVEjh/lJkp5SN08kcE1EJexH4q5kosj8fNgHNyeddRIaZ1
Q9FfVSEdkymqj/zNmSDtt/KtTfbyOOy7e6usN4J7j4yUiV52ZxzK2HzyXkc/4Amz
AkzNPkSuV1dzbYCJTjS0yGVky94+DFz0EGVli9ES1DfTQBrqUy3yrhJP48CDAr0U
bRG70Kyyf36bTOyzGzWC2iN5sohKQ5aHGvxjn0z7fQTY1JSZ7EeqN3TR9PueTHZq
NQLVMO9ByMRtRBe+NWttsVxha0zD7MUwXmdt9qn1fLdFn0Vj6yu3wcEaMcaxGXJ5
+P3PHL7POB185D1C2jAlWDIEnX0x9/8a45M24Ko31DgBJvo10cEvKJReNe+1Hfgm
1JAJIpEucxIln3GLN95rMIIGQ1ltRSF1INL01k3oFFyjwzV/Yuh16x90TzkqRL/r
DsphaMVjD4yTUUL6ZgE9zHD4vXCGljTBahnL6kEW0bQVl08uax/qkuF8y318fUtI
7ucdoPqUbGd7VvPe8Drw3/9azg4+jTVfMSUH+817PQ3DZ9OlNagSoZdKbSd6XQv6
skJhyqtLGYd8vQoCV+tB+IiNDdZsj72w1soQvH8RvnJhMiJpBg4ZcIHtNUurfvKW
xZ8mHJ4j9DwyemqzGMIpzq4FLTP0DZidmDyCbjgsHsk/GRAWoONdPzbZ9ytfqbdl
StdS7LVKrjgCUF3pBZNDQTzZsZ9VxmKpN3IJrxucB7r0fYuWUBcQkovhLQzy3tcO
qQ7iL40fDVo3iF+fpBb1DxEWVX0coTchkKw1OoqoeQnq4MHsGH2iNMZ2UrKBagYV
OeLcGV12UnsmtxxJBApddUIw+vRwIx/3r01rijqaUJWAIUT+3wXAvQhd2JQvBbVC
r+aE84FLKC3i+VeUlG6kVKUfReYG+nGqSXhC4qVjveTHCHV/3JebWrn95LZIqSne
q0612TGZiD6XgqXOYLtWZvNacSpfv2MnrihzNqca8+7Kqqie3AykcosvOTLA8vlr
qYSEtaYVHXTH+uTpxKYJf9XruSUIy9ZDf/TFEDeoj0q2uqHJ8mIPcES1iG8zF53P
jbFK/Eyve3tc8AmcytyAWrTGrs35siJQjzCRxP7aIjgjWpkTTFTRTdbdXP8DjLUb
dn5zcJjAhh+YszuYKFk/uyxCK+sK4+84ll9FsQMbcN2rdjzQBKWvnBhbQJicrLvF
vjATCv4oNv31OtUJ/9MS4QLUKRn+1tRTBQ2nWJTGUi8Q2FCvU+wxArY5ImEVJXE1
gxLA65zrZUGJPxrMAWnOiuzB+Uu8sZqKiScW/KN5PJCrAkxVhayOi8ZtZD7x6xQk
KbSN0zNz5QqcJxauHxpNUEN4eDMqEgHXHjCmtCTvHZ3etqXnBnMX710WHEnHOq73
RidA9llEqbhiYEA3qdtQaw9BvwSYSiHhikFb2abmpB/hBzKM9gwcNnt08O8kaxzP
c+tzqsYj2xNTJ7a9PcG94K6vksgGu9QK0BvU7El0HcI5wqJQhH3X8x/9IR10Ll6e
z/b6vu8DmLk7YKv0SLvOs6GLHLBPohyOdo6s38XC3uZB3maMewMhtav38QiarvSL
QSVmzbBIKvaviSFoO6is5RDLCkCBUFzAebQi0Vp5HFYZR+3JbYdhyjMoJpVnLnIa
oAsC3XFBBwSn+M66KvpamEeUJ+tuSPeD0tZAWEdnKFvJg/bbWIwvJjeH8jPZsDr4
MTwPtSBUPd9Fm65EF5LKl5bNVn0w4rEBAI6oGWFECdeU43/t7eN3kp7aOdDPFKA9
5Od/1EquebK53uRLobtStLP9eDznPSsa+97WtPm+gqNwke7qQjRUUsEXog16/AVw
1YVK/pN7eHZKJNHpPA2sILrCUlKZ/Gp68wvz3EpYOpND1h/5S5KsZ0iPU1RVdMWo
I95/wayuZ7yOdm0hObUrRq/mhJSdRItKEylE85F39POuVw/Me4541hW9MLR6JiB+
fs4DVsxwXSS4tJi8KYtAMNDdk5IojKrQU+DRp30OeXkGhYYxR4C/DbbyNzucYAna
1zEgoggiPW4QUw1PPnlKcD/yTan9zt5AnZ6XAPFHPh9Wv+Gl0nFu/gTJCzFdWnHS
9Wca+WqeumgKg29oGPlUvQqOUYOkejIC8ZB+eL0EZkJSxMBY+5Fx10xASvFEdLrn
4zMXM7kv+SUq9EFI6O9I8Jq+lYhU14ChNVQCC0nJsHESnpoh1dLc6Krn7JL52Wiz
yPm3J1eOVoZrFkvcfzPmtj5L12/47h+oaBh8iongtnDNa4dBQIBm/MBM9o/WgE9Z
s6b68sZ5ToHJzih6MREOgcgKuQM5fXBa5vGNjnazbXTrRQkVILq7ePaxgSmvv+wF
Mqv930ciqrBrkYrGmzu8dz9aGi6BfUspzCxRxnxX+JRgagdfeE/nRk9acPq1/3Hb
RHrEwMqp67N7hPUw6wMqe0dTMkaZ1xv7Ye0HdllIa2+KVvgerp8ALI8WnhplKPNe
69ZniEl2pODJ3m/hW/Xb980I6EP/GeUV61VOSkkWfes7WnEkTz/wb8bhoohOqwOs
mLiFRqKoVcVsRJ7aiESBKroTRyyLah8YXYSNGXMerRRZyW5CG6Tl63nW05T09ExN
pv+KKGAvy5HJlOW/qKhsZA1NqrYDnMtIb47NwDs6Be2cLKRGYPhKpkBlV9bcg6fT
48sKNa8lzmGxpKc+KT742Syb2Rr7HXwWs8oV+VZ3Mdti/DiLIG+7CMUeY1dLfYu4
j0VC4Lnxxghb2i+II/cD0duEYU7MREV0Oz0hfbJHrcAZ8OwFyhrTXZLzL71vJ16B
1GhEhpuc8VwYY52wVegNz7nR1Hq+Jzfyy30swkPkgAGut4dT2DIBLNAH1sDKEY+Y
lxPnnj6mRvm24gopmok3ZvE9HwrjwL9l+6HAYQMvH4CuLlPqy07dOH4GzcCAjrMd
lom566gSA/MZOrOZavUCaHXIBEZGNYaeeg+qpnGnH0ou0R9+fRePemybQVLN9gXl
v3jmUw4hgaCgVerV+v+tIbUi29Ek1ux2qOHO3bWYDzLF4JcqzHZggu4bhhD4aC4N
lCblHi5T3p6xke9ln+G8HMiOEkKotq5WFRDzyPivlaewHnNikMZ/l4/iM4ghizWl
Bsh+QQH825JPnRAYbM5eIq+F0PM3BmFhMWyUAjwAVCMCndjvPdHOiXTzaJyRHJKF
LifLh5CvfiRIm84TR6Mv7owPwMS5Wqd2L+DCi147ZVS7QWrCt81Hhzk7jFIIDCaD
HWUjJj38UPCvO6R1PRQboQikP9jP2xhAjy+kYl8tdZmJud0jWvBDlVJjzJFaypaK
JTj7Al1T5GGuVTi7gochshJMToYWCMJtvzgwvCZmy6364fpWkzQTG5oYsAWEjD7J
dnbWuOUVdeEdrEmdi8eLksC8prshQCzZTSyjJ07n8L8v5hyOcq9zYnt/DxqXAEa0
RmWeIrxlOq4OJCQN4PW/BU7LTSSarrJNaI+7swa7DFKZM+pB8KkaHZt+TRLDm4Bj
msOfZ4+iN1Oga4Jy1mxEMtbQP4S8F6+HgAkmfQcc4Ij0jckuPxlHcsAPm14Zf/yM
aTcik8YUrcluwFrHrP/eqDcfSNCNmn9RbgNlfTzuaJYBZjQ62vWguR5OSQfEPr39
IgGkZ3vCHNvRrDC/3Xq57HAHY9rAk0mcjoC7eVAQFNQn9RV+/iML295/wXMR13rY
WE3mynP7lEkUypGp71Bu9gytHKSD3081hRK5Cl5hM477zpSKIQ9+yhAMwKro1u7M
Q+BQWdpMuJnmQEcLuXk4YX2jcq4k1qpP29WL5i+K9LjUEsXOEDb7mhOKPe8UYNmX
hBi7oNOCUO3Sxs0eXQL5e3OVaPcmMixEoibovXbQvc5uPgDUQhzJ8V1YeDG7CGrl
pkYSYc1rZlDWPL25RZqd8XZbo7eERCuBFhLDfZB60WXRuCuqtpjjEuvG7xEjG3g9
bpTPczRIUo3OktLzvribYnpeioEgrHHCscHqi6L/rFzdDBBqhkSnB4yRa7x4xBF5
XsaxgX2y9pBITOWkF1f2rPqtY0Nf105iJD+AYx0F4LMbEUoJpbfMD2xmY4mhJxpI
ebNB3TTU1ao3GAE55XBgt0iYJmQuRFzTo98MPSjXX4r4Le2N4xsnZeLHy4I19FBs
WL+sz1yUE5BJ/NnttvNp3zht+7oN9G2nZy71w93Vda2z/b0SsVmGYeBe5CLfhM7j
ykoKU4tgXuwZlaJiJCdruwNewfNjoy1/trXQH8dcOt1K33SGK87Lofa0h7rMUm2w
W4c6zfSuidSOSQiJwrlNAU34AIQ5C5KGWEnW5kBdtYqL3M/QmRWWAbQ01X/ow9tP
g74PFTDSoUSo7ZZzB0KclQm8jl26Swsg3tT9zj4FzyOymv3d2X1ZFpt+kbtLlOmV
DeLL8Xi0T+4s0kusuxiVSVBO7xaQ3glR5RQ9mu6ys5Np/9EkrPpX+OUieSAdBjBu
0NrQx0Tvdw8tJQnknedhDE+Tbc8wGnWh1yUnoL63cBby4YsqvUU8STC7ZGP563JZ
BNRrIlm00qNcUSEps6bUoXsvTY3zf7plo3t31UwO5LrB3glQwYxhV49oXGyqqoje
fia9klJ2n+MQb+zdITe/1j0saxYJpTFYNzbMLhT4gihiPd+HOJ3k1FM4m1ooyq5/
a2b0VaKTRlJrX2uetHGEnvUEig7orLUS6+QVHt4S3t4Y4eHrpgcJCBm1ot2xvhi5
8SogsCX8cBslQeJIG09IO19lIUoiWbrSb9DGeOb6D1DUA2Tjls9KL5udjAH0Jeft
cDATuqXxRQZ0VLXcXJoXnbY0kmlE16uYGtfa8YY9TEZQa1OLvZJ3gviNwAprxYn4
8Wh4c0cF8tdaLmOqCXbIJ8L53Vls6g5w4utFq6YeU8DQmqqeAtnTeTq5ARr5WG9n
l2cO822WEGomm0CT7AbOVj0gZPJfPSPDZqMRCs4j2dYxNaV99lw4PP8WYCf42ZJk
APXw1YGVpqZ5hq+mcBf7MJWRTHRI494HgkjNdZOSrErbaLVto3YQEwSYbQP6auu7
8Nd1stp1YR0Kd2BAmexUhHbSeMex5bQ60JCvc1iKHb1sb5xBCE9KH7av7+0p6EFB
JPwocm9IdNksvlYV9K8CZ5P/pRjC8x5+31isnCpStE7z2ey/Q3Z7H0v0KaOyhA62
1m3/vjHNsoREkHEI9tDQS9etTlDhRj6merP/2Q2qXv8ovU17uk+7rbOdJGtFCguw
AqkHtQDuUTVyyXbr3Wi79+4DK/QUGCzV+83E0+xmAW5Ss/I2gxR9xJXceNHYraos
4Ssq7sB/glgGEAY1dEv0b1/vfQYTdISNpOVnZU9ob5g3kxxV5CoQVs6jRxymkUTU
I7LOLvqFKqnEOuAQTday7d+UO/78Ap6XVh6SSaUs1hUBDgvT9OXmvGjUjx9w8PL4
SMLKgic7THT+kBzZDjTfv9gJpjWiHq1UX4tBirQjFDkxSf4UrJujwMNxuQ0hcYZx
iizl89vAV3aQQdZEJ7lCJQwxNbe8Zy+JdyRZXBGBZ7ZUmGKf6eSIsTVJV9iwGvds
a3ea/5gv+7dVrB6Xlxsvt+AUXOC/HpGaXhx1ogtslvfcBeu/XcVThPl6je9AxOte
2JDE5V45S1ojv3UTrql+qNF/r9fVGJqcW2dCLeVPI+a9zXJRGGA+PuKj6VVmVrvc
2PKHpVMPLc9cET3/RUKmXHWsYzXrRjD2DymFX6eb4BuRljNVkfxbpv11HNhEa5g7
2uYU1yjxY9EvIIKXdOmq9aCKxjqQ9TV98YuD6ncP88BnoM5h/Uwdps0IMA1HGECm
aEF37LuvWHljZtO4ic2Ja/mx+bWMtYQUXSeEt8dju/xGqE0xLuSD4mgHuvp+dnkg
AVZL+rLZu6OGZM5cL+Nmh+GfxNvB5H7nTvsXWVwOX3Ox/N4vy68X8OQccdF9yoRb
gZvNj1xxGVIbR5FI5ozwL3UkA6nWCTd4242CHAFLvP1GX6MdX19pX5cizFeJrjZF
l348ZxRgUrzpSLygcAzCBP75YcAPHzcna4qM+/nKhLMt8yuDVCGqnK2zKhfy9GN7
ixbN0yopzTnmLZ4iwAajAfJnBxiU/lhWFzTvzl6CDFeAqbo2/G/sIt6ebwvwlMqg
Tyu7TvNAoFq9ECTVI3HbBgtJHO/ba5G/aoN3eNSmVTPATb+KqCjYze6ocldS5Zmd
I3Ef1/cxjpFn7v4lZFaeWI2Qq3cCyEcCJBGwtfJpFblW4aahSlL/dPIH7BwAY9vX
N7aTrxrxlS6MdcrvTKu65XVC7CF2K8dfsBkNaOlSmWUnxeSTOaoJHRCd06DCzhqg
gTnF3TP7FkG+r8/8KYZReMN3RhH5HNfer2Gnt8zPdY53AxMvxNUvwmSNA1UmGXD6
cSlSzCiIv7oQuo5qijHZ17rVULFasz3t3VE2bh1KI8oKiwOF3a0h331Drl7Ox2I7
rxPPf/2hqwM6ZyiyIQ3oXUTIkYb8BaXmcA3zMYpjy3VOGVcu+Crfx15TA3NyFmkz
a6kftRRvF1WYuMptnKhiB44nZvcrHyd7yjGphu2wc5/N9wu0SBlaqocyLR41+C9e
/Z9VZ03Nuvo+UON28mr82waGYswJu8c6CFEBjYYVKLD/eh7AGAUNKKzqm4KKt9TY
iDhGBzs4LtleU3PyBqh+BEvWJSeG7F7SdGLo3Wg5cJ7sLCHUq/okNhZzJFgWH8BN
GtqvyE+2Mf/yyiCkssAnxO20rTiC4wxmqMgy9To+mVta9YLQZnQGlTID6zxDUlnN
zlONaF4uRIy/iC78Vdwzct4wIR85vyKQy7bLA7D//ZYyhRD1kyCCIcxTlpnONKkx
/8ybIccp+UpNKwuKJV/3Plfnl9cOPr4BbgA0g5BzCiNCTqnNsMmAsNE/j0+OLovU
dF58KbaX4HJZTr38djZzqb6JmOyX2mMd6IVGl92er9wSVaGj8lFLGIEE5MOEjSeP
sWFQYjaES7JQ5n/lD08Y/0yFEG0XXBNpd7DjPGjj/E8ILoz4Z5Gf6SR0NjaFRxXK
o7Yc5Lh98rseepjzXHioS8RxYdGEeqAoTaKfrhfv9WCLCewHLjouTQqYrfKEtKE4
0Bvhw5dYHZjbOW/jzZXooOdrPl4uK6+LHAScMOryTOte0btsW6Is4og1QeMbUYtE
wKB+X42sJWmru4aYbafSXawUfbLfa6j1J2aUQJv93fdIfsX5fyCPRNgaNmzGHdcY
x3cv8EUgD0eFXc++K4Nxgnj5OirEO0MawZlUbloHXR/1v2cXwl5q1t8Wb5NpOWEU
b2leDWPiyrFj37IO+z2li9BOCOc/C7o5bkLi8Ttb+8YQdZ7Y3J+/htjkDFHadDUr
6GhjVTJZ+YficyWA2Q32v0o2L7y8H8adHfw4dv+GWmArMtv3czTZzFsgRjgHZyU7
PuL/tvaSIX0x6lNOvAO8aeheK6cKTKuPgehZpIWn21mLh9UXaAviT8M3M/f0u5Cr
DD4h09Jm4f0sYuSfJBgbECTxr+k4JJOa55orqNH5Lwqbq867LFwxIBe1gsEzf9iU
92xIVk+zvJMUBXwdiZphHnmXWvcfT1oGQgdrpJW3nNnA89RZn+gJF+uxl9rAc9JZ
28RO9xrpoM/SV+Hc3ajXo1askUxlO5X88MXTznGbm3jJEHEmfg+h0h5x/zz8PlGz
8V4/KCcteF1Np3x0VVh2nyAHPRnOo5JSI0auh1tvVP9zNNb+7KcA/MGu9l+gpGZr
PFPC6o8DDWyTMfQCbDC1ptgYplWna68AjiLoC9mWrNpEHrdO+vnRPyCDQBXQprkh
bgQUFthc0eyvBgPgVu0qGIRK+PsTG+ZNZMsJnR3yUKKeG79wjDZ+RWjr7sScQ+E8
7Q01ZlBYxyQ6wF4TMPc2TiJ6CAeGnTlvkDBTjGj+TPVKs1W5HQijnOzBW7RLyhBX
sRCNyY8rNlGB7Sk4ZUER0pghVuZ4P8sE5z9uwo6fprfujAaY5w9K7YFEzsZ7qwqs
Hjm3ksMIHEv19APehJmYik+9TzwLz471oPxjROUhENkPxTPFC+4Ljld7LLf6fRz7
GNsWPtk9e0nrgHqA9FgxS6rg2xqb7dTxOHGA6bT3aIqw+BUWIHjw79bHGoADHCRO
Vsq9A3u0i/9BD45Xh4Ma4YRznCHQkDZUeIqs0lMWrIvbaKJLMmXq58Gu91DEj1Mk
d1389+WV/GbYX30KmP83BrlFN/K0B4PmxfSPMmKUePvEStIiVGy9HLjVuhZdhhJZ
5CH7vLVCsRXGrCJsxLIdcRLa2BNk+ddoPuXPAVuBn5Dlhg7VDxUJiGjnSLteQt8e
bjZe8EQLjVnDEru44vArIpcvb36maUOI4bf2+qTFFzGYUC+8nTwic8NbfeAXXdj7
WSsTtl8zzOiZpRUl+lMsBSDgr8AQUn3/1vRB8P7mrYInD9LbPsb8mXLNeaHB5cNX
baDektoGXjERYZe6y3LEZX2OB5YDUTts5nizfy/6udxUBq3Usjx6IJxFU4KM1Z0I
m88YfJEnJEavjpWXmy7zWDyvxT45WL76atn2qtCOMB9/vou8fWxkkqVDZ9Ran7CP
zKkb+5EAPfchkg59HCB7G4TwQ3N6DouW+ij0qrgQLXjDf7Fdr67Zq4hPfs+nMKkq
1Jr6pSl8uSfhzoaAgH+NSJLwCPJlH6aIZXyCiMYHCxCgBYuxc1lcF99ErQWeqwym
A6mIQkeWvUbWQXmL9Q7U4v4SjSiQDtx85M0ac+TO6zrFPiz9KOvA+5Sn06LcuLwG
vhQc+87bKrPenJJmN6DrhKT2BTxge8Pco6gbmOMf/blvYqQRl9z6QwY5Tzw2o8in
wU7jAGO8ESN7lVF7GvE95XJDF0jAndwnuuhnx+R5tQPLoH1MnYgEDxNiz4XJHAy4
wKRPC8JoOTFoLQmGUfiu8/bCqJmYDEMYjgqviZaVHoJ4YI+rKPdF/HdM5T3v/cdG
RcZnnxO5FWzxek6zNwO/wi/SOOB+uPInWzB2D8nHGxwhonuXUsNIouUUc21aVPR1
pLcb7DscFFNDPBZwhkWyzkGtECXIzm/XAs4HGpmizhqAY5Mvgdpj6yBnV+vEBO/b
t+zsILBVObbvR/yHbTIXUzmG/vYTS35X0tAI089seHvo/cc3Sfk/zSfFxvhug+Ga
4Z4d0qUrcZC0gAmZkk0nrZ+iTom/UszpFz7p2nku5HFZJdrnzmXkKCTNvEYQqqf/
cugXMQ2jhQxghpVGSserOjF5+DS/se/zbxSYTNC/P49b77AGfBcagEVRSjxdB1zc
QJzYQ52gUq65FdThzLgX+7fJcMH6/xYv+NZHbBmH3u19LIMiryYWi/zyxQpZYh2v
JfL6THSLeL2ggl64E2v/DX8iPbISm+Wdxr4gn8nDHk+lWEPZsTgbDwFvlR8eUgEa
L+PBQkQF0kmIiBf6L+SL7P+dqXgn6/uvr51TjGaJ8qUaGIZ9GeUpvBlnZ6GqoCaN
y7mXl9LLSrwlt1CPBko6XFopXPPEMkPtyKRGOsh2e7FT8d15dn96OvS1Fub3bvUe
+GqdIGmNA0hmjBG4s+IKrA2aEuZ+nFbBhcOdXAQuRRNMAPsx5yZZmBRZYwOV9eb9
wDUIi3GBcOPqbmEWNyL5fbn1rsXATZGYMevDn35/wSbstxHD8fqewi9wZP35QkZg
JoczlSxlJHm6bwEDNZ+TlcwY2LvWfIRhDDPkY5e9rqcR/dpK9FRsB0YGX01LiVFu
VIoL9BTgnC6XjBzS1pgGGFMmbuBUqKmf04EmAQH4oiCv6PT8++d3Xdlz5MJYc1Zc
GFJYdmcxhTaaODy/gFeTwj34LntnS+cM30Q85XVZnHKojQa702QUKV/fCAMw3U1P
t7pM2wziDi103tdviL1QAirFgKJrql3Nt11UCIP7XIBF0dfBTMrHIW6kehPReSv7
GEzW0gq9a3MSWtXaucUYGWDr2Egh6jsMmp3yf0bY1IlGMUiY3PEHGBa52cXEcPvl
wvCcRLVBMtsCiOmYuV9rbMAKV4zEMhB1hFKugnmSvyMbY+0h827MRql5dTfylFIb
RpmDNHFm7eYgHST9XYviVh5bvcswyn4LNyIdXNKUbtPAfrKydbS0/o4XePEX3V03
+cZiBVgiss8M/Hc+y7LjqBK/v9TO3SkXnpYsL+Mubp1t/QnDVYo/ZyTYchWIbDCE
dEQZnKChn+siB9GRdpJzq59HL7iTkyh1b+TZd7rhWQBdrdNwhwD9Iy5rgQss5huV
sFHGKAKFNXXKJtbwbgMIzCOquU4Iw4xYFN4/zBpMGZ7bcGAXK226HbQ6Opj7azwf
Ta+9JXWzTUqBLHAI46GtLF4cLa4XbyIemYWPR/bSDPosYtNNWSBGNAQkcJeHQVdP
Nsc65Ld89ie/RxI5hQ5t08munHJRItSb3jM76qpm9vblksxMPdXhiyhxLRnnudan
bnV0rmkXmR892BEC7Tl0pbHC96pmS8BfT7zr+ecGZ9EzLklIJW04lZN6VReax+Hj
mDXHWeh5muIajiv29thZpeL/5nUxRUlOwd+J57HwOPM5yQk59/ExIIWLidfiK7/w
CIFr0enUidrYdnHkgoxLLqZgUwx60e0sPmW0SX0NJ6hPjKeUP1F01a0YLe124U23
/7oKCL0/D+RacPJLpBfqKbfohxs47u612FJ7okpGi9dTCUAfCMbnmWdi+n7WpI10
u9lG+Cita9FUzj4eWskiRrA5e1FI3fkJ8Jf2QqdCVEu06T6J6GD36NcAgiBUwoxT
xIVCCY8O7hem1Vgf6mvwdnMeCi+iiaCCc6kJi7Yw5hWtg0SKjPR9x7rfgxkapLnB
ScdYrsLtZyl62CMuDamwjO+vrGam0w73NcSWd2IkU9V1w0/ow5QduBkEQuYORM2q
DKc5swqI1tFYaAOfDsK83KzLZfWJI2KAsnV3unZqN4tv0SXZNcOv7zl1jsENW5eA
gruSY2DUsIbg0tM3oY3r2oPNtEYanx2Uo/kohc5dE5Qxh5IomQvP3LwJODRMZfQ7
7MpAiFHq4y2niz8OQjK6ijuQPXFmaTwIqLKzVNufWDLJG9APmJwW0gvBicN8UZSc
tTtk8lDli1EACfU9Inrzfzey0WZibBw9itWcconeCBHo+Ec0zFpP4V6FUWzgiHuG
UpM44II+amwQmGIFwiEEMlUTU0uZ1y01X0yqtq6fKkYkv+Y+iqN7Z99JkwzoB7B/
LYwFGP8Nd2YGi8UE0/WfZqHvgGVbcnp02vFhixptYQvkXltNloOIaMTEZK5pbFOp
N5x3QRPft6V9hmDOwyMWMQ0T77fTTEFQX7iKxvR31m5haQIwqFu4hl7lUlumKlv4
4nuWzbDrm6Bk9HDMAfFIDTUOTwCQKG4VLtTuysFrWuVlHn0Bo1NJqsiYbRQUF9/8
I0O8yFCrpySTcep/0iCKoaUygMtp6kUE6vfQk2aFRb85FOFki7gVYpeQ6p7HPbTm
b4iCcF5APChXH90GCpe58tznyhrytyxFP7cmdR4qqmP6BR2G6ejeTdKm9xd9lDpH
hanGDNCk9dWFCEU8PoSA/HyYi4qFe7ax0xFS6wgKWWdsEm8mUq3ULMTI9kTehaOX
iwJL3ryAwdvOfcfS1fUPm/ea2R7D6qgeevKZbwTpR+onN8qgFw5bbvna1SvCXde0
ez50cmUI1UYNIOA/BRbBgnz43/2CJ5iMlPGL3XK9QQNXRsnaVSapJmgelfV0oHZl
V70RbJXuq7vbh3DmWcSEDGv50WC61hoBsqJeEy467kWAPx+szSKEuZyZ+BXEULz6
IHehiNagZ1Q501Mwb/Q7ksUby/5rQSkFU9VsvsiIDrrogvSt+Qnyqyyvk8MWcgo4
0IMqicDv0qGILivsIs5/1Lxs+ceDHVl2Y2KKdtByJFDOtEYSN/rMksvv1W3xWMSw
2xQ21NlJWRbnKVlnofl51gh4rAiq7wDq847/2HPz16aoeRJ3h+QCRbDhm6bx85GI
zrhzRR6XQDViTDgnCeUnwFsAUgbJOMZEg9yJBhlZ7d6ItjlRDku/KOl+QJJ0GyoN
LaQQrvKL+52Ru7tIS2ZYEvHwvPC1UBWENjaZkurOeYDboKqf4v4+1HR3+A77NTqp
xkBFcapATvYkvp4sN+XGC39vbrnVl6iMqxeNwWqoZQTDFFs0bMZLSKvp+znkLmov
002gTXNSQXQQ+N+IcKuzgwIjBWnOLIdUcDbw2tXszaDfZPvjxlacnO+O15Kyv2Ix
CFt5WeD0RlDr/uhz2Vo4bUmujlY5N355wyhCzunlIMEZ1GcrLVd43P8cZ7H4HN18
qj3xdZdfj2xEZ0MC6aMZLAuqI+NDN5BjbwadNO1O1AKqfPUreElRxL79sE+4tID1
b/tfHGfukj854C1mmv7URVeDbVtmR3LfHa1fpg5BPd1huHtCjzrUgJdpUfIuJaC1
5oafev6m7Ck+/EEG0Ru6BELMfw5MH8da6ESbrCQHw4ZU2dLQEWFUr49SI8ogzPkL
tU+Z2FDCjbNd8MACU2FGCMV59S0xcIjt15hk1/9rnbJZkFNC+ax/TJg9g7nYJR//
aMyl9UqSBq1cpBak0RMvU4A6ENrF14QgoSVHa8/3njHwxeZygx6X1lOGlQtT7N4G
xaiXw0t1eImi72HBI0o7lCVzE5/4foR0Qp04KFJqyVRoveNVIxT2RoovS85eQ07k
R9xXGSw7kugkDn/H2BuHYxFZb6JTrVIdNWF9tB7KLXWBJ6sXjZszEi24Wfp+fPAB
0n0GxSpF3+oYyUfcuLVXl9qrLkooeVLoxjNbJnFn3qgv6EIHAf6fHwFMdqqoI/N2
4VaY/VVRovf5QFub/W6UAZE0yMGv7oPUUua8dQq+XieWfnKAu63TvQOGv6apLZ6q
+a4//V0uftjT8f+U7SkYxOewSv82BCGL1ROFiaU1ktxGAA4K+ATwdS9zKUJvHQxy
X32vu2CLsW5iefnypNsMEwJhdnczQyBEKfcIXWd/YrptqJodlFFWPbAcCLlXY6BV
FWiEy3pG9rThqqU/5QRbm0KBS4mzYQSX1A4YUWybXqxIGrJJWKFOEA2T1j4g4IWm
2QdZEax1vmshOOutvFj4n8K1HkzSnSbGvCBKTHCqcdDJqo5/s+JzWKpte4lsb/UR
7acDLSyMMiQbCvQlaAFkbJeVKji6OkpIgaJAyPYcy/d2X1D8bOyrs1iqngvGxBJr
A2vuexv1zdu0PGC98/rBRFsAjhRFycZqEVAngq/iWmKq+kf4JHTNdqmkuUJT8zsP
lY+7DiT67PxywvKp+MNBG6PchopEMfL2ENgZupQjXFVRaG6ezVtCFhtw4rsp4ws9
KtUhL7NsOi+Sgbln/PIrBJVLkwzQJKqbWt/8vFHKOPPAjMAAiUSwvUXkKE7VOOXV
iiFjDj+Iy3nTSeGwV7CkBkTPA+aUYW6tuvR5KLH4Z4Xp13kqFFuxAORAfjF89rbk
BHw2v3/hiZo7QlP6MaEVJ1EZ3PV6xThYL6FzjIbdLhVG9MhLqOw4gbuXJ51ha4mF
Q1Yl4x2M+KpIpjh6BUomQMzQxHIMAXdqGkRhrQZ1AtTk7+CFVGbyhQiOSDjmIczq
zr4YWkF58ZpIOiw4wNG0IxV1v6cCftFW9OY5U14W9Kg2IclWkHjM+2oDqqkQSjVJ
R5U8KBZsx9Z7HTq6y6ZhLxT6S6j338QWuVWqIrhz/14Zgw5ApFJBtEDTcVd3Q1Di
B8uVNS28365nxAdST/SxOe5DSHBJDeWSfEL3qIElu+4JGteNxnBUNgFb5Ywm/F1O
rTgtNhm14NpoluU2/3s+j0bAuEVRX27U80sGQfzmm5q2wbZSWX6NFuzuHBPX/gi0
xZoQLm92nYnmLpo+Db//9QIkNz60zvNXcNAGwH5x3e5B4dhnMkFhKbNiGJ90gOfa
96FcPWwC7K6/c1S9fiJeZxlborjyHsTNONgWPbpvBHNP0HXUsYXZpjDpx41q4km0
nDMBdsqDdWS9vr5zr0WdkiQC925TKLmui3JuBVA32GxyOLj4+ZxkiVG4uAHrggeJ
oSPD6385VsKCjk/lbZ164SD0ff5ktkoeVuDUS6BWrla7YnkXn84IsymJrWiWynRl
9Tf3mKDN0tlFRe17BETnqGA5pEgIb9IdnJjN+LegVrcD02CHmFSaXFrC+kqaAA5g
hJpgj/LkmPaSAQLMbY/icIhA+05FQHmB1cxcm+wBHEf/hDN43Q5Y+U16lq0z0Yt2
jGgkAP6B68lEfQSf+tiEpX4SDMeOqGA36cQJfGepArT+n43uvQEZ2vA/jJ41Ec1X
xSeIxfWcZkHMNrcHlq/O7AvyZeAPCxBjE0zWWJrxnK9l9DStO6DsKamYKadGD8BA
4Fhxd7FlNexkEOfUTaG64J/JIg6hSRoA+oJFn5sw0kcZPs4nB97yyRv7AnLc/755
ULasfQdZMQKW8Y20ZgsMbyoZjY2eyxbmzbwWucKmXe50t38BWt6HMEv2hJ8xHHzq
o8i1uNL2FZEFRpTpghv+mojXRFRL3rGwV0leJg7QB0mwERpKY4qK8LFlmhqCGQK6
xCMFU4IDX6eKzD6fhcRwCGdiDpORjz5Y/jyHtAdrrn3I5zvOqeyN1xXrH2sZwaV3
u8JSbn+2cNUxpy6xBWEyGS6/TlkoaGuA8UsJm/GtkijT/NjouJeYYRqP0WAgdllf
dfZBIuZMX8tIRNIjUktjPnktPDK2Nulp2NbzFK1u9n+nJzBG1IATaG5DAiGB+nYo
k3Bv1gSSZkZmpqY/PKKYPPemJ0k3nUP1hVT2SMa3NdFkrcecgMf52MHoHhmu3WYf
fP+Qp0WcG3xsaamQuurdDWezjMxYdb/xNUyvwKrJNhlh8I6ccbvHtqkK49QqdETU
CXLynKe2oRxgmoiQdwxsH8dCy0UvVdivijGsglfJIrFal4tApECx+Kv0uuTXNFnK
hv0jbayB6ZZpNyic+GvB4Dk4r6iLebFAXorBDa1C/2yCNAxRsz8KemFi6WNOYizn
Pqr3fBezWwawg9+h2BC6nL4/HlgWe5n0Et/xcXFWp6ywZYqfXxRynmVjnIZXPwnd
JnZqwJZASDr8vla4GuKS5CyWWPSqNJxznlSeFZODI5+EHDLqZnpapuxnOAI72JYe
Xv886rZ0tPQaDY6Sh3P1k1Y1HBTKOgbGqf7VW826hhskDE7LWJRBqb3p7FdkAFrY
D9lkl91Aap+0pSC018KhJ5+7Rv92WP8+W6jx6Bz8rSPJdNxP1m7prTdn9RI5t7Cs
SU5PoJAaWw+V52z28GxlndJVlxO76Ztm8StvD1Q5dgR977wiREjyijPaxjdTq4X3
2B1sdgdMhqSqnEx6RJrq0El1abbXEX+0ERhIo1fLBzU6TTaqmq4QiIcHr6Pwhien
fW7/nVz4FDngglM6ZV/R/UVS1kC2+JIzG9K7+KXGrEqtsAZO+tBYVdgPchu4VHbd
qPFnq7y8qhJ6Js49MWIK2jMClkQ25qrN2O0wA3ujOa/gnMROxJQziOO6OHUwSYeu
F+vW1zAVld2q6iWKZp6pldh82MC+h/w8yjhT8npe26w40plHijuj2LU9/rJcTfGX
Q/aHf9pWnEzJp7pD3wBm0c6nwYluPfF4h1PGXCoo80JpE27LM+tKR3BhZlnwBPxB
BnT/YJLpOvvefexWOkL72lk3lojEWz5/GOzCA/8N0ELVu12kq2vePJMZyrQReZt5
/1HgKYNQSZ+OBlIvbIq8ZUkPOOEPG7by5oO85jFSeZLalVOkiGj3E8CZt7Afpkf2
0aJkuDDuGPWg21DzcIEClKFn+OlDRny038XV3+TJa7Rmh0yLffZ1VYqzy0kDauwt
U2Aw/CTiXC6p8Q/DW2qtqNMTe/TYeKQTAnCbpoyFVXIsU0A2jaOwT+5QnZgF+cup
NaYRrJsEMd6ZOnXBNWxdPc5xClGRcmOM8RNcWrfHInUeLX8nG4PixIm2WWusLqEK
6h/SpFxIv45D8lDQwHxIUvjHsuDEYDaFMz/uMX2u1k8lSNCX3EmiskimdY/6pzWQ
CjYcSvFYJiVQsmSmEeuBzDr3W6d8XYK9E1m6pyies2iinGof4jFMQlrUR8encvAE
nJFzT17L0fTtovtBiR12QgnK8D56Bik8Tl0Hzxq1Ac8wcSZeBGvGgLWcIy6rHyNb
+rw0vyyBwGtcp5ly7H2ga0Mm34Rf30vZLeUIxeSJJsoosQUSAspx2UTV8U/U8x29
/2VcNFy066rlcUV11ZlE8J9eONZNBV6J6/LUldibUUA/1fUZlvv0RQ8yc3G2gKaS
CTqLyDiblOCgdImXBlkkWnfPprzFc2miJGhI+F0tFMP9y2/jhhS1Q2f/klqFhpgl
WkHLk/rMMbBhXEiqOKsmwrVVPCq5977V8gmPE/wkn1iC/VvJoB3naw5s5KC1+ZAE
duqoOA8Yb8ORrmGXZCydp+JeD+zd98K3DHSDz+QmSGxkWav5wAeD6y7OOa91rUxP
ywSBT+K8KDDKRHl1mnjqL60CdOtZA+uuqE/P3FJyQqWb13TRCLTy5xGIKvThamMy
jeysYz42sbqFk5qxAG5+8IfpUf02vGPhzSl5+vZ+vE1wAjkK6iHMWHeF9+1eTShd
awB0M2R/QgRrMNvbxB+SkvTW5wTv7HJ8f8Vv5ZoBSVGHLz2Qhmb6suZPbax+PBm9
P2J04/neDMdmOtOqJMh8QeYF9BtLyw8pwYmrG9uMxcVLBkDQgSi6y6gBBAIlguDI
p/TEMAnYW0NgVHMHbwiviN1/AQhns9GwSYEdOy2qYrPW4mlOiGVQlnTI7MJDb67E
rQg5lglaxtQEakXsGZapgu0yLflNwcfEvCe0DoUNmP2tsI5aIeuiNrROmgKqaxQg
uSeGamol5UqyDSMVtfhfF8dUqp4HRYLnUHx2XmI39t7CKR5tW1Nr3fMIsYXo9Aj3
O3aOudrQEtjcL7x3wyCYf0PuD3VoOzrB6dFaXQB0zQBbjsV/iRtD3gxUV06ulxrU
fXtl8TxS/e2o0D+6Q3z+gypVSZ9iLLEvFTGTx42C+RmhIOTM/PDthglMT2HKufNy
Nnxwk7/rrtNfPAWK19anVhZro23j/o5rJorZlLHI2bTIIBqIPPsWLJm6iVM9dsIa
jLJENf+Us3M/IOS3ZRf83cxjOPi31BWuQjD6cOULPIcBCkrnivhg3r1glytnnbNv
pxkHgzvPZawJFBVPG5KKgn40Kv6CUFs99YfJ6e6cpXe4MdeLE+g45Q1PW4IwrFHu
y7lgT4XNNL5omQuoISyAzCfDZuJsjTEVIWawwLIf04SzPNxjtSco5nEzqV84TuUY
sDLuazksRYSj6FEpAknTIa1pHr+F5i/mxUT9GYet/2zexHcscd9cVXzqYoT9ZUiX
4ZotmqHAMQPIgzTril+H/BZpLmW48L6WoJ9LZMj5qD0MShVXOwFD3YBcLZU+Fxro
5UG/Rx97iC/k5HRnX4U/YP7Y9DPdiDsaR8LcOn03nCmfOXnDGSVBjYsgKB1Y4EES
mRj7/PKGJIe1fNoQ0nzj5nYecGoIE4hjKYYxQ+a+pP3DwXXpj87J3epjwYGE3W++
Iami4AqLH4t46JK9q9BM49KHpe20bLcHaxMA996r1hviwyehO6hA5soLZuBQ8faz
21HnnaQIZvFqmXuSwtG1JEhPJWFN7K25K3x+ai7Q1mxOM76LZER94SzvEjX1YvbB
61dDu6vmTiQzwsuQ7grGzBGeRrZ921f8KP05OKLW49Y1GV4d+MgH1PnpWa3CVptS
twoY3nQNxUKXa03ktZnyXj5yQMRcJyK+qzvorWEUauxmmT7e5QMP61kOapMiT6sv
r9mUC/I5okrC8thSps0uDDnMli8E085ox+VXYhNz71/tU6uYO1/JmcnkyDonesHg
5RJd7TcVlI5SAz/vl5Z5BUd2NqFS5NVUjX3H+ftw/JGVmeoDAIDP/fmPA1srTlmX
QQlHyqasp7FCEHtFd6OsscOJVI5OikpB2jNTC3/VPXxphxRi5NIYNql6k0ogIzXh
t8xgByZDwmqNDEPNMVGNIPnrB5Xr11XR2TrHC7ekkV6bI4RHHe0c9E23mIUUTe9k
ZPeaHriAi0OKbKZ7UJxm8JwD8knapPSf4fdjbsbI8GA7yveF2kezcbTt8fzwaERM
MzEugun/vrqKME53aWga/02X/Ub32PEF5qUBF/semF46F17kPPzlhUBq2h3n/hGX
6JMY6cgIBVTpK31PGVG/+CZqS26z6ZKcgqCsn4362KzURMnZOyAlCbqiU73XeBE5
86inYkHyBLBlVfNn3y8ejjaXOkDH0F9uxxVgLeCkzrf/6ptN+bfvN/WEB9dUU2+A
9mZ05e1XhEfbpIpe+VjJv+LaOwlY2wTSNRR4tI1NPo/dALz3oQnmt5shiSVY9B6G
GwzA3VbqOA61fw2dGf1bWOs9qxQ8XbNjcrvGiU57zHIUJtIaNjCBL97AP+oZnDeT
2BbxAatnT4RK8HxtVfrJ7JxMT/8lCYxKRmQ4d0UKp5byAEqkJoHWaEfPSkR+Co22
N3bkOzbVDtWNxUsfuIbMxX3Ahrce+APEcRuASTLe4cfFL6mHWmd80Nc9I4kd00/4
9yYveN4iuRMdioaEHuiTB1OXJ7SomfVrNawxnyZDtlilmD2Q4f1KO1XGPQUzLkg/
y+soiz6dIPEUaGzK5WyN8/nIL/ZTad9m4Z4oBGLJAyIjz5Faa1mhD3sRRC+CE3xq
TuTSRyEfS93R4jkAJKBJZk8Qoz53NeUZRgGbk55+8KXHacrdHfrr4SzHn8TLwvnt
ScvFWYdkXxt3eZ8hIvyOkzmqrxcZ/8cTo7dLReAN/JnF6IjbhHZytyp6QaExzAHJ
HilLrzYproBXo1V4hq7DTlR0sJslOJ4WsysVRLmqaH5U1skyHC0Qkz5U1AeBaYgN
L8Jc22wFF5AMiNSd0VbaCFgT6/oBP7KvvZ9z/F39vpDmpaVgSkQjphkX8pm55i6Q
2pMPQDwR6c8jRhl560CYb2ELxH11EKdPi4Hn3vvsEvjr+10OKpqtaaY4EJvGw2OM
4JPlcFtvXLX451ircoHAvQAmfLEINVO1V/t1KeNK29kwV0KMLMwBtseQiyN7Wai6
PGrPV04IDf0BHsMOA+V3PlM40sJkrBmTeMb8/vEAPKp4+5kXP/0iZgllmYofItLs
O+onmSiV1WxAI+9RZE3Lh7VfRbrpARoewGvucciH0a91UM8RQdPk7kTYB0ozFkMh
Yr2Pm/ZGL4P1cm7k9LCPNpIvq4u/NkP86onsi2UmrQ+Z6ukPmrL62Pz03ctGI23U
guT2p2JwODUWCBR49dHFKKS7cLuw4ilL3XhrtPAx84l/WYOK53gGhsI9/clq+7AJ
MrjCDY+mxMZd0bCS5TEktLQ1SNXcAbVDA82a77eI8ATzT7TrkhOIED4k+4bPyCrk
H/kIokxqstkXSkaUiCbv4dRj6TkYWFlNXlnA7gqnB5gB7lJ3pSCv+Rv0zxoiR3K7
h7vOYhx49a3Sq3FrgzRZA9o6Rh8tQApYBzAG6HafmXqMywKzQF4OdtZvDR8c2eqo
vVa2iB1pz5hLFbco+MIi89Sj7/fAmgJgC5F0DR5BmH6H1vk3GIezthT7M9ToKwrq
gbkxQkHWmYw8AKWho4Y8nIhslBkU0xcYoiPCUkvw6HquAmX5nYkF79eFCqhujsF7
oMlFkSuCc+GRsdTq12ciVt/RIvUNMbc1P/2DH9eXLWmb3wtY/Oe9mXM4PA3kQyqN
uSjcJ3CHxoR+pF9LyHtqwEdPNku1HxvCDVb+/NOAyeGAA3XnNcsO2WUwQDJK3ztS
OK4p1nXvpYUf0tOgjEYZUsDoLz1ErpoimD/ncPTBKbO1uTggAx/TQ5bu+6AINPE3
uU/7ayc3zhOQTkns19gUIJdmUI7Z7CJN6dqPwtxmwpcqYzCSNRCu3bXpHB+NaWqz
RPb+HHk/CjPGKWKaT2xRYkLaoMSXaURGIg+3C4wtYXIDemtYLw1oUg9Yvcu2s8MD
26ctnOokimioV9FRg2shjR/wxfjhqhZ487eFH+E3RopgeG8m4n3+dI7fx9yKi7jT
4W7SN+ft88d0jKUUoIk56Eer4U+zx3x4zKFo8tI8ln3VPC4fsteuJqR8QoiAV5pX
mDjxvH0OgJapAQV3dPh1eTp9NRI9VGJh08KsUM43PGAVcX1ehflP9J01KAFZcGlK
0IqQz0ACeKbTvufDoMeNS3BvpSx4XddbHsGp0ACK3k94hwI3v5xBaOat99k+Jkrh
xquz7fxs5Gv2dtGmp/M+YT4bzeAwALI3q9FXbzuyHjKeDU+hqzK2DY10jyYCCF+R
9j9mFmN2XU3T9/uLoRrrnfa+4hDUK9AIV6HgkvbhknuiL/Sc7LVUz28sl6OOXfFs
T7PaI4lRUtWhH4ArWV0CloZlPM52udq3oXuRL3Ro/e6aF11YrPzVNj7aI7N2YI0l
XMB1+QSBzlTINfH1GX5goVGWhUIcWu5XZ4KzOwoxYKQt+wn1vCalEMyFTue6FDiW
FQZrwXDUvCilouulX67L1ihqg3iUtq9j+X/5/NIlBFwjVbkw0zr0gKgD8URiilNy
rDjGrNQq7bJSpz0MmRfi9mYmtBldeXjZGY3yyOaBaGvK8mwApGyZa/s89XFAHOP0
AHAdo8oG9fMmHiggtCCsLHMdKOvHnR2k5t5KZuP7x5clq+akjcytV2gRH/oDrf01
jpNYtxOAx/4MW0z2UuLNkkeUK5A7A6rDdpfsU3+UNUc/fKdgpI7JkIBdj1VoaUev
gm3PTerdKhC6y8+HE0IiobvDWbHWwB6Gboro9kYkuvhSdUOxdue/1G1ZmlS2f1CC
QPB2t6BjYXQMmHuO6cSq5vO9EsRV8y1M6imnwk3I4X2qO8hkiKt2m9rCZhGDj7yo
U0+CxArpPGT6/+66UrVY0dvMJ0uZt6ac5Pz14Rck+bgKWwgGdo/Yx+O7kbma0Q5i
cpv3ydB8RHb0F4JGSk+yg7r656boGrPs/8rMsgIL19FETmLGZ1piZGGBit6AdSXC
8ira6bFWNVqTs7wePy7SfDtRENtMinLgSRQKe8Ew8PM5CKuo2madOc72RQx+nfZ9
vlnI9GSslcM5Ohh0N2fe+LlOvYIahLUS/RVZXz+V/P2BYCOyJ3ykaIMMC9LhyZFe
WMHQlqRMxhOt9wim6wXJPjtjFTZE6W0K6dQ6GNcAlPU+SMx9azkboTk04FLJywbE
MtPm6rZNWZr0W8Ugm/8Z3zKd/ySa1DZ1ilpob7ZLXfMgabl3OY8XNJ4YftxG4YCY
JFqhKnZN/wgJm7h12y3XmK7xTRqG4JSrSpdlvFeV9lhdJJ5vfhtiLvyC/Kd5nMtt
uUa+dPp4TsVImzcbeQNnxL8HhKRu1xuKhZG64ujm2mKPMSg/GtR/SQsQ2Y/DU3H5
a9XvkVi3y/5SlPMS+xL/EjijM4CRDi6TPkdI3Jge3M7sEhFr08k3vuu0yE+QoOZ1
CITy0aJfA9IY+mZ8R0ymo71Uk4pZ0Xk9B/jiTNsAuDhsllnFTdbVUjauDr947tPE
JQk38GEaJokve3AuIH8NimE7LaCUK3+s5fWDQbBuoYJlwOfDc7un/h1zlWkdYKhx
gbPxkzPx229nJPTiaARaeDy7WQcKW22pKxa7KYUSoryzRParOq3Ul3+tzcFYTY/Q
ZKwZ2tpfPDARJ/Ee3ac9NOvXk9TMUJVdEdLDx9bkCF9w/gSD57G5kdkiAGI4RtBO
Vh3pSn7LSuB4nszv+S9itW1xbboudc1dwtq68OqJIMwcld9d4zNSpzYChA30c34K
IaquoR6uqKuAzZUDQblNzXK7289C/EZRADWUfCpVuxZ5EHjl8myvpA6QuXikp+rl
nCAGxM2Sr7gWnGn6aehZdA4S5MXCC0jyzGk+3N6oH90TnP00rNqnSwHHsQU7EOG9
F39NNUfaO2kNrRnVbzR3cZzCIwxtI0SmKHQCgqkBbGQwbAYR+3XiAo1o4GKAFfYo
aXQWPlbs5W3RiI2EVTwsx/ypUem1KrRUIlj2c8ACzW2PDgRDMSW8Ot8m/TviMPnT
JSuXFUQjfwxYLWiedjS75YrPvmwSCgBnzwx8U4/xngnkbjnMnxvi4dVxSKMxavAh
SDqbrVvGHyuR54/5EBrpDTBCadEKMh6QYeVRFJ1gKSR52S8wEhvL5G32sXQm2RhM
lRQ3qxVRxJD2O6U+OjUKEy4RBNrH2yzsUjyxxYH4LFdSW0kl2MzaN7Np2qLAAuFm
xfrZK8Ttzldfqp/giPxr1FayDhErwYg6SPOL0FQZKmzpu17sDLy225fBv47Tv1IS
AfHhyRnS3J/XQ67Dq+JXlLsUHWJWoiq5TjpOGlDySA7eS5/S7TcCOx4UOY5LZVyZ
/H3vhIHES7G5dGWZObXSLpa44ZN4mdBFOe6FFY8LxUClZpkq3hC6h3BdDzWeyP4i
q2edaA2gQgzgum/rdeZSvqjjhEVWAoy3oPgsf3DOPKIcx+2YO4GcwbihOtXf56dX
5Bh+hV/W4lAn377rxdxdRrbW38zQbk89zd0/3alZvPIs4E+WlNMPqytt0Vn2eLeR
TX+NA4mB2BGdaKp4rgKbvk8TW9rrs8VEL14FjoYDRqBIaeSIAksUdaXfRJJRrPnf
6OLQ0AC+cSeMxzdezsBB/OSNheuHcbGZwFxhKTB9ETQNmgtZvt7cbEzrJVkyRlVs
wTGz0gjlCle2STQTdxFc1iiSuI6YU+s1ixnju2wwYlsQr3b3xSgoEE66cBaXU5Eg
b6h9EhcBgB5l01Hnoca+cBh55q31gQKUMcIO4wwnF4y04/b7BWFMCPxkyPzmnTKa
T+LY0b5mFEOSVWrIcwOxtEwczpNtQpb4sgfjjbvGCXIijgTbv7yT484FQAGyE68z
54rivWdJWZb173bH1rmozGn+Xcl6cm98Fs2ocaXzOiSkxPmHa7P9YTV1GqJyixn/
iZTv7G6X5lFmlZyFG8Ijq+0uFy0iAWaaVmiVF1he2514HGyi/HS9lH7MaGhLwazD
nxb8N6FaU+ucZyr99VQllViGbE+YZg6/WafnzBoiADRewRt8n0AkzcfRGe9Utf2r
3Q4HicredFXZBYapN4ZV9k7lNzGhpBWjM2ifCqFgL7XsQ9Vem+qofbwGjjye5o1L
u3G/2ehOk4FARxmdu5/OnLm2KfK6yhbbjSqaGIrg/qeuTbibiD2Kpo5ivWiSuWVk
dzuaXtmRNrV91ffx3vIg/AIMQllI50I6Q9gEmSfPkTkr3f/vw5KeaOOy6X524ugi
qowyWpl29AHSms2uKZJkU0OBPmzVCnjMYOhB8FRQzx1yJ65ZwYpop8NSdBml7zI7
uAL7TewLDkRZx4EVF9BsMGR3Xthvb7Mhgrjo+mNHGnvndb4Hi0Y1gomJiLCpYTBc
NF6UK/gjmv1AQNUn90/xouLm5hm3IyyRgt1bszuT/iMl9ObkmUf1RAMqvNxLJCp7
m8a3vhJsMPCXmFg2Jhq9HoP7Sv9ZMPwSku2OJjDjN2VZ4wzcQG3J9FdTFFOZu9XG
UMjmZSAO7J27YoIvRT+Gr4mrayr3FhRz2ZiXlzOInJXKXkqmlGb5uMKqmklO0e1f
yPIy4QbkboQRxXTK3Rk8xzT9y3CgsmZltII62cLO7+aFEnGmVFDau4V9frboNssW
ODL7hCR6gc078U/glkj0V25noQxPlESunm8H2/gMVqnuSBO/GDE3p2EFP4lKZ39h
yySaV7JEzsK+PmAIRE9GgZCb+Wg6qChjCNzRWqZ0FP0HcU+LLiVDtzoKkdiPzN7M
yFaQg2OX5LVfN+l0i6kzhZtq/djaD7BclVm4aTh1V0kCrqi7/v3GzXPxJgSStlLd
sUcRgmY9rkvM85H9Lw3ej2thS0l4g0eoQ2/mU8IJvRyWsPmvygI+x3VZ4PVIvfX1
lRw/C6ruI4uYxh4cXeG1rwSpt+vEaQzBuBglvDa7Q/i5r2VJmQvpfpeErBI/RHwL
VIH1H4ue9wmiOdrzUxjwrkqzcYrboz7vHtdkGtZehDyEkPGq89rWpiEui7AiiUZD
HDNR9eE6suzbesOHFgbtAQaXHeeYmbQRQUGchoVfIQ1wpCDGCp1D5Z3Q/DmKnBKn
q0sArM1p4x7gTzbjjCvz79NFv2Z27hW2YSy2Ss3QIB52GTCmwxaEDGzmUNfs7l5M
L5PFhn2UFKkCExD7RaukEHw75AKB/rW6gB7CmBhkfs7RjiMi3CKaYqctBko7W7sD
xYqDKXDOCLZwMpl+S+vncLIBUY2lFMeiUPhyQa2oTgkif0pEejY8It7UuO/E5rV9
CxdrVsStOqLjUcISAFBZNxBP9wX4yigZr1KuPsTaOYB1rMM/1lproDQZG5yWQUBt
JI7akQsk7Ml4Mv1lChl223IIeKh92hG5fi9XIIorB0en55o0hXtYYT2jyRT3hAtw
cM3jP5aTT4+K2SUad/u2LhspZSS79XpatbD21Zm0KDODalj4FTM0FrEa9zO7nhpz
+XsOXlcnFlvqGvjb1NU5Aw+p1Gv6604NO3GCS32xDdHQQYOH4k+uKtHBCzESIA8/
kNQk5nOhS77l2d/QFPgsywQ96RiFZJmvU4VRPxTSiaam+diz08GLPDvHmC29CJyO
+UaDkHX7L3Rif72KjvOdbEBdRYtVUiycZlUnzcP0muBL+3l4J36DcQ6tqS0ieOPG
gCeri0jgs+b2A/epAF+IKbaoIM0iyrJmbkE7Hkg2b937zUlxZZ1mBGrccs1OzdKE
U5PdyAROWGPcqfYnCIwKRZxf1Ofyvt6jcWrk4iw5/6Kwc8NcqK3lRgy++nA7I17I
onfuMt6LlutG28Sb8Q9kBBY1F7uCxCb2X2u7dayNTc7DM8GCv2gpyFaSNtoC9WYG
Uw4xcT/7ncdsRsGAgfgwWiRF8wBY0DOW9nMPIeKIsaHCU7eKdK+SrSWDTzN+iUj7
mMU0/cm6Zn20sGan76n4MjtXdrquTA0L3YQAhzbc+pilZokxgCwiPNddsGM4RjsH
srH0kBeFk7RH6XglG8JNE4QbGnXNgkSTSqfXror41bOkfo7gTz/He/67D/Is9ZlQ
DJYTR4r0Pl67BFxy/Q+rOFAVkdxBTQ8yzWdjz/k4IIDBOIivkyfeAzQqPuItItHM
lXyJfYlZp13wRxPn3b9vxAnyTMsh264rgWuS+OPSmgaDO+3LY06Ah0M8Scycep4q
P+CYtddEDj4HSYnMpIZVdcQfJBIhQ8l2EFtZS8tjB2OEWqqSipL0R+uxtdda5Vak
3xaWqNov+7Xzu6QWnTDp0VkvgwbZYZ022XF44R+6XvNizo93EaRMOfJg27Jw3H+z
TH3OV1I2kWgWAN6nq4h0HMgmszgqBy1ttLW289nOvO9fYpx9Y/pbwVe0prudxd7S
qDHZ/xN1yRqaGMrvQPJKY2TFs7YiFEZOSK+6V8jUonckIrPQlV/z4g8L16Gj0Efj
GWX5y2UfTvRTYb1y+ZBpAEWUY8c9hl+T/TXHPQDTjqqqJB8ZPwf9w1SQa2NddjCD
GQqd7k7Y1OhO1xbl7Yylq3NrRb2IjxeZMQRObMVdwYbav3KTXwybaIMYwEL75+T+
FSTubgZvRzJciy/xshCxpNawbypjE2IQrHlvq0c6+Vbc3DxFI+CfbcwVIHJC+P+N
OCa0GCHXZPtkOXSSX19LpWtCHEHvdIX+BRi68CrUkxpdjlUnAwPSc9rLpBVfamOp
aKQ1xVOlc4T503vv3QqNORjO/TAH4vzttd9+fClsIMVbNIymuL0N+zP9zRSfpoUb
i9N2wEK9JoAkmufEpphUKubmY6HRebigruvCpB6dF1yZpM49iHS5f8hiUYpGnoUX
7iCaWDaVSP/7CCAvZXxSGKdJsYre5dIvnrywgdhtxYDVyrG5jOLuG5PEDptJYdGM
ZH3/Cp0B8Nn+AgUMrijFoTdH+4xCLlykDRUM8L47YM483fQiZqVzrPqoTOHs7/mL
vjskejVohOk7gxc8ccPQt3LZz/Vf4oZ3D/ejK3M9op123lOyUGFEqWqAO+8SfC2f
mz5Fvx776paQdqqDMDv6J2xkFPSdkFpa3OQ8yk6kejnvf+Zt9yc7GSKiCf4pBVV3
jbIejfCSCg46YlmAxu8PzwlioHbTQMcV8vKJkoLeUYpDrd2Et+Sj1zxiOpFb1Tzi
PRbZA9qTAi/CLxveWHcmP26fDnJrNkfUDPpO4b2sfpsrLpYDhDdWM7a/Bru1NqAK
OIn449/Y/HNDThYRXUbYog0yw0wziZGu69u05tQB65l/hlk8Z41eEkE8aySBJ+so
RwN6es5varfYW0fQoLSlunP6OjofAmNF8G77zKM7fhts7naOWOifOMxdIY5FwyqE
za2lJNt1AcQYyuK71lLOTUmoW61iNYJOTrfNs6IM43CxSSCJArux1Z30c0d4jl2O
9cCncqysYcIaUtcA7GHuj8oDiEthGDjtPKISp3G9vtAjVPFyu403DU/oxY7K3dhl
hMkYYfNOLjylXnu9mUcdscp5JHWQtDM5h3sPxKKqZbMSrWYRjZw/1SR9jFcGgfOx
n5Qf5tS7Ix2FQa7d0w7mCbxAEAediY85qKN2YAWfx9RJlpd79xhfcstosIRg0Hkn
faoKGQ3RClkQeInNxA2xUVYHv2MN0QgpU+YBw9SoK8mNVu6Mn8ELFn68MN4Plsar
f6AvakKgaixNSDK61BeMPHy2dE62w+2gAMPm2KMEPJtho3y9NRpmAgGjA0g6YFAC
D1q+PTTycisme8FR0fDijG6rfFwYYrAYPmGnB2TufTmRuzTs3fytmLsfacCrBDp9
c34Td+UDu9Dc4Ic4f3jCZtCXJpP40SYxTmHU99l2hTwT8pisuxJaT9O9jVXizPXo
C6dTQxsj1VyLbpuHP5/mevFzQPalMG3ww+Gjxc4DtksIEM8yjqxMbAf7dfT12V+M
NzG8fOfnnH00OO78aqdTslYfRX3yQvKI7jwCOCMZ+dYz94Q+Kk7UNRo7pBn4VZ5j
smj5nob9CB3WUULVdkeCAPz86eiSNGBRg1TG/CrZCBWycinaxHMD/mRof789+Cys
gHLcScpexfNQcBbLnclEmdDCejvsFSOsK/Ekk/PV5jEhV6r9QHZLG+PcnVX6Gif8
XWSRZMQHRHvXKksAAM9EXLpFp1JElACRrgHyMfn/Z7txtgeXGRlx9RRDVrNwIVFT
2PHXr9I2jY9NpGv4jRvUH21k27NHnMOcZT37hgdi/xVljD4ky2AVlkjnkBuMUo84
s3Rn2w5G8uvZ4H7N373vrAoEchXDwK7Cin+diY3nn3DQ++ZzPpUrvW4aIOsGUhz4
DooB49w5bbcQI8lJPnMXp3bX9AMfXLI/2Gr3PnTBWJE6BUxMjHDugcrrPi/Po3Ov
A61mvDUjtq5mNiLvBdLbAjp48EV7BTX8IgX4kqF9fiEKsuJbzraklbAc8DGyDwO/
Av/w/icq6RgazXh7qWNgPjBHQAApbY77lzSnmlW4cF298rI/Mzz8v7XuLMpZYZFA
OnFWYa/wFXm9n2u1UhLA573/uVdWuPzDXIpHsuU5KETpm0vmFePImxM4CHgXksSg
Xm6/EBdhUeHi31fAxePVP9LhgFKRrKO1D0Qw4Mm0VthMvwhyUXwa2SVHAxF91l77
9I/bYrdwFuiymk/6cOwp9ozWlTcPUQ3YW4n/7EINZF/6lfGtuzlLMgfaXy+Fw+jl
ruy24lGMLsYTM1NFWubUZo5FuxWsF+aAsHGGhD1YsVZM7+P24gYeZJD4gaR2uRWY
OiVUKBmwHgQcPlAkThI4JLfrWZUgRjvalI2FOLJhtXCOhj0u2wUua0r3pODP2aZ6
rH29N6/UE5ZMfmfnie3mqJ/Fr9XWyuxKIp2QTzzmD6j3r1kFm2SAydCtKY6BGdji
n1bYRfM08OZMv67Pg5/MFeswF6fd0FBurdYPQEbu0CRJb9Q4XuGxt5A2NOqrFq7v
k2zoAJuTn33+MawIWaWtvs9y1j4+bbPw9/TTLGkV6JSIrw8IxXWtkzhWSLynOc0p
6V9GnMObE8ST/u2kDxlBOQlq0b7CXzHaspeEqv5ul0Olp5/4z+9R0XJjrD/BsnSA
jVHQ+IHJiD8DJVtMslBDdp2TCTJ/uCdwVlEjayplplHfqePcf3Bh7fH4BzWhpgNV
smajBz9ZMHP1swU1ABA0/piOh75xpj9d3VGNoSloKccGA/k0CgpHTMaxi1kKikmb
2LavIN51oZRbH7qskjjmtwATz7BtmV5/xXeCIUJ9kwJYBngAhZp062vjLUgmnaIa
lBZlE9e7f28FrLlfH7QHl9KNbtBT7aLZieJBG8Jp1oS6GDYSFCgShdQibL6ri54T
IgYMa/bl5zXy5PaedrgZgaf6qK+c5PtdM+7M/mKzUQ5vMu0Jh8MIv9njpaCCQzwG
yg4tLo9k5h2IN59dDlK62+LrlLHuW6w7qtOwDJuwIvF8WyMIPjL23WA1LWbjIqXD
W2/ufgBJvAv6dfW/qiZNCHO9oJlgzE3bTcPi9ZO6WhMDciTxXrZ/fttOGx2hI7gj
L733ljz6FdcO/3rvYgwUg+Q1BOnY/M+n+2xkI8gp+vrqaYxVFX8u8/gez1nwK1aX
cZrF2gl5aKA3/nLZZhzwQWxsHG3cRhGRyE0qiR4B5B/vwvivHptNHLIP9TI/RtP6
0wNBNRzSTKxFYIWeU5nmztS7dvh2fPRz5hbseU5QgBfMDXrxar4aHAuezOghD0cw
Ogxov4p66ZnrQX1Fubm6FAmBz1gqLcaZkI52NHljEr+wi+xhaLhdQF/4Hqi/4MfA
wB2mhoXgJYFGhxGBb7ear57l7vbu5KSnQUmm2AXe8fadOBBfiUQ7UBGn8PQVDFwh
Yo7kmHENGOwh+8Mej72OfYlHiw6eX1j+8xR3NPg0/sAkMuEKJk+U08WxGcVdBtNg
yEmYOTVTMEKhIe6Zx/clrBTSWOQwvAf8y5FqwYjSKN4/PQG9Fpiby2/GePpRgfkc
ZdMPmvbDQgDeDSRTF07PyQDrlMhpNBC3LKs6TQHwWeJCdTjqLozp8Qaetlqya5+z
dVGG4NWYCX28TbFnhXGWL493AxFZxFThlLOBvb6vVytxXrNVzy6MAkkDY18AFVkj
OePF9Azq/6PzXlZH4IbKei+3iM2pTLUVBpny3Yn9qfloNFZ6BnObVHOi1RAjWU9+
jWrRY6pjccSRTOKrB8Cz/iTXHCM2dWagcWBHuSdftKMZxppr0ER+Ji6sz8TrH2Pr
AfoR6q9EM96GkJj5y3t1CpGZfWVDWykA5so/vg4ux/OtzujVIydXnrXpzNuJLuG5
JQtEid98pI4ls7kLsRNJTmzyth1P2doCPQz2fQhrYxddlO0cpq0+pLypftol1ogQ
rKV8KCku59lzAw+8zK7FVR0C+8kzkm/sRtblcLuUt09Mi3TMfJW8vTU6HN/zzhAY
hChK1uxCFThhS8EECfLwNUXrvB6p9z+E3MgYIuo0eEVTeQhqu78x+qDl/G4XIqxF
qw5LZz2XqqeWonSPb00DNohwFO7LRKZYnKsxvFzN0c97x087gI/mA3J1wd2bHS/D
qLHDb9Qo8Dii9MYnM2/f5G1DaVfgPfUQCjRkU5uEFIkT/D2nLsua887356LLzIvO
XUNizTF1hDfRMPMMQfpkgElarY/DkpLs17KnTNUIpEu4U6YUC1PmFlDWuXPubNyX
vn/3TcBxurqqfX2Oq6ILHJugEpEOimicGJ919vZowJjflzdWricG3QH2Rny+N9uE
I3IcSSD706xzxuiLKsh0QaK1AvjxpfARyczpJH//8iQA12M0GWA1M15qWqP2KHQK
j1cyOPBOClyvkmYedOZN2Ayjyo4nAOsYa0fRhWUn/M5dIKZm8OFWZZC87KX5A/KF
3yCG/9oVA1rSpbhy8+z026CZyh3VS3W2V21ZkzaUJyxAZNXyDBqcnHi7Eg35+hE4
UxE12SFyeBSfUE4D+xuw8CnBRtFAJGj4/nf6B5FyYxj23BQPP8qY1xz8cdX6ie0z
Ssdeym9aoOaB+cF7wg2LEheEJqW3qPmivPEPrhPSUkiwGAgeS3g3b17lTndvJiJi
FU1PJA85K3pKkxEIK+Mcb5yYKdWVYZcTgUx1jDj5D0peVmRrvZxiJ5vSq73fLWCs
eRFhGLz+iWw7Ev9nGY/Pu0DdXWsJvz0clevWIEf1AiLFOuyn8bybbEIJACJ0+e0E
MOUgqw5VcwKsDBMEEFCg/n8xuuCc8NAzJ1OAk3h7/A8VeSGyVI8vJDDasyJFl1ZH
3UVPR21tFcwImaS2mH2jY+xIwmrnfp1mUbi5JPEwYXlotFocAGrKqwK8Ej19arNv
hdEs5fl2OWn1aqcjkXKVvdFrof3d1V91vaTuobiuR7f/TqelgbyiQUMFlBJifoir
dL4EyFgJxj4lvXXC2atS4hUuTjI76inpiPS2A0tbui9fpbFO0LubkQGI/Hrz6H1o
mVFZutz4a8cVk3NVowvlY9avps8VbOdm/5vZtobPhSFjXF2It9Wp9RUOvHIj8GNT
k7aU+G8POrQqs3eW1p5baYHT30kyHf58W13sC2Icuf2a3AcemmQdBZ4rXrPbr8p0
/9qSWnrPUnQRlU9OKdhWcwCBDf0+skU8IXrPqiZHAz9x6sofxn8QXG+hjEBd3GH/
EyHj+h+SiEHE5sBQBes5LJQA+49MyXraQwCzcK+X15kgRYzEy3H1nsbhDSPXGEb2
mXrzKw/TQMXlP5LxqvDmTxMRJY7C/zsvnotE5aMmKA7MyW9wVwXqV54e8zz9ip2O
4iK6vGNpl63dhUDKd+0tmwwOfwrgCeTPJupvO40+h7a5+EbsRonQShrsSA43/BCK
O6bwvfEz4MbffE/3bvPNqp8ly4oJaPtWiFyaI7ESo4JkO7o62Rpc1j40trR7K66L
3xy6XoMl5SntJ+KKtnxjnEff27cEcvSrwC+lYr73EnTwerZP2gQXfxxocBcjD9dn
KzH3IQ20MV4Nq0YS/F02IJyrqPExl5IGAkHtZ253CdUGhCw2PPTZghn9DsfczaGv
wcg1zmoAm7LuyNErYmRU4KEkS/wwCO6JM/ZcWrW08+tuqDVZTIF49cp2JbZ8vM9O
zb03bXVmjQUTIM9sb9dpVznZRnbaYKdENT90CGQNrxK0V0OHVtAQsjFnPJEBhs4I
SxgMj0Cx+aqAZJDZvWf/x7zq4kSkH4ddFggyaGMyJXK4IEdlEAosKpg2BOdJcatk
fhD1lcxdk6teiq2pPiXXBUNf7owIi1qwO+7+hBd0e7sMWCQqFc/gN3xMFgTlQV6E
4VttD1KYFlGAXyOwdGJFwG5XwHkWCo5kAlJSKZnQUaq+gjHzi3Nl6p66vy62pKd/
hSfWOFRb7vzjbhMtwHzvDHIujZhdCMg2lnztlBGWo1162D57mNLE8oh2PTQvUtdH
3aR9GZ+3ASG504JBbKwu1PwnZV+4TTypUlgIcq43nzfdKVERNrkoWhntMryRwvy+
HQ132RjpXzVDV0RXD35cKKM7KM8o4eC0W+wzjbO2qZP/zESd3Fy+YtCcrWzpFodb
um+qZXXbxr82igTAoEtPFE87yoLtgPHDiKY67Qc2xQgI+1KXypILskpoXL/n30uc
cBz0v/rQE42Q4seF/K1yyNWIe3vJe29CgSGexPFR5vAi7i4sHWdJTuIGTbp9oWtH
R31XoKG5jL+ueETubxrucFI8nnXevcGlq7tIi5ZILkyF+gk9GOXq+RocXWjX8CIc
uL8f5v5lbuNNN7PODS5xHt4RLETQTqb/fa5VzBiGHrn4b3nau23rZpOpMyvUNJMk
Fii61Hoh5Yfb1UHRuAPWgvCWb5JPvl7o2UAi0FSMQWEKCX5g/7rvUPchi+JsJrIw
OteYQst5qRWniEYnREddmikKjKNeU1sG4OM3AKMi1X1MNS9gncegVtATPan9wlZo
VrKL65wQq0KpWq0ime4mdTu4RwO8KmHQpvKy5zROqfW0sLRU+2FPGwA3Hrzswhcy
p4wsK14i3XLsgEpk5HWypEad9At3k/WqRrMgp8i9+cX/6YQqfRqe4Q9XzBJEaL/U
7Ixktwv12ZwMAHEcgNXjjTv+pb1YI6V+EfSQxza/qbUEFd9GaGsQ9HKcznctKRer
zhjJZ+bS7wbVORnr7lleMwo/CeOAFTPvATZilkWn6HmrxlHUHSClACatXXvelt5B
W5/7drgox9qccpUQmxNccC/QhCTaF8ydUOAZwNZaL4z0yDr2sw4sBU7laTB6Y2Xq
y1kj6eVSela7qj4YYo11dlh+Pc8OcyFhu+cHt2tGSA0IU25czxI8eY6xLZEEUqrA
GjwoEVQ3U5WXd5VkX96FuUG4/32X6Vwv5Ydw2s0GdWjpt6cGrRB0K//yzRZ6Bu+H
6KG33wNwl/Ec8FFMYCR/kEQNqgO4i22v1s60leo/1t6luDvPVPOEWOSI3VYXTV1U
SCWTLgyn21r+pulvu9ClGAJv2bkC9lOqiEh47g7xVvtw5sB9IlUbHuqtdwLm9ktP
eDtivFVzbSdItmVirncodKTjG+GtKbIIZd6dGlBNhtofeDTct9BWs3JroWVXB8zV
N4Zoe+whp4S22J1/4fTt14ObNiYIQVKzBFj81RtQtKRc8IKCfSwy6EXJeUkfrX4w
CKWRHsByoyNMVI9yubmS4ia8RKdvrjRDdF9DteTMz16hSYmwZezreulqvnUQV4uG
jgs36+vn9i591SZhkg3u8PouaMN9hFR7E4tdjAqXe8EEC59+JaKIw11NPQwDRR6M
f3qjIYUdpQClxIvNXpCCdaatF76A6thtjtmkcdWkBObjZCZBC1JrVRcWSn974rFi
9ImzIoFMHdku+baYtXua8JerCk1WVZgIUSspwcmf+6hl1MpSJaldEOrdT9pw4G+W
aFpcpWva34Q7cuMrUn6Cr7jh5b7Ve6cPQS+V48ieiMYfcrvMjwPV4Y7SXs56xRGV
Vu/PeToLcfwreRZbwutDa/844SVoyYy0lWi6f4U/iNx2dKlnSSBayK3+EPfIK5zP
SfkLcQtZCpGSMwlS82dtAuCgsCuHQCmoBPV07+XhDabFzUI5umFjrZ6EuQ3gvMkn
cXgRFI37PbkpfFgOh3C5pUKkZNru9y0r1/4xGl/E1be9aKQqrNyT8g1fh/j2je/9
G/gga6XyPSU5lwHwvY5T7ZEYZXnkV0itt0pWNWe+FnTBmvTvzJ9sYeEUwF3oSVh4
1X5Vh25lJcIHUB8f3n5hilWpv9zX4vayrY6TrfAaTVTB+oaOAgqz+Fyk4L6aQCyh
JmGSuMN6piQljwCiFCdT6d4x4MHZXK7CrTiVO2Bu49lxAUnb/U5/rsi5JjhwlVQJ
HRUF8JG4D5mZZUAnr+dpYuaGaXncSczKCilqbk5Gc6o5pidjrHLbukX1xxvAO8BQ
M0kbyYmOoE3z/N97XCQc/6uZPRwQzPL3wdwQrShUsi8e0fJBwThG6IyBGk6AJjDj
rPPfpZcSEXUyTNGKejwAIUuVtpq4UWTJqUIbBzPJol8bpSKkLHvXjjHAxap13iT3
NKpWGBIflmCOEMIdHev2fIl5wSASTzmDfD5xidNaH4jvsDH8PvuRWGqpc8aC55U+
bZpJofFm7rohHbLtaj3eqWVN49CSpsoom4W6anP6dNd043CKtyn/ZyJxXi6hgpEp
WGauNOPqg2HTLPPNA9WffIrlvP+8h+WA+oZifKev3GhRRfCGyDcEM0DIqSybJmvx
0YSH4CYdxTL+/1ewFnciBnSTSGTPcIHliqYofz1kraEZx+F94akQ06nZQ+wySyFT
Sp9tCYlaRl7Xg8Ceqp3EiewZaTL7oleMcDlLsyP64L9o4P3oh0U3OAQhQVZfRyVB
MOpU6nS4I6x0LwNXpHW/wqWUzb82LtGfqpQmcDWTTDZGYQMSvQmV6ihnFEYWhnsB
hb/2699kLPBEog3y5FSKsLk+kmNLLqRAS8zOP646nos/fZvFUmpzv6f/GK4hsOUa
9BkoQ9N50xeOwchcaQMsFTDJx7rw61/vMpgXHjVD12mfR0ionlIzgjfcsomY+nTZ
ky1YTZ91+xJO+anAWMpYxcD90M+wsDKavoIAJkznf8DM6Zrczpxa9CzagOHglHQR
WlLMb+ofn1X1VvkhL5gw7QHgZlRVwrOR6pzdYKm+ODuTGMZKbrxmrcuccIolb1mh
g5iXH8Zf+9D3gPRCoyHcrWZBCMu4/fNHSJlpl8aforFvrxgXGSl1kWmtYjVIUNqz
J2m+n3U80zkR6d9MvnERh44lB8oNESW8MrFwOcpudL/KLATAyj5kVX3bdnCwE1qp
fwfMiiW/JTdHXqLY8ajX5iJyYCXJ/ujsiVoRHgWTycEVH9HIc2daM/zRwTFxUBY2
6zmmzjqtz1Im9xkeJzz9eucwcUGq/qPjOtPnLIHk8SwOB4pm4lOtBbq7em4Nm6MY
+LHUWI/AoFRLHIO3ucY+28g5vIP+82iUBUvtXXffVA3DbVnI0akaNARemZy16Nv7
W8i0+s5ZtnNCtJ4kAzvL9Fm0gZS4X3/Xj7kK/ZmKlIe8lriySGLYycL5yRw8Im/K
5u5xVJrOzYZRAcj3LkKmfvUpg0p0aQWggWWJm4uooX2mPiw9sc7DiSgdw7iXdfyO
dvTCklTQ/eACFjn6RNNo0Jqrg3xz0fPzWRiqMcujhKdBXpnH1Dgt5eavhM1My/ca
+WS9tAuxwSulplyKNFtIOKHvzuXDpvnVEHnrbU5dMqtLHdnV+ThH5Mkuwx6csdRE
OMKXNSre6CLjqHrRGmw3MiAw0eBkvGTDO9Css6ISQOP/DpJDScPdSrOG+RvlndHR
DTcqp6ai+oaC6vB+wqez+dhd+xKJkzH8D5iTQq2K4a8tNZnTpcb6n1EwVVrerAMs
TTTyi6QzDet+r/W/1tRBW+Y87SmITVqug/GrBGRoEcXSt87/WzpAflKJzuLU3a0q
086uSo52rch3yIhVNY7kZW9jj7kNq2RVJuq3DHsxVFiUl1QtLu45A95VK1j1gf7S
tJDh5AtnGLdOMwUKKieUM5Ln+C5q4ISaMSX9WtyXRiM7j7xu3tEQO+QxBk+4VEdu
2uM5RJdoQ28LPFNwQwJlWS6e6RbZ4TglwA+8c/igVtyvshtkZ1CVtPNtHk91fbI0
zOXkPEnLy21Pm8oNQ35S5EbFb4NFBVEwXWvNnzLSBv4rWTwi1d816M6ModNe4omy
FmjzNm1Wc/sjWLN+Lwdoj+fL7P2P428rG7wkYTPQJTfi7tYz64XcR3Fekn2JJFTw
mUCK4W/dFlq3P8+6zssnsbcrRbj/rO2sS+gvBpyHdtkMDcdFCPJ2deTIOUeOen1U
HMjTCZ3ekavCcSU6XetGvFvCQRXCuHV3pLekWklZY9y1V02PqqKoYPJH6zyxstYi
0OIfmCgDaP9EqJU1VIUMFtuBkn/iGsjlBTJkCm5CCHLZ4Eoizbf/b88g9NtroWtu
7GfP7YqeqJrbXtcFzl/V+yXmcNgpux1wyG0hFzBPdDKVw4j6yaH5UDpfpWRPHyl6
S/+D9wfePUMFYQMQOy3n1z7FctzAObaCUgpwlYXN/FCHK43EJ2GV5sPYvPSUOZ4n
j2i757sT+zT4YcceKZgWruqX0HeFGu6Lbml9tlfuYAGYVEhrrgkjzDogVUV+qZGd
9/Yv1NLJrIWYFy/F3Sx/6Ni+NMJHgWjAJQu3AabuSNxw80jApw54KnQzsXmoYuU6
dHJYgIecdL/IiIKMheqjFgK8lfIt+eFWTgnSMaGc7SPqS2LTUS0K3G0SXoc/9UlN
ekKisAIgrRnAYXYXIS2U0yu/4VlDq7aB/M8LDfOlbwQsNxDvCnNH6YPelXwM+1fT
qrSnZElDC3iVFaTsvM3NuuWwX+gCA+cO16XVWGmTnV1k6puNT9U//KNtpJbkFNCV
bt/KPDSNvHkNDb+Eg3MY3/JUCJTTKt/Y1IVMt5DXr2xc2R5PVSqJXBkaS49Od3oj
+NnNH9QZs1k3+D7KYOW6wGUtwDwZiP5NMpuRUKWcmORqfJwoHxflvSbz08gJawjx
FN5OQtNQALRw87I/LDor/1iKyGyJkMSpazuNyCQjw4OI7Mt+yCKkyg1OJlhVfT4Q
KNXsQ3YqsDextGVPaAPA3xAr1HO6ytWZUHr8SzvcWZVuhT02mBCCTnnqAqnA+NnW
e/NLdSORm7SC8iZY+iqpurIEaGVg+JNFH6FJdHVAxirqfc1EH8AnWZNlchUppD1B
Aj/9uLNczk943UUPf8dAo3f5J+Lc7BvQ7ZjPIH062vw+aLqbA3t3TgzEFbWS8Q9T
5FjXAQn8UdzyW2ACXoVfcqx2bebG9GD6Wo81HoSpIzpvLx2RCgnHvjQfCulmOcES
qj0dCSfNrHMuqKBd/8PFUw1skap89FBb5Txh0/Tt/ppGPasztNEcT9Hcsk+ERJF6
5IjEFC+N9MUGixlRrrW8Z5um0c1hUbfnXHotKwEfAkNWieXDCLaxby/g1jEndpFk
qCzG6+JpFXrOfSOtaXIQRRik++LB50l62FKRQO/NpsNH6K/l8vU5bWG9VnhTZxIL
Ti9rQiru4ChIANl8x0Ec+398ipOAdTCzJi0fbP2vhk5W1OzYuBSheRqwkL1X79/m
IHnvshRz+UCq2/P9B+sq3mYNBSzyYJE8YrBThpMauTl6fpBLReXTzZCeHmaE2KmL
AOLv435VACw1/LRu2ecYSBv26powFeal3ze1NzjgcU1BgcFdUHAXBs141xE0Ou53
FZgogFzMXaBVY53qhWwA+4IiR7hUDYmZCTDBY9I+w62gUfRJ5x6zub/VpFjgJAcl
LS+5iJKj7aSMIfi99IJOWRIv8zVg28vbmmGxMRfpOJsAbCSdlWEsyvw3KPod2AX/
NkIC8dGky5+eEN6jeGS2Nc7tWQ0gSSH7JwqSl3KbkS4xBMZvm+f8bkR5dYc3yXVQ
V/FTmgMB2ucloRZj2poXBkvnB8i/+MGKgPpUfOyrWEYDFMf1BM/1yatWHZO4yu7F
0C/FiGaXO1B8JhG1XymQG/VavpwcmrWP5UipVHRfxxRqzUhTszeEKdrvYPu1eRgT
uUdSWySslaLQbV6nLVP9M5g+rwaZbskvxVTxC68FTuwj9sk0+EysyQKSQMdTAQPY
atc0zBA/ZvWBYQFBjnCPEWvibbXvFaCThA1/wkTyDnI3LKD9rV1TF2qvzecqORC3
J/HB4sDZ66qZvLF9CwVrRpqNxz8ix8Znm5pP8e0lnprmXC8s3NULT66YPE3i5R7A
OsYLU3JIbbVBo72u+QQFDObHeK0d+u/shUfK1vE6/OXTCK4U053L/oqyuQei3kVX
8EVa8CxRfzY9w14/Ltb1tRgg0P7FZJxky/taIhR9qPxMaZYnu4XDkRc7TyPkPeeb
bDxpzjHecKxktGfR5oUTgbZy7wZTEusTZxk1tdAWzOo+VUomxWDmAXM5kHp9S0Dz
U3yBCKe6XZjyyJWdf5atujTJsev3k//MeG4hhCxkDaQgTx4AVWu81B/JXoG7z3Bw
5asMiVlOYrftqaRQvNYMcDqRpnsbUJkxFRrAddiAeBuDigBtHWJwV0XNBU2rnWni
ycz7lLLFzN4uk/eiS4SQRwnWnqxstCNzXzBnh+CJ8tAFMcuvxfe+Ay3V667hHSTY
jmgawvcJFuE1uBrBAAkxowAeuz+HvgJTxBE5KXa55Rair2vydKwcNmn77Ktk+rbw
Ufchhm0SQwReu//UzE+7CSL3V4pY0UMawmbhok87Ch//pkS0Imu1xRXfCsaMt8y5
WvsZ1wr8QF0Dv43bGTMCx6whprr0hljUk6L+GcICUiauYs4A7jJ/iA2ncKC44lth
mJK1s4pVZwlrXrwZTSp7qMsd2ODB+/ZAkWrEEoFxcSWU+eZ9MJ0WoYkS6246bNwm
bEQgxTSvjabub5hsNrUzdbqskMH01MjIlWsdgGnNCGUfL7VQlNwh7t0ruu8aKaoM
LY8jJ7un8RGkZgUCi0pNrf/bZnHjrMqfbTCWdlLVWh+h8zppBvyCngOvAguNxxFb
6vNBvv1A8oXK/5bzaOfaVDSbSOBND9lybpCNeHQFC0vuKTiBMuTvFqO8ZvdDQY/x
WYQYBMmvBQsGyH5VeIpk9AXX+oNNTWJOfSk4jUzmIMtjiohfmcz+Srecg6sywMcN
Rue00FLAEDqrQvMXG5xovIf2MTm4noFkdb3mn8a7nH5lMmRPJdt/q6JdoDwWvq06
E4ndi9n7tDjd9ePkimwYRN/vVCyXgwcyPJZjIRXrERUtjZ3dNs2jMJPz7sRxDryi
zhQiUJCTMaw/5JVmuO1xbB31m+MrtVys6LR1fGWvQO9mnzoB1q8hSB3iBtn/ssfP
tZEOdWZv9c1RS6o26cU0FtH7oWn5bsRwG9xUbSEYGZvtknhYjjPOHXOryvl5csEX
J385Hx/fBlw3sy6Z74THiXzn6LJI66OcT2VqNWgRR6xfyFz9f6Ewm5YcqaOpl7iR
JeR0dvfmcw7IU6zK9V3CkF+BdtNjEu58Bjjb8uMa5cMa3D5x4gd5oUMoIbSbIL/h
eNaY3FiZeEjVdLyM3TcZq2CtS3HdPPXZWScKI/FU+fNoTOW5OGwoUeqG/Obnvb1z
Qg7B+eCJbZXK+gvLAbDyphkOh7sbS2AipMHVsW1JnvVoSFsi7kxofkfHLWYl/Z8B
BFtIfGCPxrdmVIKEKzpKMgfGF38Otj5oaCWyhrewB/lFP/lmpa5wp+8CahtH5+KJ
YG0P1Spyu10hXpMVhgRSWaANVIS4JD9m33avq8EQolAbTGh9CfCK+1iGL3onkDGM
76ZdHrFt/xdTbKBi7hTqSwxmD5fhPz0RT3cGyhRUF2oOESGJ1IRIeDsY0gzjcquM
40Ss449IKhXkMDOPfgthoYT4bUchyFaIMGYzCmql/9vjn0TJrqPfwb6diR6h3HmC
kU2LBNEDzxf4xp/lN7R82EG/P/P6UJvc2vEuWlEWlCoOUihraNaUU6kszOLvuKF4
OJ5guFPVM++DjZ3w5QD25UV3t0DyzSSHZQNx1kOTqfEj3PLyaWPPtG6AJBGvlhUs
UFaNg0Wy8GgjEnnShU621QcyfAVkyytjGAZpURdGqZh9FresMXHvQ/O4aJcPkhpU
TKIO9QNdXlb6QSAGX1EHPtlcf41HHi+NutBizbFMR9pdHquYp5HhTmv9a4jRnoJr
Ft/rLEmjcGotkh4DMJSJnJ8nmQY3V/E3sOsU3SL85wjc1W2BSH/+V6kDec3wOBbN
SwXR2RNZYAbYsRQoPfrP27tvQ9tW1SKPAW91OEUcwpq36fOVCbYJ42n4yd/6OxXx
QDwy4FLtJuLAWN2Qbln3PmBNZ4ZwkpvVZbIqAI46+fMyD5qPNuYIFBgDqbygr1TF
vquwNQXKlTmduqaLFZbOA15Pi/z4myeDBQTG/TWWF1rPrnBdpVZKtUQ4TNJUBkF0
Cw6c3bbsCmW8kHT6tjYBMsuujaApJNwK22waLeI00pAtffLoSQIjMdTIljAi8947
tjCJbus+YM9UItuujwvCLkJmcPj7RxIbnp6KXnMbavqY1gGJ9KRo0evvf50LlAqZ
wdZRKznns3+P0cFO/L4aZMszXB69fRc6rGQhuHfUJD6SFOGr4L7QBAK08BjwVRZF
s2NAVnmQn9pk1cTJHgR87ZpSDZdMyNuO1DobzoNa64sNYzpilm4yNG16eyON1GMU
zBRAPeNscgxvmcxxWiKC1U6o6MSlUtZsrzfHszKBIi4COrBX0hVsx6l1F+jixB5C
dEWraMzB/QZG01vceILrzdvackq8QSRUqPWusbIcqG5stxKybtUU4HAKCFkm87VN
YQzMnifvdsXAwwIM7VYw5j5WIAzsCRrrc8YdLmicDijTVPWgzkZPNVBEKbrEKDEf
WlDLBvBN8MOO9PWPROT6Gpp2mChdzysjkiqEBB7Crs9uFrv+MOqPZDOtGRJdseH/
GDTbdAilMucJ0GF0cFkJw4sWonn8AJfIDok2ZfgjersYNlKb0V5xPmQgm0g2bZ/0
G3j5uTyY6c3W0BAZ8+TaCy1+VL46fwmzXHqF40nZsrWC29LMZ5k6KZppTxLOlYwO
I8JW55+pFzeFjLwIpzcuPurWiUu6yLtqFx6tfcUS4LRSoq66j02UWWDW6rVuIE2I
gIJn5q0Ry7+W9xF9oM1Pdan9e4/9lxYL2rEXWW/NtGFphnOjV6pEX4JbOh01C5sW
fHP5d6+HM0CvFDAeW+Em7jQoIkNS0awtA0uZiaZQFdcnwb9nmavtB4Zjt51mjEBi
iBkv2Q8YeFg+WdNndpI3PujODb/ZyxiId1kXorz8OgAJV9LjQ1H86c3immOqxDFb
O8RdmTlvU6q3OXKNBizUxQsmr3cSBQd8z3m1B5ptEoIhzyPZAeLt5/2viooQlgo/
yZBcD8SezoGFsT/hU2+uqcII83xWwBiz+y4OPsDLqNBsk63T9iwwdi7ZquBUzi2/
wAXrXOCk5aDkqfQ0t6lBc8kjJARMC3YoKTqm8rAT0rs166eDoT5TJKUvgkey6rJL
GMpn9tv42JBkAm3AFgW+4UVCyGPH9tjzF5Fe4OfHiR+hJYOrILMBWcSgkZcfuOW8
gJt4kOMxv3N9YH7+vA81+QWvulkpIMLU27VvWuE/BeL8bDeHJfIqNt1VHotXmCEg
pfGBBhDW8GEeSVqh1q4n2dAAcoak4bFs/FP2AC5ws1ZuU7miKJdooBfAQx2wVJ4S
HiMyYrH6gp7MwBkrL7obkGlP/TNDXyeH85yuXWSXwSfLihMFcTyGjo918qdU9BKc
kDcQiETde5DdxXVKodPQo284k52scSuMzS4W4I2BmcCQ7Dpxn21KHvUAurtUiMD7
ga/3lwvRyg4Bh4UaF8VsJYa7JYyF2yem4njBVe9n07aVx2DOyfGzGAvEyHPayvxf
9zdC8Mkjj7rMm8PPxAi95GbnzZhXHTs+dgk1Rd0r1gV4lgCpsd21YsI88QVrD7FM
mXAUoWly6ypZ+sEqEFi3YU16R9U/UpqgQpR0A2Qq7vKh9WjoWoK4N4go/XBcf61O
URQuBIxfODBZAzS7qc5cbQ8EW0NNjTZ5HNm29U17L9HPoHQqAigEH5RrXcpeeWRc
DTbOgR17KvwpBfWuxNRniBtZkjsF0w3DkqBcQ03bc9R1ZZAS1E/4sBc1/c/FnLaT
S+c89tnkJ9g03BHy7O+mo5+00ucxwtSG3ny6xaJm2nz0sSuXO7r+0DEqiJNXkBft
RjTlBpsj6vggZwuLnf4Q3PVRz8bKqR/lDyKm/72QJQQ+MMk75VxAtrW43LeVVNOv
rPkzm67U1IYxBskkpSK4fsAP8nDQNWkXrqdnUza8OLdO2R0YHG+d9qbMVa/Ki8wa
QOecY0AS84lvOTTElBnOP8RGpKJVwvBHrBZaVg0NLq5BOifNF2qNHMksqv1a9lgH
qdX95ZErMdl9sWHStXbwJNXushpVIHmGvxEGMnalOkj4kt+FQlEOnx2qRiAikzGM
6Ji5AePgnZR9FwB0ELc+LATnp8g4LOagIark16iexPXKzemtZY+ZOXjLghY8oE6K
BmFFSro4Cnn322yInbws0qq6fG2BqT60ey5tn0E/cnpSKUpBTT2zjnVC6pL8RA3u
Sm0IYOpv2u3fDsxH3ZoHKfu42Hjn5rKRUE1pROh58cxS4d1MxeX4x6n5QeNdiM4C
6W1wBrvuq2h78rL4YF3vJtxGf4GNU1d243rl+aITFEfSFzWg+/+4S38wFW8ZdhMq
6M4zsKIwAAGwBLBpKrkOyJcXiCQ/CTj2/4MCczq7BGibndHppZCUKpVGqZOqP5f/
K8mYHopPXewpwoG4xsOFjuwKXB12kWH/iv7z4ePa90lIjLrvwKrwoRsGnlIMsKqL
eHrIzlYTEYLKjnKWufEW15dJ+v5TaVgefVPXLi3a81n8qvr50uPyhee+xALTwdl8
wd2Hr7rNkJrOspBca0VNnntLhmBSlr6IKppwSSfcEGo901TAbt7663zPTS5oIQYr
ebXHZZ+d6VSlYjfzwAvZKNBdpbc5LdJuPjf4VHiconNusbiVihTd3d5Oq+MSh0Ji
lyUWN4OSdCHfDP/3PiOXshsmC6nbJy8hiHC4jzfaj50wmpOq+UmpoNF5HnnQWuyT
9ZtMxKldk4E4HIYxwiJOAAfyrksIULGFpV4T8NW/j9OXhspATcxoQKmd9uhVRjhH
/AVMSenEhta2GTGfPVf7lLtci90R/lZMgqdVvYquPZG1qgJX38YaYJ5taB/hUNpR
ZZ+l6EijdlmH8ERtQ4Sxt+HNNvcDtkeEUTbSQ6M5+nF9SWoAKK9MGnMvzEXZhUvX
gJ5VyEeEhkKkOUdLvq2rCkgAEvZ90Ix+Rgwukyb0TLJBweIiZYEaiCfjm+abW/i1
kamYSDcyf70BdL6HgGHc9FOWo4HYZwm531K+O5QTUwoXA6bscqHXATf8wzTdz/3M
C9NYwmZNeLPi4wWUCpH5DoABx0mImXE3J1gCCEKaFJincw98G9gAJAg00QPzXEOc
SfVrpaTB6uj6WLAOCismKE29yWLadUUGVUfS+pfqTcShtC6dpOo1v0kOJw+sVqGW
nqKppX8lYtc/ShVdo2sbgFv/ch/Tyek41JRQqyewDxei0VHS8QBRo7WGKNoZ6nwQ
2g/0P8yfnJj6r3n9hpVrSTpSY/15yAK81kvAkYuYvUakzGmc3JExNOIjIxh1LqLY
Vi+EBhHy3Bzv9OHeHLzp9MmlbV3+VD15cwx9imB4LVGW5mGbNVQuzH1D4FO0yjJy
PwXG5XNmBN5P5qUBnkpjWJc8VhnivrVgpN7N4me1pqINRq2+dGp/4xRaosVyfBDT
IvOYYE59h4VoF6HyqycSAi7JWmXgNRvrTAiSaSpsVK+86Du9/5LmPCE4NXt9PfjR
0vtoC+lp9knx8hNZiNrs7zxgG/+DfrOaWzXIA4+nJ+OLkUxpSMNmDb87EwXuP3gS
BbcgCt9B4d8BHzxED3yu/LIOAjQWVcV06Gaqx7w/V8NlEhVwfe5pA3f0VO/Qy4Bo
KxKvoUEbIQluD/JKvEaOrg6Vd9ND6fqpVHbESxBk4mh96FEBnzkRDArodK7wFX1A
sxsboXENOTggKSMbS91pqEhEBHtc4QrqM4GktRmwhyER7ytiLTRF4Mw2T5fiAWxd
iEAeIDhYP+sWtAjAHd53TjPLMDdX0+c4UAj7kkDS7RL0W1K5RER6bSwkoFt+RaMZ
qbzJXglWmzIW+4801HQtGzut7X8ESoGFu8C+spQFdt8li6pKeTdUym2BkIqK2wss
zSpqkJibj9M2OhCUkZ0/ikTi2Oglq1fdYyYePNhrvMEJ73tDcmQv64Fv4jkh44br
j5UTyINKeNN9nqaztfAKDxPTmTGWt7pDbtw6Y5LBwNb+dfAJ+Y39mhngArBqeNCf
g1fjzsNNIhX/YLHM5oDSAFDymP6Dx893U08KzPA7dT+SFbf6r+J0824prd+qmdGu
viVCC5OJQh4axqvo3MhBWpkty+ZqEa3+UjUtaKn8GSIobOm/X1tFJEYzaE9ZE7gp
Eq2bQBx34mhtg5x6M9G8icBtgLC+VSBc+937Rbt3oKrfW6Gb0c+HMXIipc7m9Sjy
iXDdyoC8GHGx3Q4shzGf6cpMcLyuhHMKi+kiTo8IgUczY8r1UMMTMSUd6KBkV2AY
2rK8JS2G41xsnoxml4yj3Kv6dmyyMgzWB2tz+ugKDZDCxBNU+aTkfOaeonegZIbK
z6RuetfPNDGTg0DrJJ1NhyUxwyNCfWrffwdCyNGCOkc5XWZtF1z/4V+tkP4Vor4L
p2PzFdd5LG/60Am3tTQTr992gEf4lMgPvAG9X9ktYYqUCw+Wyn1W0CCExF60hBBZ
bvDF8v0jdBII5DIOoBwFKa1eLEvkn3CQJxmzdLEXBGL0rr5OHXfa0lB+xpmCAZix
fMvnT+gMcqv27VsVmerzMY/0JVGtgSnJWAOZUm+MX6TGvvBPGyK5TH5zQ/uVbWyE
5beCjJRrWiMs/6xvy+jw+KtATXQ1Pa9FIWTWhCOpm1ldt6yBJU56lbsvBUWYNtA5
q9MP+1lFpZRzPY3R4xSbuC8MH/Dsk1p6LtLT+Ow6qBfBdLj3Kj7lnLa6TF47v7v5
OHjg/az2FaQWKacLNCOPMjM0QpS0zKU+tOcZhJgY5/xv3nQTSx/u++ivxkT+zZ62
9EUqjzNz49+0J4evVzTR1+UseUTs4fv1OSsJ+CRfsxlOPaENx9jdi7/rW/8O1cqi
EHvL72LsXiAycee6sMnIXIIjBYmP+9/OdumSqheuzAOp3wnLTlmk7/kzZeAY/k9K
wWt2TL67OPUqcYX5tavB0u3LP+vQz0A2FrBF3VmWf8ibOhPbwI8J8bE4A0sPwEAr
DQ6T5NzULEdr2487VJezajAzflH9khjMOt9+OVS08+dCRsLL83zNCwW9Oz2LrOEg
qZhJ+Ont2UNsxLyDbX9rNYhGEpuyn2Ckng5A2M3li9hUAjYarXi8k8p7KXaKjjOC
iYPazGZOayOcAK/eHAY7RgPP191rAGRFn540V+Xr9FUC9iigeN3I08J5AMDQjoXJ
5+ucKnjRGLeFTl57llf1KvvXHNaFvJpIFrcVd9lswTqSPiZenHn4E1LQaynhA0zL
kdJWY4UVTstfy9rDzsfZExmV+wzv6tcTTTsB35ae28z+hDjt+Iy3PojRATO90okU
JomzzxfIcLmk38rMcJu0pIvR2ixoDnAtMOvq6/y1KLVnjsiBQdIUr70d0J+Q3PNB
an0SSouKB1QN5t9WItIUpyS8e0NpLxDQ/0AYu51AEs2uFPURIb5fsKDXPUIJv7kh
0XJDNTTkz8zg8Vyfwx7GTAf7Xq9k57vsUx4fH+NnayzGEw10IrgAEOSlotnFbKSO
21gSjmb7X/AOieHH0M4K6xUmlXCHJeBTB6RLuH3KtOAq2e6J0NNoHTwnLqUj2vzB
cGwGIS+mB1hzLJTwiwDqHaOWcrihkbgtlBoeFoozC8sFSPMJQryA2h0Pawz0pUfo
u80zWUEmyLinX481t7MLfOUtAnwmazomi8WNhHMg+Yss4BiVIATwJMSlIwBxzzLV
tvvFkZbrtiHIG1VGdq/5EhZJar5Jo1dCYsuUSn+lDXR1VLhjWf0TwRmKr+fARfj3
jFQfee9WnXGwtSSIr9mQ6NenPH5znvWc760M+gNIXm0JuRDCwvAFDCv3rdM4sgjS
CKZ9pmprl5yEriUDz+D/33utOXCpJQ6Ifa4KC63qnTjcgbYEuJ1JkFGkBq0ZTfwC
IuFGtUo/+DJaicAMoGIBFMJqvQCosD+XBNnn4T855czzIZMg54HjvC3BIuHdEw/2
l2q1BgzB6YmB2vbNvxaj1r3bjyHDJ0wkWYwaX8cBKbCUVtvDQNwbHqeE8TMDPqnY
/FtBL5tcA8X44AiKnAoLibDDXK/MJVH24iyhPuwQ8Wi5LjSx7b8zPR9HnkZo1T6y
aHAKLFwEFfrpfQPZmdwHdMU8RKOL6JrsRB9ZZIddKxFzMlk8mtvKR/edSbExEyxz
xh5JRB0FvdIz4ahzF3ATXuudtAmnupSANPkaRWVYbII4fsZ5QqlWBMs1SLeUVnOz
X5Rl6Jot7HOtnYT2PCtV2h7B+4xqCAfb/Lhq/QYKe7vwscyqgVCM83xo0bMokfFL
f2XurhkPzSAEd3o9LlNjjvsnvQMeEYkndy+cKuslHTyUHQ3KStEZo2jPHlpxvYcu
RQE/dGQ79NLhF5+urf0XBimG4SYSxtI16RRGIzjmOHJ+L2EYB6l5Io8npXOqWOoM
FjPJsI4XqeTgA/bRzcXKbs2Ql+gzOdQJw14wd3sgEA5pHd/RsCDrwrdhA00pXGj6
uc+a19yPD27ESa9ArGHOhev7M84ciUmA/ynjsz2WW/KtFjQAcYuuABLrKNvDGnvJ
hj8LioAPFwVeG81/hjFCPCeNJSVFYEKcOxTYg+LmwdBIl6ufaKo+sBNXhaVSn/mG
e0T1GMdLYFMnecWQmj/EN6riQZKEsF1S0eeJcf9fvAirayjPHKOEBOhf9pGuHWQ+
j5cbtTYqNXv1WvsO6L8ZhKjzDyB8poZzC+pNuSZr81qAJMb+vbBcKyftiFM/Yi55
b+xQWBGxCeAZDHYjFgUKhpUdItlob6yJkR7O/GPNmYHyEcyeWCheeirBh/dV+t6K
v1h1sFMpHcARB6etppOesDrSkv2H0138oGKm1gJE9LLX3BMbgsp40qMzxFSnYBmQ
iHQOcTknCHsTaczyTpxazAhEpr9NfO4h7HMcao0vbNPcIPc8SFvENcE6gL2+Ju4U
uii4ZPjtt4R7L4BBV0btkUO1b/Fz9R7ssMMzSmnu7LelVmG2W6K78+Z4Q6PveuLm
eayvDFrgJDuQ8ExGG4ZMBO/Efw09VM/HQ1x6kn9XT+68IwiPDvcnhYdnawPrdLl1
tQTbcmKTxgIIWOoiEp2eLe/AnYuD0zjBAFWFrIovWdHUo6/+GuTT6nFbOW55DDpH
wHfhnPkpD701Xb6O2KBwxz2PKKwpX0Du3ZgiqYamY1hYm/nN1uJGgFJyFOMLXNq6
qwqPLrdvCpvaglGdLN9tzKKGOrrv+Q9Z7l4t/BdfWuXTbcM8DqMwRdxaqBOjeg1K
dPSHoXkIkwA6YZF3iO7F++aAtBSFsT9Y36eGctuOyMMGA76IUUkEGJHqv+qEItU+
h9/gSQmGK0p5fRcFGFtJUOFxeQl6og4TQuxqWi8eFR2z7/+hLPbXjag6CjYFNjZ7
nuUm+9fJbhgRFPsFDcnkStb1WIhq+YbBTVSVAaQeHcb7zW5Afa36Ob4luTilvrfF
zkWyLWS78cz4zrbDOmD0mGa6r8IzpbJ2qA6o18gG52cIH5DJmCCAAWcAsshNY0PD
Kx7Z8R+RcksXL+Msl6WB+E2Wg6j8GG6NV9vjiKS8yo/iy+UUBv6bp4jxvFEsONQH
0VtPBTtTBDG1Np2jxo9kXaabJJFPMQObpIYpZhy698g6a/8eQQX0tWp0m3F7KpZZ
6MfmwRYMixZqzycIsvto/NuJuuB0YE9XdalNPjMM/dy1xE8BPKmozs99+B8C5t2o
dTvu4E3bI499wTUuwvfpMUu6EEwAmD2mYzSpQLREf/1OaJXl9GvzAI8eiasrjR5g
nq+lDTKUk+q86j8+Sxf3DA1MpK1ca6FcxtJx6TBlV8nzj8UzvNb7xHZfDFulXjcG
hKHSS4207RMq+HL57kfEAlMXCZpvZylERhrWAQNZVFra0TfjfEJi5v4rYToqVsN/
yYzPB1vuJw0hQQ675wYRilce1XTT+iFKJwwE9g13iGGkd5ncUGG4F0JK0LSzS7E0
+7ilH26p/KBmylmVy08B6/jKwQ2dS4p4xwpmYvtOUsoVHKD2yjHylPRIrnOM0OFy
/vbQsmz3C31I1CAWd8W8+0wKaov9aybyzyZIOzVglg1EdIsAxDH+sM/P1r6iCBLu
uWo5H0GooADIYy/PAFGp/8e+I6sVEmNODzdFEJ3P/QRfFw1M4jox7g/765ubF+Zb
TqD/vbHSvKgxJWEM92szteJZGfgptzFpcz2Qz235msNMCGvOMLXy4OppNRVH48CA
PzKHoWdG3uoYsUkjA3+/a5i6aArkt1ncUAQuZhAoB3vRLWIFmUtBCwIPPIfe3C4Q
l9ipXbbWIH56q17suzbhIDbgQ3oRV766ri0WGZq5gsW7+yvQtPFG5G579p1ilL07
OJlICtjWj+6u/K+ySoYqDGS1T49VqAVntFxcG1ZhQR8RnwKaqcBeomCRjvve8YbA
PC8UEZXfYfc/C4qWCTJmmUFqBcJtCPSseeAdaQubkVTDydvcdhn7vXMIzsaCniEl
MDsgBYFuu9GaBG/Iz1SWQeD7+ndc1n1C6ROE3+a5VRtyNLvTpts0sNhSqG+4stVe
71nycRf0rLqshgFxMzXHNRkvwqnDO8cfHJgtIjmTHxEd3NybZaQO4EAQAwxvUWQh
Y5YzdFjL//7UymTcOODBX/P826oiY70s96Cqmye5CaeZ67q9f7Lz01td2AHg5a09
k/T/uasD2eUXQaBWN8PvsToXgf2GJPA9ksQCobtihOJl7s/4u0w0trJQ8VLTxWOT
7Kfk4yD794LjdOJR0bH0QK1qrZOgZ9f18+bN01KBvnUC1hhjXJaYkt3dci5JUric
WIkPXtIJiFtcEOvPp8awXyiFHRGPNsomfiwAUICQwl/kAV+lbt1qEZlOmnDvn21b
e4iNjYAH3kffpDJnTpKY7EoW1KFYgnHMrvrHnBqgczhUrXikcllqpbvznxsXenqP
+RULFLKjkE+jIKrlB+cGqLe+rQYg2VMlNA3mXZC93RZwJGn15kc2QT3CfsKwjutS
KMlQFrcLXUCIcp9wYpRycIAJho9LhIQoiwKTfMvHcN65BscxyYFSLomrQM/oOLkt
GkPP1glzR0hkNGWcJf5C8OQXRAlKCbjTag/3gZ+cywhx8N1wMrvPSbvtnnvHIXuw
wErYmh8Q9Wlm0pysvpHcv1FsK52UMpKbSNW4cY28xZ9YKI3+bu/wXkO+1xnMTU/j
xfRgTF4Im3TLDk2/8K9N5viRA/CovDWWGiVhYrDb6hspflP1zu1a2u7ROgKsFo0X
zik5lTOHI3j6qv8nyRzEq3WjJCobI7VTdf/pusQhrzg2NOMeMNAthG0WJ+5oF83a
xFqcR9KwMkO02wkccpK+N0hAw3cvB00S4L/lEg5SkH1BYsKEGqkRHM4wMglTgc0o
GBE/xaKLF4k+Ww/RQg+lWYSo9ccmqxt41VkrwvbGbhO/4NWEc4FJqV2GIRIIiv00
vWAUDlVybzr214Kq2iQRKrCCvBr+FVbPW9G36jKXn7wL3XTu1Wrh7CPGVGn1ggjR
OS58LLAFDfBBspxsdwr20bM+TkzERT2oKHY+2m78RMQCpVjgkpWMoeZ+/GYzHS+b
JtvJygPyojlpvEn4XxdTDJtIGvjI02vgrm6CpvMYT1m/P9gWbanYgfB2QMGuc3Ee
qmzXs/gybGoC3gUKUD8z1tPF1p+/noJyHyQhFPqzFvczaIxmOYS8O9wqJGrwmlIN
ZUQNpDUQR/vSlTPhMKFrILjEWifhkL/bVLETqK8pzRgSQpoL/XCgwBuPSzLwoJ2u
zds6L+TtRxESNpTOxqFvv/llHH8KpT5MyvSXcERGl/+spVNnnnBfljsJAkehKO7B
UPK7i7KdRuqP7lOHm9ZI6s35Fix9peMMbvOVtWeIpmKPFqGBBuCLLPFi++Uxz9ut
Q5urVw0/R8D10b4D0V5tR2fSZve0/0zKTxsqhiRvplcdPVg6kBDBJzPLePkz8TCU
eImUu1npiJ0muV7b8f8ZoXdDD7yjIeC+4MZnT0sr/mojJEA0Ruyh7FRKluC2LYcZ
GXgfUOduXrSbJmphZynad35MOl/R8Xpsm/FjI9rGpGxX1IpZX2ijT50WiXFGP5h7
fern/xK4L/tFlu5Wq2HriLJJ1pd9Uv9Sczb66jNJO7hkqKYnFesmr4d2rMUpAGQx
gs0v2xJUlMFTlJQWOYMhkfcxGtSte9hVuUTDIqzpSBwq+5WLspytP3IY1fSm2AiE
Tb+lvUdhDNMB+q8wYKi6HSUp6sdGVhyKfsDjsImmQ6Hgcor7+3Cy7EO5X2bvCctP
MaOOoSQzppF0QrO5T+tQqM3xabwXN5I9H1tpy3K9iIjw+W5YJkzPZfnQQfhQFPlo
aGETJ34NEVok/7k/JsqvF/bS0YY/LEt5PLxXk/vp/wc75hX8E6v64kVROUSHpivo
cMMBlTmfnbm0+zRApxMqaS7fxkaneN8TqhbZVaiFVjq7ZagohSH4WQUgGwzgssyw
LMRTram1dMY6C1JXWDS1WI2BkkuIR6+3ZK+XMXHDLjQ9wVbfSgCDmNYROSMBW6/F
vhFMlT+vCsXrXdb7ms9AWiVNSxRXVoxrlZrKU5h9er1FTkDIuI7azfi+oUHkhqCi
/x7Hv27OeW60U6iupqYgTKkzm/z3F/FDjqeskIiatazxRLcPampB/diiztteC5Aa
PBBZcrj8cR2bWqfKcr6Z3w7AoTesXFZHEifdn51TDN1X2PmHGtAaA3Q7uyEvctzr
ncsJy20Cz6pjc1d49RFPIx3xTkpdqOVLFiibKn1G7AQZV5WjD3Ltp2KvYtV0iV9g
0jnuHcPz/voObS391D2nsYNc5fLgf6Cgt6GOKuf4qqHx9ju8qQyefRKSx+IC7ub/
4rmPL8sC0uaEAH10GElo8EygoTQTFiwmzSJlLYuauagOmxtfMfa6KaBG+JJeCGzx
gpKOCPHKO1AK0t4Fpc4Sv3lcoOpXit3y5SDc/NIwD0NvljXH8bqO1qcelfQXTflH
WG7McQnGS0PQ8dMrnomwqe8te3zLOT48PeSD3KnJMNzX7gj1jV/SV6fiwM+vzE6M
awae6XKdIRUFNMiRCswVQs2nAfHwHwbevdV9VAdYPaL5Qai5NRjRWFoGQB7w1jes
RiPu8co6aSpH8rAD7U/kc930We0pN+kWfQLxtevLryC3p2VBEi8RvNGdOx4FbYAd
dzQJo7Hs+xsyTk8ad6oy9X00+/3/wNYf+D3C6mVce9mncyQDYun5TxXTFDUxmixC
uRw23zpX+6/HVj7E5Xp/sgr2SenwKpzBQhZWB9vlUw8rmROMfuyf7nKQSU5K0czj
vHMGrL07kQGBSPGA1gtQPcKde7BWtWETXx85Ebwova+SSznOGLyCs5/4S5Y1462S
q/Fy2PzFmk9jpCja7TrdTofGUhr54KfqVtN25dKSQfNdHEpzK27kQL7NFuRx4Z9S
mySI5paiqTU/K055rUxDAtw8S0dxWYazj/RP/uv/1dMbWKwAcO43MwWTua5Ho8OI
UdabLF9nAKQN/UD46QxvVDF23aG6a35xQ054Mt54aN/NOwwa9Smob1m+k70Q1dO8
j5xmQMV8w146G5WDxZAShGDn+5gWwFinbDUMbnMCjHTUAss/5UHI63shRZJuplMS
YPeKD7IrE1qVSngNQUxTxpPPo9pNS8r/ASf2FusOo5jVw1H7lAkeFI4H3KaaU0kq
lm9semJmk3gwnwRkRPIb7jhGrrUWNNw2hWKLgGcQu0m8A7pyMm2lHgyaf6HYxNov
3Dpg3pFVMY2UVZmQrbgtqf+xoF0yuGzPiLvGAW69DWXK/ph+WxLbp/+HTyDSOANS
6UMz/EIFvaEw0ojltFlWn0wQz1PMojE1ReqIAUl+qKjMInQg1Ut5xYSQwyPC41BZ
ywBAR/lmWiTTYQuaiMlsX8b03L54jQVJsRuZ+ZsVYhpljw1yTs7n3uISlm+82bB/
DK7sjHk1JXilfdIj3GFRcOYW8AHXEso0BQaYs7q4EJkNFHIQksiP/eUu9Bqx44X3
LqyGtnyQTRud6HRLBYux33PuW8KdtXEqsIH8fyXj+S78mgAZ1X9Xzm/d5zw5Y3KB
KdCvnoIEPvAH4GfWfyGThnlnPBi/cENUoGMN3OIlzdR5SgR++uF15P5RQzRlS0Po
guqBZRRHlney1s1HYxffEvBC0qIvkasq8NPA4gH7GCD1VMWCDLjqb03un7CD3q8F
R4/oa9V/H3mdZRlcyC+SZfEA/OXk9jjP6sJEWwMd2haVtJIc2Y2w0OVljm6dKD0W
TPeEz44hTY5sxyEbYRLBWdA400j5yTzZPH207nBNPBjHhtE7IS5LgKN5JSUWWR48
M2D49Wxj14AnRtyrV3VeS78V757Nh9d2gvp378G5VRws69c+jn+/ySJg39PhVWHi
7HkPW3B/YDK8yXVk3KKMZzAi4du93kYIBOkgLl+Jxb4RsVDnHat7UT17R/jbXmxW
wq90P1mAyLPLS6oms5vpEKfx/C/4JgwhaJoTu3FIyCwlFrBK3k2IGJW0SbVaUeNe
iUGdZRKp3Q2CIwvNUV4qx3SNz9tsoludS/X1/ZaGwBURsq286lGtzuy0S5O8IopF
BM7UmZBqPcqySvFY9U+9M9M5BBVRSOvQdjWKI8aTaNMkjiz6/LIZpa7hCOsWN0Ab
4VmSfvb356ctj1AtCyf7/yVptoqhWMd03o6GnOYLsPz5+2j0Om8a10GBs6YSkP7I
g62hUDRDM78plr8F9cXGcZzqMppDP6Q+cRfxcbvEZJWkJK7GGLHDPpKY0k0BANQd
5HxK8vqEWCQxmsq5Qt0ExB769cB217ncy2mETZFpQFpAwOapHsLllgBYaN3+LBXd
76+EDIWAE+yXZitx+mkzy6SNirnl1Q/Xmv0jANjLepVEo8fbV2xmfWdENw0X5syR
3VWw71g2QQpAchPMuldim59wuqif3R5xXJYbCLnl//JI4CAO37pQh6Ja6tvO8wXM
lszIaM5KoXLNwYupu8bYadRqB7WHxVXPXXNg1ebKZM9GFBShvkgoT1v0TGSOEaYK
6H0hZl371brhV6a70/izBJUfasulgjF5zVgMFatQBOTlzFSj0+AKVoPN2D0v3mJJ
0+7mWVIhn7O1ZF+/HufCLi1Sm5G5KZRfcCYKPnrW8xDxBpv2vKOUrA5XSz4XXHGP
4sRzxvhAP78y0Y5CPyTpxCrv8zqwB0ckoiL+1U78JKrvkiETNke1Sk40ulJRk4d7
0H0K3Fm8wTjp/d+kL6Zrp4DSsxzboc6IJLO0PaAOHuzOEIILoK2IxT5PPu+W87dY
z/rYyuZxrCCex0GekPFrA6fa5oi9/VguTxbdn9Ad+2joyZL8muxHXK7qTK6bvc26
3HMAyh9bAIOHQAvgzCB/ls+vzWYEmEgSHMrzhh8dU4I4znwAW8+1dxe72UfOHi5H
AVEY7NTBeSUHSnpsnC2hBGs6cVrxdVH+knoQJL1gh5N6ZCYF0bikL0n/aQNsCFF3
/TyI5rN1OzDa/YsyEr493+BAlfyb1lrjrz10rOFh/WXpYTl6wNnuKfxVDolCkVh4
/E9xNRlGiqusMbHkTchgJ2jdCtoUbdyxBpPkp9QYymsLDEZEeiLwrYYlCh8XtFyF
fNBh8+0w/kE1T7e31a93i2C9yap9yAqY/T3DXDQScAcit45fSdkcrnMegiBMomYC
GlKZStWFQw/C0mZJgaOm/OPcDtLzdNLutGp69oovpJeAAEXy4wvGmcMm+ynjDYZj
Tl/y6cuOSXAuM0HndtBHACqbOZgJMZlQahEbp0AAdc+5ajWiEslaeYdZtIWZpAOd
dAnjcSfBksj77HEHU6UfoDzlBaMYA8Ot0Vt6TCV9/TqgGdMuL2ZzNQJKYSkCuV4M
ipYlBKe0aVZtz+H5DNCo/vaLdmBE/syxwnrNGep0s20JSGq6b4Lz0PdUMmm8mwH2
vRjs210NqTERkVboy9mqbF6q9xhpOwepv2TW/oixmrI30gzgBAAfj1+Px2l79DeB
WbxXEHutCfxBZ/vY7O3Rh4O6k3Bhki+mqrcF8SecRozrMuJnUOFelgreWzGx+Mad
uENTqRU2Kx62YKVrkp5pXBHRNgON8yYzCQtqm3UGC9NgZXVkPiQ0ITzPmuLcu7zG
94Yzgrvx0tsowkW178JgfgTC1eRuGuZrHTYLNw79MEfR4i5if+jDIc7DbfF9rfCU
dYoZfO5Rdp9w1gJyJo6tMSUyrUyTkQ8uo2vF3M109wras955oC+Uw98pebiBdjtL
mP6vAv09O71oGTPnPmJtRtWjNKHHYwb3JMh+4ltDV6Kz4Y80dR1e9+lVrCwGeJQB
QuktOrNsshkKRK7w/oYDYvxcZBD87QvwanVFKo4wcypzRhFHGnW0AIeJJ3cvyli6
L66LhchzTjxGEjcAyRFQQYDJq5ptKnBC7i56qJadK8X2t/FWAV6C7/YeOdNL9qHF
jfDYTXQKHXtbKos0AIGPXTi/Aatxukx3nApGhfPtxKkg6lyLvY6z0z1U9vviJuZ7
VZW+8NsTYHhUL6+WFLaaunuGzMiM0b0p3TB3YB6JGG7qthHJo+2YtcheDk/QKFl+
I7Z+6k+6gcaaUsXjYwjjC0iyNf0S/YUtStCZqqPq/ltu0F12Y1vrLnGVvx7qU8Oy
3jxu31xxeH70mr0IZPCDlP2gH7gYYNkIFFF2sYFFPHY3X0czgbMaUx5KzgF1nFQO
3RPUiM35SkOE7kcjhQkfwIChfkZa70OzNS+cVqlPp7FnVw2kO3MFRdUod9Hnha16
SOX+1Khw2NbdlHUd0AOB3IHGMGE61R/hU8VJyCHrzviUEcoqv1tAuBytzeeTEwT0
y3600vAoog82T3oiVOk40GWUCSLYIZdnhrZxV/FybGV+zUEUF11LxyD1VjLR/NCQ
qsRmJkQngWc/yXZW34iz62OmusZP03Big0W913H8r+HFeCWSd9Ha358qrfzXsRyQ
p95/0mjNJPHZoGchiFogBG1SBz5xue/1ijt7THdSkKJYtfwPHSbcMT+VLWh7UYk+
CvIPAZkuRx3AdJh18J5i+MBseoKigAXGeEkfZ/A6B5o1J7F0ssurQytH3bEX9Xb9
OhhCEu+d9Nc92P9b5lmNZIks0Y3jNv9UaQFh9y0jcDDiTx/Sdl+W8p3G1yTDw4Hw
iuYmMCeLo+rcDVn4Zz6nmCzhgzAuQ76vjIjP8UM6U4Ekx7bAfwupLjzjZAHCE6X2
ztR8bGOIYPBn4enkVgiAEPJ6wjO23PLWEOurFCuIOv95gUtHGBMHPXVaMbTUN7pW
LBMfO5tq3tEuFLyCVAp6yFfVaZTMgdJ8MIualYGinK9OOC7+LwChsD/zrC+ASDIU
jEKpIrhjx1d73YcOLQToRiftVwAJssysy3CRpL6VZPq8S8iffqhT4vFqFSNpTImE
D/kN+adn2EQs+sFqefNMR1GZ4WLg1ei0JWgdnHKHY8q/Q0uaNuu8d3m6J/zyK1ki
AZZd6J5nL4ets3kNlde6jv3VmyQzk3q8W1msIz2nxIsbPO5VdeM474qVAZ7VQf+j
7kp59t2ARVq4+OX2+sh/WskXQzjf1Sm0o7gnaPFNksIpb/ICXfkfhV9VArVbRQhQ
1/eQYyQxRYaOgv3S3zKQRtkjdDooNpd5C4wsXXcu+4+qB26qoVO8lpH3w9JIfByG
KNPDFeHQmeAjlOvJU0enaGqcfBBBMiXfA32mt830E3JI/6NS0xqcF9RnHuA1iij6
sWoDkNc8Ku2zp1Ind2OyF7k8K+NlE7N8NVPvDmeHnUL07wsF8yRwm3ConVP7J1GK
fQHbQM/y1XjiALXLmi0gr/b/n+jBrsNR6xE8RpRTCHASVvFliXsHoeFRGvqzOohg
9jpcrhXbGZonTwemANz1IyGZ3hCoJkWcskj/q6jLCQF0lIQVy589U28Ke+pkeCVq
d/4YhdKXIM6VcPJcNC58HKt7CrfzL64gzyqJ597LMVynV/Uqtz5Fn3tOLUkvlLR8
RDOzNIwwW+mwN4dNMUM/O66mpb2B4kyn5Frkol2rh9V74zWFHNbAAVbPgJYLIJar
zPN2bHxkmgzvVmutRRwh646ye0NGp7g0usIMGoKh29/JkuH9b341b8xtBsE7G3kk
FkCVtAUe0Z86jxSSwG7YjkkOhVcq//a1qbuFxKxi1w7/zAEWa8G7E4FwTGnk+BsC
KKl4J42cZDeRwZ2YCjz9kX9htLMQcT0Rd6cUUburDeg/BOu7bOu24RS9sByntPAB
0yNPlTJzF+NOrPk9PJnfCdZ/QL79mbYRQxhUIEGTIoHRO6yaH1qU/3Xv7l4cT5RL
aPNsWiyb1SYwNk/obrwj/uT/kla+ZLEN/SdsgK6t0wiLzVqecQhq3VtaCq/T1Nug
ry5ic/pAZrts2QJKoTunqR0OvPZrPv7J9tCPJWqu4u6RikmZvkjawBzeG4epDvwt
9//soy+p1UsYY7sIZ5o/4WRTu2arEoyrD5eEusT6kxamtgi4mFv3tm5Kasp/xank
Yg9cwAeSbSFcBJSvgaYSwPfY2+ht/YXzqsnR7cermc5MjIEHUqFRGXKrjLaNkkYQ
Ebct/6YRHKBIxDLJ0QyHnAHtRUhDwCbSKA7LK6cjDFhCQgMKsqUaGRI1GT6MI2qR
aXNt9o1Ff354yELRRw+kwvQ1jwhwWylKhCai3yGFZrjjUwFtOPmSq8VrR5pJXhP2
I8ZAJ8Hh+oV14yK60nEInM/QNYAoKRYU2PxO6i//+QgFuxyBv3xkUNjCjMk/q3cA
kUwsjvvuzEm8Nz96U7OhEqQZq4HCpZg8R/bLcIfJcxS7X2RVH1gC1sEEktp2xXbY
3wdbJFN2Oh77ElNmc++19GLqXGK/6gOQA7Ar1W2LvD2nlzz/ezLn0+dLVyIWNk3l
2WJ92RR1jsx28p3wGF1pxwjzaQJTg2Y3UsxJjn2V+qnXtxv5U5sDLB2Ft7DU8GAn
02T9udi3SQsp63x62ucVJOqeqgRg10B6+4hyZy7uIGN6MvBy0HVI14bV2+Mbgp83
L7O7QgL3QLZBgBGIkG/w5uMiS6A72a3CDKy5fSC9ufaNJ3iHk8D0wt8SerXzCo8C
RNzdelsNFillBXeZtVomTZZ+58JG3vzE5QG0s63oPnbLzogQcOOmr4gTRKUvzvYF
mf8gVPe6jObJKLb5QE5LT1NI5eJMLeOpXlCNRvpLa5xRlu9DrItLsUdVBCCEJwUf
hwVYY13B0WWqHh7cukZJ5Acf/s/bs90V03EaXRo1gt8YoPQZwYMOBAPbGKZkUIs9
k8ZrjHDedOdfNheNBBlHwuHkFwRxwbTcOzyxSxiMAYjdKDQ34m2Wdve7TNhi3/UC
vPoTcL3a3Jgec51TKwK2nj7yHrI3nt1CGRjlhSag8kfi92OFGvjOTge1BLlChJyJ
guAxSndJfiJCvbT5uw3eIzgfMDf1qJuHOI7VUwg7UsgsxVSxTPd4sLQaVzUtWwlB
paiE3UERCYm1WYMQ5PwZYboeBhzF5tyGx5BXoWP4Bo7hoRa/KMftRuyaa1cWhYPR
3ikrNWE/L6OLFsOff27cskwJ5Hii0wJhqiniWaA65z+MAt4N6mIIV2PmDpb/ghEj
/UWQvQNFBrRzRDWX9Lrh76ehmFkAXqsoeE/qvXAIeQyYKBGd4pKCq3QEDM407xh1
08GER9t1DApw/qfvB/xMw+ax1LoFPuPg1MyWGaP7sswkXyZPl4T/3z7PjQsa30h6
fI6xVBg1hjnjXNJxqrirMP2mzkcOxJEkBnhJ3vEYmd8eHHkLD5m1E+Vy/ImuEGAj
ddGY4GRWR/DSjh7hASgQ9e8Fod3ym9fnFSmxzX7S+g0vlsryBv4XR7juhpONKJPR
A5cW39fu7o60tizWVDIVTWhPoDXGkf6D67lEdgKjf9Uoi6AaZDJuvpGR7nF7Vc65
Q5rdckNSJRO1+7lyX1fQc3o6/9LRDVZdnNE7dcSiJ80oGxAR1gxjMv3eING4JuuP
HEk0inuR2xw4LdUy1W/KAR23kkYkZcb9+lFzC90dNoDL96Iiuaq65VzAQDrd2pFl
rIoSJb9ftN9Dokbz7NEJY9yRyDbZZMBLYjujZFBf3144VLGwASjFGXQQXhbUNOyQ
7eZ5QD8PM+FKhf0WMYwV/1VzKMdNPtX0IZoyOS9BJoMTtm3lcy4gElxArHgmUa0r
nJoyt0m9FxrVFxxj5N6ktLXCiDMJ5XlvW0kmySH1LZoLcsCHl+rUrvlAIVvxP2/p
uJgJjYgFIX+waL7QHFjaFWUK5Z/GEmRa69NoBNOI2qhhtcO0BfPcJXhwb3bndYMt
hco0pEAiPGRInSHHymgEXLPU6qrMglhmWO1fsHgrUz321ghLB3btmrM7aXd5ck0x
ShZoqKG5KHTporYoGNx22XaRrk6GhSpFNAEuPSBjyPYkQ88qnSiGwmm+DnauaoUV
iVOJK5yQrFUhJDPQQLFQeziEx7VNjAsb0+xDGQSrJFo6R5EZBpXZ7NcbMOGB7Uu+
RgFl2rUY3mOTcCRzDKCMG0zd4g+OMC4z+r0nI0h1rfovj4nkIqaBGJR1TSfHfZD/
2tKgE2cemoty/9XXgCXGRyB4PJkHd52ggroDPH/JpsZIM5w+2nNDDfWJry2XCman
P9cAV4jqZXXYa9Qxz/F0zkllLyCunK0pZ7pH5hEo6BWBtPyF7RC8h51SHyMzx1f5
NC0xwhhszbvePGWTYeOLnNzQfsiQS+m8I2Gzoe29xYoHG3/a1EPlJumg+4AKJQsP
AU9eDJTv64cK/2A2hn6RiNicXGxmXWHqJts70WT65z5zkixBQrdOpnMXiL1qpnB9
WAOkgPUGzRzhj952px4HY9BoBxGC00iPQVmuNt5sYqLp1APtHYd1TO16h5icDcAk
Dy7v6UgyJ75b8wfZ9X3RnW1RzUG3ofzxZjeffXXZYTFaVannwR6c9b5nXGwGDq1c
vrd0Htu/3x1gRJW3oyxmOJ5eBKgK/7pdZc2gQD1g/iMRbQmiJkVGSpBHu0FiUNEp
73N+DQhhqSmCPX+qOPbhvEOSmc/x5dC7y7K+ieKoRBuNxlur80X5wnH8yJ50q1vq
Hbi837y6Zg6zh73jWCjsCo1gRwjUSCT6X8t2Cad+2WFbCwqxJfFG2W927CgqGfDs
s6W84IrtQ6+MHGmRJNYt1zJ9vjb5cBdeZpKjR9tNHej9Ya+YIeI/F7sXO0I+9AYt
wc/hSg4AMYs7ANGoEVmLIl4XCeYxK++RsXEDxdosaE3RpRl13bUDkU/nuk1hODFW
gFR2K1sAo1A1dv06pnvCXXX07/R7hkCSl07Q6L8QymIR88tNPzJlNT5TtOnhWOk8
yx3TKRPulRDK3b/g++npNHwDiGmqi1c8wg/6QldSxQ02pD6EtOg4hqPXJVgIV/W1
lHaLHudyiFN+dxFVmxwHqkUzUwzk7DxUlp3Jil0A2/Mxl/BttU4VSAd45vnUbnfN
ubvfzcZOo6/tJkIDQnAV95+PhoMT5fS43qMj8Tm9MnBZQo77xFfe6o/4havSKgHE
rOuyai4lMsVOkoh55thhO4wS5FA+rwTILgyN+VDMNUtoFZ2S5BrZqllk42N+3G0/
15rdqP7U63i3zLCyDlCJ0e5nWayjAwaw4x0+EJ3Lamojy79GZikk0UEnUSzEL5sG
rBmpMklreWK3VSDz/I6X3m5KMRYisTL92CPDB11MukFDp5LNcOuejT1HNV4CkNLk
lTV+pgeqGOYBqZ0wSvCbFgaCW1loPYBbh6d9XZHYE6FhiOsK/djv5laNQS4VX9FW
lWxfyqlXL2DkWXSpeVQhspKAvWp8ODBPkfIrcyWdQCS/UuWUWBLaou/l+XEW7dtW
WxH41foZQGTc0nNtT+pTshNz6g36GZsdYd9xkpx7b0t37ZQbfgJOd8MiGmFBJDqi
4lgtUXvMq2Jws4Qvuq3nDaAS9IV9ZPODlx56EzjQuqx0/Qn3wmxb9MAsz0HUg8l4
gJm6ZlJ04HI++X65mq3U+WAypgKLnZdh+9QSJRCyeQ0viBadh99tcT8D7VWJ36os
37PjbKF62OmUSI06XHmmFM32rwov0utX8j3qvMG3qPXibRoHJvl2jT/KHdU2vD0N
E3Ydw3Hltl1eSulFWXeXaODHCbLtvHk65cOn4tjrlPE6h4Y0KKXlWj0P6G03dN0O
eFpn4lCSq8lNKPbfP9znZj5lPFBRKt7o86EAZB3Mnn6PsuNHxYnWe2EJQdJJKEjb
umVLCX7msrcDRM2S3XnvxthpBI89qf9+GA/Y10GhlfHtl9fLZ1o+AQGSHhpiy+eb
tJC7XrsVmcH3ib23EWUljFdAS8YTpn9sNeCtU6BmVGRenGIDCWwyznEismNAaWbR
Uu3f1adTtFGbD02/ulbhDPr2uyK9yOdiYQ77c6qwJtRXfZvl9NAjBPh3rZL6laxT
e6xIg94DIszZA2rrW0pFJPDjEdtepRVP65CElT0FOzINAf9iAS7aGda3BOlmcobY
lGoN5aXgEjrYoPce+bZQxGzOoot89HYHFdWpbph4kgxD1tuevSeyL5sXqYZqPejA
xkJfjHILYRkmv5KEtBpc4RSpxtg4CIZqhrsj8hB8q6zSNObG+N5xya8nAt7Veq6G
RZYAfYL0oCOSyzEwj/IPQaoDP4GtxMGbiMW8DI1g9D/Rz8arnU6ti+Qh16TC3OZU
dZERWiFAnQaX13ao3u2KnyhPjkdmTsajQXJJ26ZcWl42g4SLAYNKNSCiEDlWRKBQ
JawZmRr3j26jN71KmgBkH2Jvm+Pfj05ge43ZaTn0Wh7IcKtwIF+rsDomeQnTpMCR
yaWhCUu3O7QFc3vds47gObrbJpg7KkRKoNa/v5hvlweSzkK9NQFkl/xRGhEqEC2H
tfynHWoIKOWHFKsLP9EeeZjOP8t6VslmTxagF+UMcCVLLuZtA57uOudk9oRLb79W
FAJrkPSSGcniw1PzZC/yQFdcSdcypCzYrAmWUMm9Arw6/WTLuYmbn2ZTK435uXIL
4Z12TevrXvhSEilRP6icIvG+J3ztzcfWY8/5knKRdvldjE7noW6dLPOqHKbsLaav
1vihHCvV8ZJrrGeB2VmimJ1mWuFuK56yXwJ426SewrPKwycKLoq14Q6SSrAKqagf
X5KaNN+E1V5b32fm2+U3eAbDf9EOHx6QP6N0S1h36Net56iyiKMkzgOTOOhxJK4G
nGelPcf2NVtHwgwxfL4Rht5gEyDMBGTXBtCQ2DMlbjg+gwGiZBZKPTBLv0gvWT7m
4p8KttTSHfy65K9wsPeXavyec9PclwKvKlIu+4i3+XQwL74udmd+OEcwpUhPVukF
Gjm5m09MOfK3C+qmtw47999eEkh4t4z/gzny9Anwzc0in5OgTY5P1EfPVcbn9GcZ
r5Cm+pOg8Mi7NEQlo5RoZaE6yKsOBLiuc/1PZDyp8fw1+1Z2KiTp617zdSp0ksA2
/X66ZdDkJrKJWvlq922Uxw2z15QJRrN/NQGzNJRb+T3cpNcZUL6ko8N1TAZHkLyB
WoKEwN2Oui75z26RZS17BhH4c6tOB45IhKrt6k8AaEZbeaR8TXxFqh+wt9TaQLPd
cgDgSXi+pR8Zf5mmh0lmBQuWGKBDNQ9vmKkqsYlSMgUQFxIb9qaQrAdHZ/PWFuhn
oGLguEP9X1E68y7gwmTDb87v1R6K5u34rIWwu3atK00ojdkYcjfcqSWw/Xg67STn
2csKYFUXF9vQINQu7X/2VKoSYCuOl5pG6P96IH0Akr79ZsRPeWIa9QgGtlVEP/Ch
B6fign6cuUGpNvasK7YXmty8CtndjfB2oVZzVk2qCr/Kmu2JUO8UiasiBOB4gmrw
iyAiEQKIslwEpkr2I/5hI5N2cbg1ihyXhCjBtCikVkXak7ydAcwhfMXBx3AatqVF
Pdo3v/J+QfvN26nHQP/kfd0ndnpFDSBoG7O2R75h5B/5CwAqwzH1E2d0HSTK9ENH
ubUEPzrbR4coJTiyY00WU7KMFGrf2L8m7FRz3gmk5qV9lGDqvn9G+mwfdJn4R0/c
zNE1BL2iM6jTS1z6/ElVXKY5WJan5ksKu1FbCkUprkVAc/BZoeb2XowiKQaqAwgw
y3kH6Zt0/EYpxW10z5LoOwUK+N73kDxh7H9K2BvCLWYlTeHM3WSmJjDghzWtYzgp
UHZCPdX9HQw7ZsCg4xhfhE4IO9LU/JdamjJe1NFV5PNtJd3YpV5bP55NEr/bAw95
9nusez0CDot/AymTwxE2ysZsMg26nOh9ov0n8xD2YBXpc+k5RzNCsYF5pX38u029
xCDXDxnANFnNGOp7209za4+/wKoonb2i0/RIX89qUO3cmy3bigGIqaCuRWYLTOTF
WUOr3qSrndq/5GBZnFKIVyErxkpJcBly1QQaaES3jtBPyqtC51Q4bAfpiomI78M7
ABr8dNXwSJmKSSzbWFylIArUJ5anSgCAagdT7YYnkr/FzfN97QO6QjtdFKnozP6T
G2GcGW80gxdehSSExvXqjerPH+kqXLoTZFJtzPPz7Q9FPJqAtsp2EmAHcfG8fMKV
AhY44q2QIAfR+y22dqhhMwI3oatTiU8sSJKGX9xLj3ZOI3EtSx6XGHxTDwajH24f
4z5w3srPR/k/1b/g9F7XbaN4mEYzSdPc+085mdfqHIELrSFbqJtGdzV8yzT12zh5
OwJ6eXlpNPv8QNviHc39LEVPs5oLBMMkqhUZZDTqwUEgTckNVTrFivfUQwe+UiNr
M4zNdmLJQDQ84yI90bVqQF412klXH14HEs7ntYEPlhTePruUDVxf899lXQvOBBUw
LP6/zlzVXDzCM2RuOlEBDMbH6hGJnyhrIgmUFrsuJvzloM8vQ5ciTwFdwN1327Tf
f9Gb6DmZrWG/FO1ZhiMTtDRb6Y/J1WP+oMJ1NI2HuDeeXsuIlqK6qa92XFb52N5f
4VyKfWuezc56xePFGlaIqBb+7agdb5TK7V3Vjon1bqzGLNe90/0Ahb2YK90fzvkR
8YtUF4FhoDKoryO7pEYmRUHIW6H7Sl7017ooJy8y5O7+w74ghMZPx0F3PU2//nCh
Sg5V4hRAWK1wP86Oe3Pnjpvvflk0Bi7PRLDXGQu1E7UqyPqgk55jVHPwGC1rfQQc
V7Li7QHdY3dApvcTMLMovcoiDq6pV6gn0vOL0+iVMuqYyRjGu7UkbDvaMZW72UDC
6SQUGA5mFstlQBpJA7ZSHdzf6tbxolIuhkacJKkwsdm1h660qBxv8EQv0flDMqIX
bcwM7pjSaAKVvfNeGsjCmQccPVY3JVIplvidOr9sC/RLxS+4lxeuJsUHkgTr88UD
eaCs1TVmTqos9SIU2+9JnQEtIQoajOGz2NNXBRQL6WcsLTFIrrnKjAJ+1bVocXKL
m4n6sbpA/BgSjuRvLbzBplGDXWMMQCvQhh5wum5R3AJeZBN/vcNstrQtwx20ayel
j5i/zre9S6o2QxbpIZY6cD+S0Ydr6Ewq0C8TJybgc467T0KJSlDLr7Am4CnbhMpr
KWI715Hu5KdtDH+fYjht3f+k/vjRJw/PD/DXKbCKsnq2cGBYDT3/6QSEgzU3Qnyk
U9Vx4PH+gOS+iRyqNQ8aPraXIOic58fomy7ioe8oJ/MxQ10o++/fBzt8oQQsRsKs
UmK7vkA/hzDHObRpVC7x6AwvxGy1MGS8vBKmf9ougPFVn/qgfcQUe84UEek+HDPS
nan6TngaN7olfhrbJhlU/jgydvklVUQZBvuRDFFQUzAcF9lIw6OqjV95qWqOzAmR
3iwoaRqSgGSSjpxlMjSm4+N6rRTQbjLlWyfGNo1fVLLO1dOexG7dBwVNRQggOtR1
kdHTbaWIXPgicASjiv/D4FFn4BKloy4bMlBw8DOlBmYcJKcWC/C9BU5TJVK4x7AV
rlVyaf+E+Wi+n7MH8gT0SfrQc/up6j/DVB9fIih2fEF2tMQ6WLJtpLpvAh9wNKGg
FdrsMuyLrfp59HDPg3r7hUcF0cZClmGJyEDdQ7+/79UdA1+RskfGuf2yFgJINdTl
yfryWb1bkE8R2N4L07VGLy08cp31iKzmwEV+4a8WpcrjHBPm4UUoqqqV5FYF2XJ1
bHIX3WrCrhRpe5H9zLanlM0sYRufo2cjKBCUQedWuY7g6Li0esit4PMEn/bN2cqf
dDmfGLEs+HHTxvfuDWy/A67BepJLtKEGtzBFkhRgKbYlSurtYbPMxTWvTzeI2ACb
q8I9MU048zOO4r6Z/l43ozErKrpMU+yBW+7Mv4s1AiAzOs28flugUAWa0Q43takP
z1ne+8ruA/Z8zLbdOiSxiM+jvS/SQVUlbA3PqT2XxFu2E/4U8GwtS9ECnI2bRUAk
kywZ93GBZKZ1hFzUPgFpzXmPp6zmy8l4FjT8qLo8NkfRrtg9zPvVOo6pd2Fbr2sO
Mk65JlsQ5nttulth7b9hSW4zQz1Ou7OJjZE7yXZDaFmK2L+e7y0bgdqL/Fe65/v8
V2NQKsyGqW/9y+qhRwIMzHJfpZuksv93qGCwPSnHWZUx85weke8zrqZy3tmTQhoR
VLOFZR9su2TgtKFN49WDuT1WMXLgN+M1KgowStmZdZYEPMQT0iuzggZEkjh+rOJ6
48OneIIJ9l+W5NFVLAT2zGgUqXbncfgavXg6JeKcTs3wglzqAfas/AwHARQ2aGrb
+IFo24jBo1x5H524qM8hrAxazS/7r2h7E6ZisUOmvHHiib5yvK55yrkyr2pPOlZd
7PwkfgIhPUO77deh4QD20bV6X5uFb2y2zs/QZdSmP8y1PcnVgWY7CrrWJq70JXhb
1Ao+1cnu8GOLBAa0YmxIl8EZeogtUWx0FeVv4V1wyx1pRwZ55UUUDj5nwDBqFgGS
Rn0INsSnxe6BA7XK+MPbsu4o4VX4+oPh6Yg6GBRmV2ZpfuezqNt3Yi2nygPSG8BZ
iz+/q/eN+otjSBaDPBQnj6b8qJsbufR/ZOdCwac7Weao/wv4auNlWuqyr+lC+X0s
iKW7fQ6fz4QfDspQHTB0dxinAvHyT7MW1McUqkLVVMj3rQ0ssjDxBi+NyHd0s1zG
JOnUpR8OLCbqZ7uTomjyKGdXQebmqE4gT4G4G//mHNsEwNJyhe4+Z1Q3/11rDPXg
hJ7AfQ/VPS3uBPKqGKpx0XpBZIwtB1+F5BSiSQYdo2/lBfbefXxK8uqk0Mf1qc0u
IWIfMHLBXbzVXReMzhO8eBNcuqW3LzKQ+gZfgsDfYFVQAfVXX/s8weXNwfjNiyTF
flx6u2MJJQij7K2zWp7B3dbWboM8wDNtwkLUOYj2b1gwFYZWHlMtjc1t0hALl9iE
06DpHU0MGS3mrj1884QHOO8C/DLya9ZkLeHFJBpcLcBUqq0742/lq+ojUrtM3vuL
kXpo9ngHhlw8uYGDIUA98+vNbBmUoEsBGd/0PXGvJ0RSDhJnIcjTm406gIcrpYzx
NDGd4n9iCYCXIc75EHipRqRdfYBYBbn1rlz51ohIWt7ZHyQD2hnQYRm75E8uKMZQ
upydnf3bIuEd7Qm+4SdOH0VIOdTh5kqT8x7yQbM6q48TstXBdzjdRCLXum0UPMG1
t55JOLJDwPtatjNlkaH0AE8+LJK9XljhpFCH2/WPrM6eEYspZQ84x7CPxQHwy4Z4
xV7gvXthng4oGWah/4HtI/r7o5P/tSA8mr+DYnO/hau0//cp8jVYJi5KHsQyIQxC
IAKxsvaIlSTwmd3pmNkzI4x2LbppskLyZ1xO6wGYq9qi/6MbhrOnE/aB3XUoB45B
7NnclqGXbWK4tgMedXfYseDFk7i1/slI+sBMogZsPeQgPEMPPFr6tJ7WJkEnZoSp
/tfiptMlQ0nm2NqtimlkoA3UsGdv9ObsKs8/kccSBBf/BLXRE0Z2tGXGNoCqpTal
otUECkS30P/Xx27hzzUPb/wkF6xqX70WYxh0D7epVyFtofoIcJ/L62+Iyjb8c0nU
QUwUUplK24fw72e16jVFyAa2r9jeS3Dl4MIq+Tht+w4IC9S7oHqAQjIYi7DP8Ksz
7g1bgu4r18TGHLy9PuK/c29OMeajwuILFodVV8lr5ejaFsQFApG5d1asjhRSA5c0
nYW01D4gvoNvZfx8UvNH232BlvAhHanL/UiWFpO2cxEJGJ/JRT42INX+Qa4I1Srl
+uxvv4py+6yF9zvNjihbj5/AaELfQ8YR3Y69INhc26sniEa1QhzriR8V54uN73eC
VNDTX3TZR5GbAqRPY1oPCSYkrGYVgJwgQzRe255+sUn0W0WaeSmxSmhvRDsDhAtP
/o0z0JjXdgmhgjJ07Z7aAF9A9nHzDnhCtypRkmVqTArowxp8g0lmbaq75HREY+Zv
VZ1pLeME7eb6d2z99fOXD+O9cBCxR0a2EXUPN2801Fq6ykjKYysSYSeBhl38KysV
81wuFbwndj0mKCiIzjcdVUvmymrLpne8ajOoDC11ZW/GDaNUYPXCYyBqCTueUnb3
mfnSxsRDmc52aOLMTxGyraFlHwwlTroNpspVPeKaRXeSuonFVdRSvZS4IQ85WPVZ
SMSgvcZSqrhdDA77lM8j0exDKfGj/f7yWzRf3LDUBxR9TclOhEx+Xlh3nWhLFpcg
pjRFfokaXdjxQMxCcL2EU4zl6DKW+YqXKeLt0q0QqGgW2tESikUCSUEIqNnio46B
xHRotoOOAlHkW8uxKB3KBMgJnS8Kk0ckYjH+Wj0OiAKR8xXh/6kG+Si3G+qdqzV8
wPqbyEVY6fuSnjRjW9Z8fBWX/b2kgILGuGA3xuLBepB5xDoInp4417iqbk4tTfiR
U7yLJ8SK1rT+8F7Q7t9+2xYJUcBiHHlPT/RTs5q5GsfZsLxj5DL2nCCLK3wBdE6v
iDJ4XXcTmOIrEtwnQC4SyqKNbNnXF+wvMlEzWp/bAUFdttKMl5V3sfjv/jCCWYXX
a8rtSGfc9AVSQE1c8FY4mdsG+cW9ajeC5q4odD15Cvd4KSJTgR5HJUjA84SKqewq
ypA4j4pNrZJb1k+mzau5gvE6H6sA8/dC5Qhu0/uAIZfGEjzQJM2O2vPG7XXx+u5G
WegnF5kzz6EPUqCTUp9VLvlWDWflLX6HTqRlAveEDKyZFlA18qtiDfECFO8qT8Bw
CySwoaOaCGj48swmKiBHq9iXV73LcTbTJPiM1GijuvAaqNNgpJTRCH2frNiF8avY
4TLnp5PmGCAV5/A7PBVzaHCojoLpad4ZQM+BybNYR9nMMWcrsgTEtegMH6Br9HBD
rdRiPCbnjIPUXhUwshZHuFoikVU1H1vXA6T9R1lmjUkz4TclGCnNNnZ9LSzlLDhz
EY6l8YL7I3bWkvgZWvVeCpg/d2m0BaLH/kfTfEKzCS+aaUL13kMUFZgzxnwSQlMY
/7kzZgikNF1RU7O56t75tWPfU2Ay+M6Vz9U8kEDi2Xa7ICDbEJu7hQOFPmNfValG
wYBmr3FXrRrY8vHCWkxxSN1qQJEDPyfuz38GbXJTAYYsfcirPI4DWsl8nr164c/j
KeQB0yZWrnPVwcCyeFnWCp6iNo9Yo5tgQ8mTv1UuvBjrDvvhkzzGybeAClrTm+u2
0qu/k7A93gKiHq6tHQphD0rHfPM2zXo1ci2ChQIqOOSivvxrAhaKBtshW7M/2fHD
+9mC4TD5AWY64yReiD3bhA/Lfz/sQ495iAMfQEnb8tUGT/m1kSf6bCf23xYX2X6i
B1lrANNcxHmPfOaRJ8Xjr7JECjAsKEmySVpOI0HKkVsRmd/BXxCFzlZNQgT7W5mU
tdwrzhqVWJcdgspU8vwLydSPPy/zrg41NyoUU2yXbAb72KZ2I+F2u43xI1HxmwLi
bqi70Iw197PV3gjYwZdgJYrvFPiBLE1/yFR4lR/rDen1UPHeMpgBdynb59QkBmRX
hFBmg3Uhh8vslDDT6Ci+GOAdDN9QyTBTeXzmjIBVtOq3p08DDea+7cDEt0VRXxro
cAdS77F9JJ4EUpFN8TuRfYcGrjs1Unj0Eiz1qJanayyxAxoFrlHcc4XekptYVQMm
bGYZsgMUiHG4pyy5taVAwFkrdNXnF7rbueipn0HQ4HoI0aXqQ+32ZaUghGU+NnEB
edHK7shK61DrpWA0pDlaJsi6nLZIheGsT2RYA47O9FUcR4FdYnOtXHxbiFP05mAV
dzmmge/FIGARhdychZw39Ofn1RSYJ1TENX284Ntm2EQcOtoyd1ZpSZ1dwAB3cjaO
skwY9fsUq6ZrMb/yuDCqOycjm+d1+AyXZQZlkiztlCn8Yl41OGEVY7DqJRa+4hc7
ALqaROxm+WxSb4e3mR0DXYcf+ytvX3J/l0HPzdTgo2SeCDJpb1etIV11J2jAyO1f
0UGHyNheS7KzR2b+k+4e+AjD5uv+l2g3sF/gUnIYRBscwZVwxhhOEeU8E5AI20YI
V0U3H+135YSsCct3eYBuolgAcy7wx9YUxHYOHaeyqK5410ikG4kJKm44XXRAu0Mj
mFyD4/wZoXBcD8ktQW2/d5UfhTa5A5qFC9ucIf+slWoMvEb95fCgwwEby49IxRh5
9s48VQ5pp/ZbZ58S/GM5EApCLz64awztR8Dz+9SGd+q0QZSwqG8vcVwEtQXb7Nxk
6MoufTZGvqMUmfv2USxpxQpjnWpPhmMAIzU1C3INVHaFRkGMHLi/vhQ7oV/ei1Qm
UzlklqWqe7BrQfvrYmvbzLRTc1r5rtiPRR3cwpfeT/pEZVzKmcAak5xJsQ3a3DVk
nPnOaYNbME6YZY+gjQ6q8qJ/h7zjtP9qCpUBmeV7gglyEZwEG1Wa1HHCVSEJj2TE
AjzqOSryTuJebkfxhOvI/iCticekLvFfaGCCi54dSEIeOzU90N2sBpNkGySUxq2H
raBkP/q3jIFJ/jbLcL0tqvo6ijJ06cXQLftLE2GrgUSkhqiDepoPBL8pMiUZJsxK
9soplfxemAJTtg4rJqh7I4YVXGbJbHvDPexUot2IKKzPeWCb62o5fSkwc+49fdN5
6egte2y0INztVrMvf75fHzPcKhqq1Pg08Dfa49KVZ+uDJEarAcKZrqTIE9XfOzJ4
2A4OS0P9G5Yp3flWpfmGNzqe9+hZcVLDCfsss+FJiOc1MMWVjUvLXoBig771oouF
RNYMa3H0Ugid+HYE9971OAxYf7lQgg2XfaOtcx4gcFvFZ5cWXQjjGTBXN8cGpG+S
XhkLV42NqrbicaVDy+c2OGP+Nn0D8Ebpf40BRafCpCBHDHmNnpvjupk3mTaXmj9s
oB5XF5cw8JhTe3x+XomQ2H8k890RubrEihXAYORAeDRGEknNP5+ZazleRi78Ydhr
vHI2bYXa+N8AwwrrEb7GmHQZTP/C46qWPw8/wdDr82cTyI+EWYnCmyVE5mWBuLF/
Gav2snaSO97NMT8zmAWbplX0eDPo2n0kHcbVYOF26811YJ/T0fZ0kZFccjQynhe/
aiJZsAHbnoU6jXdYX3GDgc5pTr7zmAbY9vMIpej8NHI/EgGw5ukyLLf9r03ktNx0
tBxXKyZZygTUNwbxt6hj/m2bZ0oFEYoUUWXdQJGXflQ/frhnEY9Otok9eHkKzx60
LHjtxdCVXXIsYHGWqi8ZTpGDWIgRMda1Jvq+BdULoTXOy3OGASggdTjH9Tbd5IL1
cria0lvIyl4iKQfNb4qjxe3y+YDRFJh94j1ZlvUBCDWkoSTw1S3IiC8vBLIyqWTJ
GnPOBS6IaJFq2VJJUSiUgAU+tDoudPczwuJXSQ0WgC+lylaG+fc183oz88nswFgA
wr5vREhCYlcl68hc6wDFCOr+HOUY2SFQju0NU2Rh8FvrlSVXwEGrAHJVIwjpaTim
0yO/IMS/5BNjVW7OfSgtYCOnQw+xUsXTHFFzRK77NZf5MKT8Whx2wCBoJ0pDX6YA
m7HsBv445iUcaycd55SeQU72AhtkVZqIPQG6zdQtR6qeyumBxubwsq01tAXzejVm
9A4cC+ZGpZ7kXrV2c+IVSYgKmq/tFeHRwlk/sCnhoRVattbSQ65HuVfEE5md38PZ
XyPJDXhtPX04QABCDg+O2CmBZWBc5XwW7Iuym8DMwcfL2SBYvldUNzy1VSIloCXL
8PkDi1yfyN4JA65B36g7p5UURd85/jaRdHTW1f9ZMtQ0SviOMwWV/kgL77+dZHyI
ELkN+lK+tFSTsp2nYbxKlUlfJnNa4p+AdG7yeIuvf0sTzyOg6zw5zvTR2aBuz86u
MYrH7MmiLN+3Wm0ReH72fHzOQfxe7z/kNQjx69mVguBwQMmzlrPI6Wy+zxUjHkIb
G4VMrM+nWSzdr0TsTmDrtUJmL22c4AbkwZ5Ym030W8od3y2W2xmgL27VFeQxCEHg
P5ewscyg0A6dwKE1bdHpz+zG8H4LBx50arI/MZ3KLjsahl/zQYcsabqlQ+SaOGo0
b4qDJavCEhaHgVC8Yt3r0UQ3pXhs5pnz0eT+bG5iGabjHBO09d9tpqVBfOC9Odiw
Srgj26f1seSph80c812qvswdUHYuDlMO326yhHUDHB+RNBGrUN67NUnjN1PLXyrG
sdFZkFheYGMpDLkDPIy29ZA5dk4Eh4i1YeqeyyPG6sMAnWjJxGjmoCHqbWtHb5F5
9BTNDp1Fk8cHbvmdNBlZ75S1PlcIzR3C5rRxqlAFhbOW1FcevVmFe/ogP4JOTDwE
3AM/3HyqK2NPrEGjdMVNd9hrq5D0RHtE+Ser6t5kjAJ7DcBAymMGBgUEPeVz3RM/
0yUJEyLg5VJ3WBs9Iuxq82C206V68/n23HFmKe5uXhdfK9dV2bKNNLgUA6G0kLwR
wE7cceWvOC2pMx/OSFz8uFS7eyUBXFvhdm6VsoeWzS6boaqsDsn6fjaUdgDr6cIv
boEeYR7cknlFati1sGelXiSrZNe5b5WqBtD7TK0dt5f2g3/VNPNfyh2l0SsvVMDy
06oTaqzIH/H6U65s3VCEwFrkRX8zBr48jc5oeZOq7IjbfQV1TvmNobBNWpaB0G8O
pYIqClgn6TiVq3NztQTGiW6hYSDu+Be3J2f0jLnJnO4qSGXjA57UOcFSVDaIOwLI
uT/MNRYZE1ztgEEoDviTJLl+vbmqfZnqv9bHsw1Bm7JOYeyJGt0sY24N8AIQ4ezz
J62xl+tPtM1Xl+95twBJarvETiZIRhykmmj9MhQpBkESuLl3dbasVTRl1SChnKCC
yLFo11g6yvCc58PxCB0eVzEPc4mSmtCzMSzn05lllEl7YSaYhtp0tuSMbFBRkUJQ
FqVF3oaunsQTVrT8aiAxA4Gdc68he9XddqHDkQd07LowPICfLhtFg+NVY4h093g3
+sYofrvVBmasmkJg8wq4Q71e1PGll2ZGzZRqONFDAFTdaeudbZijFD0gHWjRuxZh
5aOUeKaBoYSv8HRPjugixtlw/4Fswrx2hzfKS+CRjtyPsOUW8BR2P/C86b9AApHY
H8TrSlGGlnlPEsSZSu8Jq5Ny+HVGccqDgVYoiGaEm3nXWxoMf5NOtWo2jJYYepIm
byJh2N2zG0Xfk5yAdYQTxnwDyq9tOoLpHNriFSUnu8dZSAgPRB6lpZPfqdc9U9ZF
ukX4qjf86WE6+XvAXUPvZaLoX0+vDTwBgAi0Xk4p4ET2VebA7uXsEu1b2zqcbPo9
75vR8MxEjkURw/uJir3iq5Nt5m0ZyFfpMYczvNuoStm0J2u+e4wBiw5khsnqgcFc
jjj5LiYjhcKEu3moSCVzrjO7hGR6W85W/sXipVevtVineTwSP7GyL7b5UzEkmRVJ
QkWU0DaNMN5sGlSGoV08ACJcRrh870U+tCOUwUml0QKKz4qUakp+Bzx8mVVwYftp
dpX+MmhLOka+Ch2ibSFwZJRH5p5UhCmvbyeo1u2S/BxMcXqFL/hrRd6IBF4nDqyb
DeOVrWTCdtWrOtXeks8IHD5++u6smpnd2Uc0tmzez/ldjMdgl1tQkYMmd3EjYzRG
I/SQTT8RqP4eG42r6C7tIXMGnyRcXKeRagXLucFQ7AuH06KRQ4USQg+JXZUXPBxT
G4bm7smIEXwmC2Q0ygTBxwjTWH4zerQjTt5MwtJDZtuHS5efPR5RvCVoLqX6uISV
8xu0eN4/DJmMIlfraJ3S4CtlFNc3Hz+Z5KNXEW5E9FmO2n/DZJGihRkeq+rDv55V
D46TnozGZzKqOHR/rSXxI63owLmBC8ryEVZJegbitA3oIgN9euSSQBgNAGooUmh9
i5F3NlijAnu/NKAiw6JzCMr0GnPShMKWwStf4XTHrrIU/TTC0HsjkHfQsczFe7y4
c1LJmjAhl2hoUkjDRtAGLRMBElZXIKknIWls3GeqcXdJ1VQIznx9/jtbElM7MerJ
k32L1lQIg/BdfxVPUR3Knw0VrMI/o42+K3Yxe1FFtxZ9K6oDaf0yovTwcNiPtUcN
U5fFeEi6peOZ9goQYrhpAk2b5VYO7LmBY1gWL6lkS7rWNsm8Hxi4S482ja2GcQP5
GvjhCGfFATXCB6pkapSmlNM6jQszh9sW0+/VuCGFUG9Zl0I7YeM9BwGV42KeKmDw
ubF3YrC//dABkfj0mK6toz58NYSKWCTrEw09YKgbfQ2FlfeZE8TVkKozevmAi5jW
xWMrkolXblTIuBVJNmZrz8ju5DMoVXsqE0V0YwUGDrkM0ILUvkcGwjBQcM3Yp2Lo
JU5sP1WQjkz0j5fECe9nbnFC9JqDsveX4agRFHaO90MlWuuYqwfeTLf/wEWvSPFB
s6k8CY1si5YgF6gHSRhE94dW6khZIZhfv/O6fjUIzh8WbEX+h/ceEX/lZ2gnbmHr
HjNsCPne2cg74GmT80BdwpXOGhXsxbrbN96Ste2wh3DI7vbjF25yZEEYVhEEycMu
pdre7wMXg1wuMt4xuqeST9w5CuMbyIBbpiK2sZhye48kYIEx1g1IQF3vgbBbA15Q
bQaEoYR45jqkrLsLpLN50g9FoyG1FzWVdiPE18a6M3kyIYOmkwch8HNScpvr6Axh
XN7FsAZMyInv1i7rJmREYJ4bIHKdPkRsIuuin8quIKNbnmMjGUBT9kKy6FE8Q5YY
F7b3hEUc32kb8rfNwuq5EMpk+ZwfRD9SMMZFNkXRbM5AXeS9TIpvlffiImwrAtxX
HQDXULD84bQdS+xJPjcW1uYurTxHI+HDdvSjC5Eo968CtB1+Yuhlc+xRi3bFO3/q
FHUylZTroiGrzDRAHVULxXdQ0wiFoLyGoAl4yeSXkRb6mGZbKBoAAWj+BicY8zVO
dyU/aBbuleV34Y6wPlgp4XCxxYG8v86Cx0eQVVn+Vi09YITZERVkCE8fpY2qVGL0
WKlNTdgfBCe+jfNOAIDfZSsU95/v839Py3JVI01d7UKH27/EC8owRayvnjXtkCM5
hTmn5YSpY/bhTiyV1vO+t9dyOJkpCIimWj6b6T9a5R5DU7VW6wPqxSOcGb/YBtw5
EOl08Y2uQOg7sqgbIbilwFz/1y4nCCw/hvhVWi3CKw0g5iWFdk1p/udXqqv66Avj
4yan+KzBK4VDQVjMdzJfolqUpXfqFRGQj4VAXi9T9+wW6pgCeteyG3UjzEi1Jqrp
zDBQvKoqwsMIIAnQlkLbJTb1UNlCqt0o5tohu5YCjsCUf98j1zpaVH9z6x/yBxPZ
8EpZyTJ0o9SInglaU3K0WT+0G7JQdWLI82SMUkiinEb+YpgDjYQpQiYIT0Rfo2du
4jLMqmvJirhs3Mtu58djJFEtQYDZMmJUKa+Rejom/tiXPwO4mLEYkrPtpUkZ3M8r
otTCzGyOfK9NdpjG+L15zTJxZVOsDldF1sJKC62pTxu4dKGXw8/O8Qjl7s7/KPbp
vX1A1GW1K2arDabKBg+QqZSfLqICyTYh1st6y0rC9zRqtHGxBzrNRGZZXI/tn3cs
n9cJcgy/RlXx5vtx8kF8mEVr6KlHQ5YZu9mZLPE8Ie0/CPwR+n/Q0CZXd56F6gQq
Q3bU0eS48iy+DjE039VVYD6iVAJjFDcfIpASSWFWxVVyZC6FQegWnHAzYwBHVpOC
tPWXpfElEm0/pR5LcEx0wVjl8MmajhfOXvfLyFK4+3/4yUIm7ODMbqoLjT7/9CRx
LRzVaqfe7HzGqU3hwIhvcfvEsauHnD2FdFGNDx0Q2vX10fW3UGQFeA4nvw9L9GAT
3ynPk2dpa7Sez0NIsdlWBqWVwz2/aa/MLdyyzA7xx3wvil33MDTTE0mw4p3Z+2HC
AhiRtH8CaSJl0gOAHA2z4cx4EDrBtKcmMuDeHhgWDhmuZT9TjwTrVPSvR+AFSO8e
nEhxdpX6dOWSAAFtne67DVpeawmlPX3d1mwiXBnqGvxSJ5OysaWc6epyop5HyYo/
xuy1o02+wg2tWZRHzei/F8lGBcD7pjVLLjwetdixiQSYM62EwO9bzEn6+kywIh4s
snOJrBcyGMZWIsFVj1q3Y/CFN+SSmXB8ZCvGCjso4CCIOelStGvpW1rwLen3FJod
8Mo+loblaN+5SQ2KLwh75JSJovPoVorZKkY89KuYMVT4JHMKEKnPBn/Xs7w7ok31
KnYX2LPGt8ftpTuXGww6jX7lR3n/Ga8stUwrLYGjFzNcwPXeSS+5FsY2J+cPMZOD
3DIcBO5Xdvg4JB+uPK9rcVMSEFqqxfTcTen0QWaowqNBOM5hh7INSEGztjpMqsyg
V5B5waMiaDomejslgoPcdF/xRd/eC2lawWvMAmPXiGVKjp6gIWtSc+KXxJ3kDsjr
8agf3FzWR5xKH8jZRh26PaIsFOxLW9qNX4tKSeg4sfMgPf8/kazYXFJn6eGpUEAG
KwIFlueiJ+ILPjTGG5uVQlcSNcyYdGaCHanpnD3Zg6cFW+wfLGMzq0kLq42DkuSg
fSlwswkU8+LTWLz4/ZZVFkMJQrtK6a64ryLBnNVlGxCe9ipy4BL6FQC5uLeouaYb
SyzaQCFyzrg5WHIUKODopharMy5ynIM7kEX6XCQXmIzQC2+KcObN6PtIdPzHzsrY
4XMlOHn8dVM+nDb+SCET4HdocKQ5wnPnUnix17TS44jqxn7mmlPBVP1W7Qs+Ah5y
kCd9DWz7tvleQe1FSSHDpibsEEMN1SqLP/UXWi28RqO3/qR6J8Jdo0ornhEUhHAR
RqL0mBMxqr4O4h0pxhEfitIoaV9Aon+X/xDzWCttpIiUrH7nsum4acavOsEqCYw6
cz1JF3jeNcmUG0eXrtGu4FOmllUF5LntdT1UF0zf/10T/A7zIDoSB92b8PVuVy93
Z6XdF4YTFdVk4Ykf6T8HCFn/WjfMJAYd5dHSRVEAJcYUfxBSRNH9j/bzOIs2XBHE
MveWWzEMmQl/Pwi9PC0IxpL3UVVVw4kpQUIh28aLL0dFmo0niIbRQQDT7HNG5bCl
DyHPXw1oMDAVaj1KTnyP7OMFp8BExO9lEnC6k0ELZ0Ol/9gq4zfsx4ioT+my3j6m
aS1961ejsDKNe3nnZ1sZ6QnO3MCA5TKvtHCTHvQEtRWzE4s2GTnRYra/Tf85cJMz
Rw8pJN+mXLasfQGgCnm2Mf4801ZTrrpuayXmU+iNOi0X/Kb0CF4TsHqxDceJAN1d
6HGl/mx1S+PFpLpKMJapUfmpX2MKMX1EYa7T5SIECoTUS34u/E5rdof/INDbIbnh
Zt23uHHWl0lDSJI/BLzzvFSf4MAh9pSKiA7ZowtwwwbtSK4b4sA58+nXAmyYK0YZ
rP9nhMZbjuya4JOPL77G4mQDwlEI9FmqzAYg+wd0qb87YhQHgR5koj2Zjoh9Rls1
OHHay+xhrWQJdeuKdzyN4+TEq51KPN53p6ISk+daO1krhXT3iIV0g+M/5DSwM8Ss
Fy+8SFqxGUV3Eg7i6xEnYZUGsDKbv8SQjbWQvPAxs8UExg+tjevkQaze/HFpBlvy
IW6FF9ZB0dQLlm3q0QuWCSRhc0rASMt2oKlWXzlohZoWbZH7PQKAE+nbss1pF3UU
cpG9ywopezivlem2U54DR2oreQzzY4u+4x3LGz08ylc9vOeLC0dFvfqLkCW5iZkt
V51RGt7Ojz3LNxsapaU9kSck1hLo8wWgk1Tq/suKAW+2Gf2GX7MHqd2qfPMnZWN/
zCKZOJtNoYVuL+ZSSfoBtk0EHJn3rbuZHso2cXX7eDDINySe1ra1mv6/6VWP/VuK
YWpLIdWTtadZw2ccaQhZMqXQKSRAeKykvDNL7ggYkjH8W9iYohdXrTx9MHO79Jba
3zpAybkv2TasmBWFWgnxKsXcq5BICXVkWhNQXLIYi6xwEG85LR8MHcYLaqoRx1Ua
cBqVo4+xl3N+hNQu9snvri5t3LzvYO//dayv8Gmj3cbjBcCLLyUhdbmP2S9Rlpe2
7v7cSqC4wdKQ2DE4f7kI60GDLf39Ph7uy2MTTm+5ovBkV5rKTW8/+noqsFB2lrw6
p55y2pNX42x/xJ1CrhFA/NcvrI8PhIlOsMPa5biapmhtuM2kqWInIfuxRODEY9ld
IR1HWgU6YPpfaQHWlDCD67x3XlY1xP240syQs0Nxkf5VvT3us8qP9Y1gzFx8N34A
U8wFEWscujrOSEN27LJYMREVpIkfnMLqEKORqLds795Q0gUefh7sL0MgNJimO9Fh
+dg6AsfWeZebuWb81cD+ieXHaY6q9MOcZL7jio4e/MJUhUUAv0OvsIcVTOmRGkIx
6vvn2jMO0GgN7Db2WwA8ME2zdLsIB0vdqHaBAxueoSgIjb4Hb+adJT7DLdf18ue2
oEAPQsiTJb6tULGCS+CqiL7VhOOPGw5BCz8XObwP61/Cc/9uGUY8SuFlBwytpT7o
hY7wlIZLbrX6cW2d6F4Pj/KBjXPgyvO7g1q+XBgQsgF1yLaE0wmzMqQCxXqnAY5W
RoUFOXFhAKwMj72pfrOxgVYOreEN0ozbgYPdjUGyP8LZIHdEAdzyqvjbhcyulJe4
jlbJARA2y2PJ3cglUdUr3MX1UOV4PkqoFOUSyolsRR1YFYwwKpWD8NjEs4pU6GUD
jv2A7xqYcoZI/stsak2zBDbxbVU0oXGEagiMv5m5gu6HSgluTFkzhIcotPERftNQ
lK5mTVG7KPcjCD4GUVfzd4llvG1uY/YaWdaBqv6XRaFHRYED5X66pNYvB+njxq9b
fm1vAH4ZJicYcMiX3exekY5ipJ7z7+WQd7l/kfsyuJ/86VqIpxYTAsQUslM2C6R/
Ii6oLNuR5A83uO6bJ/4obBSPIQ063NilJyYe+m4op39JDhxUL9xgOuwdUTeMrUDk
WvNP2LEP32TF+VxjNDti74DXT8B3pdlv43HErR8rwhsL1Qh2rQd1rQAbExfAQzFU
NuWNhQPnzIyB2gOJnNCr7pdWI2liuqPKCuD3sOHlXS+0BGiAX9QRPX84E6wLFCQp
GBUgirjnuA4u+rcEvhGX79vCl9dS4njD8a6CTtHnROKmhbcOIGOD63fAfrKh1ASc
3oHpQRJdkFSr5i+sx+GfcPJKzYqkNjpf//HP6VwEv8y/ItjJLizOqq3WFb2BN59r
1QN9lDf2NyOApEGDXD37bVAMFfkB6NbHdqM3C3ajfqhwWuZrNSHMUUAk8IDmWfBZ
zr6UfYkr0N/ysT+2D/OWFeIOuSTgOvlhuJm/kaLSMv/kmm53kJJII3JtZf/xXe4W
IqYSs94xlaGwY6pPJrO1dAJmxPcMSbVeJxPrFoS80xHfPUcwisLP/0jxXEVIAjoe
T9MZpSe6LPr9nSCbLNHZ4Zv1HxvmAUEzapR1aeKDfNL4e55GCzfj/MlnzC7FVWNz
BgmCKWD/HuO+R0cdORzYGd68FiSix/layBSsZUbYi+gxdKvIcj4YRHJEFwxX6a/A
BnYTlomC5m/NY8zWXOZqdBZZHSpBEADuWM3r3GBO/ynOHgnEGIYBdudpg8wBM63N
mBxUOeITrhYp3YVVGs9kAzDCgUcQkMO4Gwj19ya/30Jql/qsW8JwO9w6B0xZbrC1
7lLal8unb2WnUXN3lFTZmmO0Atift7CXn2U1U07aqfQDfxgQ8MhA/sUhq5jwD1tU
pmSwBe1DqB0jxqIMpqyIzDs3G9FMNHFUfbr7egXfD8bmDBan1N5NTCkBUlYYC2Tl
lKgr1b2khVG+02P5/LkU6+Ihml0NP7yVePkjrinqXmaWqqJxKjp0B49WJl3ifpXY
DopHqbTBUmDj72PQ9TQhWai+qFBSbJXBUHrkupwCpc+XE1aR45SAHcw/69RSVxtu
aew9DeYymoim62uT9l9NA9spdb2ScxbrSvxPpInwDNvyfUV1utzfy0nh5PoJJueY
esMOSj7SLOaGEkZD9FMkHpdTQC+4TW6YZks9Li8qqL8RCGYON2K92q4slviArwRo
SN50np7KLtfA3b8kbIIoLggQINfBd5eo8aQ3+UIrYuybG0MCJxYxz+SOX3WDPpZn
8wr7N5YruMBocMhD1kkH+Pkh7jF9Ztq7vz5Qok8YU00V5+KoqMXiPzHbQEEVvVKD
1Qi2/Mf12GeaNGfX2/jdAB9/cPJ6QfxbOHeJoV+xhta9CMjV1bjJx3Fdr/u7hdfa
Q4CTjYqaSC9WfObH5nE/ZzUsa7s6GsrbUVOVTmlTZFBfkjbn8mdSDq1K3YaXlYaU
C9uJ+wQSZvmM3RdiCu6C7CfXdG4xhtI1RRjCnT+2cfPOg5RDRTLygDlQyzFx4qz4
iYezQ4igPzo2D0gTltRY4v34fUlUtOYVYXf+ml8lXbYEy6p6UjA9ALcWKMVsDvDL
vWUkitlj4m4CwATo2p6gw3sKGz2nD3Rj9shSZqc6js0dvntm66LYgQQiPp18vFFM
JdDYKqAjBF4ZXPH07Ilb3RUympMWH3UJFPUxVpLUghbMeDc6AFsWdqGm49ic2r7p
T8d2BsSdI3PL2tR36dIal/6WNwKWQoCHUPmYtEoActEkoRKyXEmM41expvHEXQDA
PeDqHk94+4YehDdI+6doibLkyLdF46kWu9Fs5e6xJbs9fHWJTQgcEIwRYbF/n63e
v9oWLB5JY5irwG9pK1hDkmQKqiAG5DxW+HIMuFBoIeintj5K67GhGwJk6IdOmzLI
mMMFND5t3OU9iCUbp0uUqTiXiW3McLjZH5QjGhdmIp+T9gqBjOb/kyZp5UkBs9Bk
ykU2vnM76gvGpsH8z0IAYapfdP9Md7Rqg8WHAP/a1FcHmT/mNuQy2cbs007ntvMw
XWq1UNH8Y3kqOHAyXqjAP7ytLhezTwH5q1epfkiCCkmwxGjYysD2ymgLsE1WhNoE
iXeRaBX3jy9D1Q9mVKxx9H+0UBya/dY2Wom1N4ezNFO9TA8SNnMi2CgbriBN216c
hPrpJkZiecgwq2oI3T+77/LQlUuqHYbcr0/AK+yfLYw6kyg4FoXhMIytgKuc8YjP
sAaEjLH7yuvrYTkVDbuVO1Fsb2BDGiZQfz8BYppYhrMch/0WDo3XvMvNoTZnj6uK
LQkSClx9zCQirjFA86kKAJkU2VG4z2orA1T89LdtxpYB93ZyfCWxQjPTRoaahu2+
lKTUDJesi7vKvHhmekkTYmUngaQaIDXErP5ZtcsuqCkc7xSs/NNF3E+5umQftCBU
oCUZsfgKWDLivgWbpq2klRyRXeZIG7jvgb3cScaPLf2KQpRNZMRxSySQZ7njh4zq
f4T5Yw0qfcNSBcwd6t0abLSzXzGU7jIaBuGRkQGwCF2Tya8osRCQyhTtE/kAaUlB
5INu1fNd1j+jdJr+GjOckbAZVucBCjbr8uhdNdD6fUk1W9TGvkBlwyYiR3idj79N
9Zn3yBQbrwh2UXkp9zNgGraMLDwgq4z1L5qMo2VYoQcyQcWPGO9YPBUU0WDKzIDm
w1SKG73f/hlZOyN5kIOg1a7CdKTqEV8z6V+xMe6ToKjAGwOGjIjGOqizOPmCwM2q
fvvz3XkhhyZQeCtyMKVaAhyP45IdXd+mqAIggH9JPLeARyNA1QjU/02Tc9dv7HVu
YxRMPzq5uciJeWjq30Om+BDTtQv1XEUe+FfK4xaaXTS1yFOr3LAIchvWGIhSD5Wh
RQ987Bb50vNIeEcMWu4YDDgX9ZZYud8WUkDF+a+w/nNXr/8BhN3DDg6tpV3mGApM
6S6gZvbKYpsN3b5E3/hZ73sk1ZC4qoW+JHX5sLL7vcngs0qQolvM9EO+ELVye5h7
osTDs8T+B2GW6zr8Wroa9hn1AWb7CUKgxhUOknaiKaL+wWiCOMv1y+VOO4szpsyS
ImjDSbH4UoSvj1bJdvr28K/qDrV52oDD0Xae8AoWoWgzUg9qxEn37z0t1MsfIWCC
wwIn2A7f1jU2I4p2SxJj0JLtSPdC1dhRRW9D5MXnZsFt3zB/ybJNJYBA3ycFEEIo
V3WUonoI14HvjvpRK3MQTvZcowIeoYpW0911jjaXpTSgRMD2Z642p8NZO6uC5My/
1wE8GpyUF3v8H5v1ry9yIh49GYegGaLdQdQZX4AHXROTMhtFkRpv8NSwy9UKdO1G
mRyeg5HVnww6g+vMIG52FsirLNuhs+38BBZUa93rgU5iKuV0L97u7HgrCNxz5Jvq
DuJPiKwX6TBKz4k2pPDtu97wo3ViW0Fz/c7A9szadI4aa6TvgunIc3NS7qznVhVc
XzjmFJ2/oRGkAIntEqKUazIw5qLTt+YgIVxTCLDB/9JV+KA3bdlg95+DkS9e1qmE
cccSuQfSQocVh8DrRQ8dNTGJ008cmLkblcHSVpWszunCiNOlVfFfuaFF4WpgXiqi
ThIL/ve02490oG11YYbVeRhGfpbih1/xbxHW+Sik6ciq5oHmWyg1QW3Fde6+Jyq/
gkE1LyTQH80cTrBWrhpKi6LPoDhaQAT98Svww//VLib8fLMTAArEwKE3CZpo81qj
xdXHyCaz0oJr4R+BO1THCPgN+Sgjjfr+zQLDgDQAEI2kmbcoGo/yZxHWYqCZWb/2
jn1vEXCF+ocvwqI12dNEQa73S8uKuSJNopJIWEMb/WKe1el5M2DGctXf8LBRbjd8
L5VhixmZh9gGdFvBgoKRWwuVeH26g3hi5pb3U+Av5wO8fZQ6pSLfp4a7PicexlsC
ycDIdkxvk+h27Sk2/pzK06V2122R4YUNWkXk22O4PxzzgNzRWQ2diBKHHPHqP8z5
6D1P6mn/0aKa0jEycrHYzVuPSeQn2PD2K737f97EXC8EeFiv4T4uFrkK7oQeo6F9
zpD9iFBQxZYghYJRl3Hcm2KAOi/o4CQY0skdK8nycBtj7TZqJr6JSgFp2a+7nAKy
BHe7eve8wuGQTfz6b45LpUV7kQoJ3ZbMJhw4+DsoAgGGQnp+W69n67QxJaDDla2y
I2mb/ydE26GcAdpd37a0Lw1V+JXRIL+BriIyionVOI12QVAlF77d653F2nnlk8qU
R8suEv6gnql74JHJH6Qi2L22Mw8u0BfuoPaQ2+1+ojsWLgN/0gATyMiOIdyuEjbd
SQsOHg3o/73DgLm486oBHTTFYayolr/y1RCvIfNzB6qs/B0VvFbeVsosTUYtn/LA
AXgaFsIwzMUxmnKTH+dI6WTenFX/Vu8FYztTQI2TWxryv+Ek+ckTAcYta4fO3+Mu
TCQJILqY8qtI4u4hDN8OUls81UX/LboiZSWRctKWq+9ODVCa2fiDZ6f3Ea255VUD
kyDdOJwFHUeEK8iKF1T+u51cV5tqle8WDVWo5NaMt2zq0cAuQ0Ws0B1+mX527iRf
xV+ZQYh6O3iiZS9kndRBtA3pM3oihtlhnU9IHQLbJA+1U9DGrlLJaFYmpbwqTGa2
rezY1ct+hrr651oZS0c/8OnnC56I5+DfQXLrA7mqPSz1TjWNxVfNODU4j6APDCio
GFV9tGjOhmd1KWf0eVVzrJZdbRlpe+lA1XCplPxWdffI1qE4m8+lO5Af9PoB1nyY
SPlfGK6scCslhF3ZKOgc1ZgU1/998idi7nCtfu23YtExUt3u0Ty0XVW55CLe/kTT
GshKVfaeYDZ7/doelsLkff7haTjXPvGwRqLfpjHwdiYN6xvgRRJa4Pgd8ayMFzNf
d/Fa4cZXq21MppJuXrHDo0vFBHzBBW4Rw1YzxpFEjizleNmRziFbEEQsmZo+2hNP
nIOSIoSjcjpK93kcootlft8S9fQ4Ue3qglVpPWFaXJZJxfuJiP/jf6vzvutlt4yT
/ZvdkDA5Vxw/ozaeu/Z8O09yvQDUE6Oq5X2z6eck4aQoxIpgx2jao8Vo6sr9wKEs
kL+DldJ8laLNG55ydvDKlcPslhTaGd9hZGozijQLtM1iLSoILtnw7BTKm9kJG4mv
5uqp+NRkTr0rZC3i/Gqmytz7RNXL6NghgWWEfEcJrk6oNsrRQW57yYwQEw8zVN3w
UmaUZDJPd0m/OkQG9/B1CRpea1rgaDgLVY+O0fp950mLtlVjVo1nGEf+QLzu6pqh
d0AOpQax10f5VTxRM/ZDZDVJzcKBzKm4Q6OTsgIC3fTlgeM30MvzZeaRdmW56Eue
dbv+yy4U9QzXIg9JR6FMLdGE/iTEeji/BlGidk2KJr0/fXaDrnljDTfTyfpfkdUA
7prM+AUQLL00bgoR5OiGcok90tsDK31kYLKjtlGxvnggbf069qr5q9IqwAsXsbUm
NMiHYyw3EJdyY2JBhs9Q+P+jUP9maEfwL03RaUpumHXldytnUhQ4Dii+/fJ720BT
Jksi6JZwgHLHgiGF4cE10irrbU87zGcTdcTPqBY1S05D1IqrOjlY0vrDJdsZHVSV
Mk733IzuOc1Kke4+0yjBOeLvB+mcA43Vaap7iT9wiWjMdAaTH7UdeLViOTMHqG1k
U3oul4qGEGqdsaVufSJgV7UzR5p8VJDiQ7oznay/0qj6vcbjVhmMyQz/6nBZCYlu
CXPuHtn2YlrVAXlYR3vBKutDzYg9qdnNhhKgyVsiXxQhE+ozvdJCUn6o7+1K/GFr
Av7cPyZfJg4Om171WtvIf6vKPLNTypk4ft1ncWON92TPrm815HJ8YxYxe0+jtWiy
jPLtE/pcmaP8gjwqtn5REllIXJ+0588KfCw5pJiL3rsyYgotmCgx/ve3CfO9GoVr
qOT9TGKr/6Ot9Q/+UIIV9GlgXk2Wsb6/SwJdBtbX4uCbtC079xGWK9IKh7OeRYhV
mj5BecDZSx5+4rbyi+wqEWR7h4Nw/icNNksgwbHU/jAQ8MU900Ib/lSQl5WcOC7f
iki7nIuIpebF2Y3ilCpbmNOO4o1AooZpBoiP2ZiAZh8HRQVYOmheeJPzOuzYF4+6
lBfleQRAK0w6ORAm6cZ492UWRVxFPnSBmR+QHVEr4/9COEfiagSt2cx+jFhaTcmf
yOajBL4DiHVLDkE696+vD7/+uFOvlE3tm+u6Af3SH5YQ+KIFS4D8J3fmSzbydcfI
Wx3xGzuH9kOe3oclXTcND8ucvBXFlpVyC0g65KKXatrVynYrydNIwlb9LSC22gaX
KipuaMguL1AAAR1LRXvbKfs9PkwGFmfLRhiaakI9PQwIVe2LvAOnM3VxI8DkS9cT
eeIpoR2FbNs4uD7hHigrYr0FouENRP/fqfJ0OTCIORD13PUGh8BXa/Kehc7KGkJw
dzlWBhmnpWTr4KyVbTsYkU3gNXoK083Mro1J/v/7hpIlKeLQKPDMMgp6jyuVbUg9
Gv20IBvdUu3EpHe3aXQGxCR8Al9ip4EpSvmMcNk/SQDXTZ/VYdYocr3NVYVlLQCm
rBv/hnMv+SDv7X8wZYQNpp1S1lGcpgGZeBxqV5uAYSG8cBcn0ocD4NfBVPYARUAs
FPV57XeIuKj4Ih1fN0ls+H41xSIhyRoEyZkrZtnYjgkWr2LNyZiqmxlbFNU0ArHe
bP8TbpyVJOj8w+uQNIzto+YzWX5d4zbfDCx7CvIMxgrWPbr6qp/MLs1kO38gDk58
FwJnL0k2tiQBXDI5dAQ3OPRC/3+nDj9GwfoBdzng90bmv6Ie0zYlxZQbhgp69wTK
GvLA4n1M5O4uwG+AirX5f+prb6KPFm3qA6uFKsO58vGrvwKykLf44A5WrHFiHtF9
9w8POYU5hw3UKTXABC9r8zAvMh9F1MJpPdvO5aOxjIVmCMBzlyKTDAqV+yngPa7X
vNLNdKXT8c0e7dFhqdCco4+mKO/qtFxhhzhs/mg+wapZS6lL5gGgA4ZW3ABszpzl
n4NmYMl5+sn39GbfPNP2FgLgK23Ge1gKk2mS1UljJvMa98teczlTCJAfR7f67rYD
hVzvWXu2tPRRq6ObxaAVVX1qesgUTZmb4uDCbT1bZeIdK/shVKfnJFoaj/IwEytZ
6LHwdC4Np7wv76MQ6CXFTL5W1b7AaAOPVFqS0ab9H/M8p/SV/C6iMLbqVchgO/fm
ZOrNWfQpMuEViJovNpqipPKLMcsOj0t46mhY0TcuVLr4leTd7p0V9B40VTK3qFoF
+hXi1ozgKzONqCI+ZsFe+ZjtOLcMtMNqI52nubxGOra4LsK0xTn4dVrySoT1PlYp
HEESCus7BjgDS1OFWGWK2wXz0i5kSdU/9vhaQqvoAgibgxD5/3WEbrCxuFIrgdEh
p+YIfwjeTLz0nzHk+7d7DIY6zGtHGzBFrRFTy4UCmc9X9OS9mmUdqoqSUWmjuJj7
LtAxtR2cCuZyffdEm7bcZUuuqi9StglCnMWXmmil6mGcLsBsvnzyTfh2mXGY9FOa
BUe+q2CCGau+4WrQRfW8fdulZWki2s73cM79cXVGGvVYs/V7UEBFiPbDT2d/0kXT
h2ybTYE8y4Qxj4n3t6keI+y28G76OSUCL5XoRydkqaoNry9scVvTd867nfFgxiPR
9tObjfE2oq6aCYV8HmL0haukm82zctzFXUES7vhkfQ4P0Fhr2pCVK1zP+PLpfWrW
lKKGfp+zuSfpylaCd1Sta+TQiVtdorxgoDF7/Cj3Yi8A32m1u4VJSlNRk8ygOETk
DiCqap9JvQUnoCJkmaQYE7Pnq58t4VZviGcEQ5blQDNLUW+Pp5qJUSuGXNO8BVQb
8q4HyFxiLpiS6z8+NdI3QvqeLffps5788ee4Ni+guMFl03HiJB8jQ4NlsU/Go0BT
/DNSPt7xXyUCRlwwJdgTtTcDgckG1D1rFu2LBiw+x3ckR5Qj3K6ouV7WJXFrA8wR
32SG1h/E7R4xteyp9n9Q6Mv+7OqQISMi9jnOTEqLk4H+pqOhQBLLQXe8jd9BbGIu
BKY/vWydlixr2iXkxn3OWQOBkKja3d+0jKincNYuoVP6MhZvtytvSYqes/i8MMyt
7phPsZGElK729dILhN2Jm2OX92OvQQunKgOC0vOFtXnB088z8CrjQB3ZkryH6aBD
R30Gw2x3QlMURhRy6ounCyZIvONW70uQP5DUI+Ya7oxXNq7RttoeIIfWqji020tA
q8bscwog9G6mktH00MyfnoiD1NDz4FLnTK9exbNmAAd5fX8k7/Z32PTbLlDtSwCJ
JJxd5xKpCH6tOPhEA1zrNbHgEgeehGNeBJYu42E2+YwrKF+NOT1xSqIUqMYv0u0h
qDpqnm3znTDRC6fflh5dnYMekWcJaKbZNksFcCxackeGUAinnLoOMZXuFx4B1dMM
EwtB0rTGClbBlHj9khCqM7hckSTEteDoOFekNhtPPv2EHZvWtz/3Xosgb3gdkwfc
4RqfaKX1RuFd+Li3CWvpQqDhY3fbGqSkDV2eVyVsqZiSGrB1s1uiNBjgFG/9neIg
V8BXbHYac12LMEmJORwdwidAP1kwJTofYFD/5xK+Fg+es/gW0gD+VGomhduzvqzc
+FBJYiOIjaXwOTO1Jjj3jTFZB6fepkcaqMaqhowKI/hnRNmmRA5zzyoE1yqof47e
Dp21DnXG+y1eYmeOkqtYd7oscT6IMUcx3jd6CN4P0Lbn8IDYIUHsURhpW+IKUihS
9oSpY8V4n7aRCb+Eu3rlYAn4c/HvSxUSCNGhRv5xdT1tolV28Ay1wZDLrc2tetpG
fh5/+9kjfo9NXzfrfFoQ1Yc5VZ7jd5xso4l8qSoIY6edJkuA3JxMuoIfdBNdQlw9
DNPWtDbzC5loyD/Ht2yIYuHX7lsEftekEy5uLBoy2QmqfHN0g201hj7A59gdLhNF
b/4iikj3f38DXYgsXbJ19NbNCWIPTOeowboI7xo+LZROG5JZMA+BNN9dMaz7CaYA
9uDgFvVnKe/ExaUzmXtaUgeiIW2DYWWjPJYDpdIqkZ8T3nZjR/OLkkJ9MNH3Qtxx
fIe/6UrMdb0T1MLvjCpL3HEbmlc19yvZe+kvFis9J+zAy1JPWBTxP/UxRQ4SH/sO
5Cx5s0TusIvhuA5UMPhpKncz0GPlPigW1NLNzs05ccF6fQPsIPSMdy3BksUXAQq2
xVQB466rMl+/kfpOkD5qBeNLUmwt5CF3gWMpsLOsDdBv4DNZKqLQrkzm/zCwUPXl
BN4OAAdoh8QNylrECl3FUm2PtVig7a8jokd3gJghegHsYAj4LrU+otv17krL2pa4
LQSlJCQ1x2uHzLtRSuW2+sLn4DL98cXSTK5EWDBvSD+XK3rlE/ZqX5QLPzfrKeAf
DoGc+x9GCrqZJfzUOM+z2ULD6T5j0fz16SgN1+sP+K159tvJQR0sDpn/+7fDGhH9
0ESWpx99nV+4dRQrcXQXEadzrxW089ueF2QzJAZvdTeq+9BGu5/61UnZ4b0qylKA
T1roKwuq8w5M39K3FKUP+RU8/OWrawe86/Jlmzf7BPoNfufTf7Xwb0uZE6droXlH
ujkH7D61mBs/OYE9P94AAg4kLuWFszkPk7CaHzAyW6QFTPBpo42lCLJw/8Pf/CeO
aSJK3qzNINKFUMqp69zLbIERvIlrEr94rKXrz9ombgbC1glvafvMYQmhGj3mH8o3
/My91tIaiav3l6O1mnVba/w1zQfIhMXma3YMMppUfr5FHc8MendpZwke/SzxKryb
XyOGlZjpbgjW7tR2xwgoXDXzSOBHHh6B5gPkBysGuhblqnvLO6eegv0jif1+5WWq
uC0fPkM2+cMjo/Vi1Ch4cp6QgyVJkHxUtODMa3gMLxjWbP6t5iMzE5A8fxzjdTkZ
`pragma protect end_protected
