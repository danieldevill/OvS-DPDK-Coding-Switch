// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WzLA2xUDnQfuidmpQMTYuZ5EnheSYB65m9SLY6UJCkHRuqYpVLcZgAnBu47JS7GU
Tepnu7q1o+Tmmz0z89zgJGDqldUMAgknchjSsmP8GOFzTm4W/nKkbt21Rqwhka0k
KQLeE3PRKgcLdXdLmNjCAHT/r6ZvMgzEdY8d0XCYzoA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57008)
3h30MJmfxRdFGaShX8z5wNf4jaq0BL0hLa2AmVrU3A7LB8efIvVUasd5xMklgQvw
K/8RfWwHY+kgYtt7LA9mPo54v9VRZj81CIqgmSUHiUCIapCrSdIiyQKX2i94LnuY
mdaUN7LQx7ZzlWGt6D0uTTiejdOeFQ/i8RyxFase9TPgbe7ElkwaEVWaMjHwIKq/
xcuj4QB0p69G2ZbRQ2+ReoFfufEWaCQzCyPBFaXli7ouQIUphJqgW+pZ8V/ZqRi4
gckz/pOh9uWs2SnWvp/UEEkA1BfDps4gqJsQWVJOehx1kCqW2oS0T5gSB9bwL2RT
nTl4DH6qXRpro8GmNrMmS7CfyfnRfcBvgRtctV3dtjaCP+3CwggrOUMgSnVTmgus
u1WWol9ClugIQY3iEjnN8krA6yRvWIoOgJNJdi9imo2JguCHBUiih6hkoMRl5gHx
sj1i/PnIG9GzMgkOfm4XE7WTcLhH0rnxJrq0MjOJVmYmOpVjk53DW8WjptSw12uP
ZlauZQX9QnSg4elRbYKuqgXKG50UOGcXeuEpetQuntTrpzoLqD0lJ3wNAwgwIyRT
6HI4OWJjK37pdv1lX23Q3NMtaKGM7LgoW3FNuJUotEtJe61O4rjVVWTF1NsgyJCb
PEysMZTvJPJA8SKd3cyprDzeUlacsBNozJEgq7MO+Y/072VMeDg6q5uhdwQShIQN
XayfCM0miAYev+pLDkdoDtLCSOg4UG4AjmXWcE4sZP7iK3TyA2DByr/q3o2K9Au9
UHEg3OzlUZxaH541Lm3ukdvp6gTOCoYPpoGVdY0TD4uviEPs7VAUqShVOh6ijbT9
ZtZdbyjMKyaews0YKbwEBLDMvefvSnS5Hwjo6Ts01MdHuITt9/sjOUDGMXNpiWxj
AtBDV63T1H/pn3YHL9052YKCEpr0lF+SJP0S42wUoWhikgat+tNV933iR8Ijg2Tr
hDfnfCbRyPMYBz6UoEuDK68tHbXIsleou15Z9/06a0HfJAZyN/loHNfOdL5EbPqs
bZJgTXI7F3tlqrjj4YGvd+ApxGqM94wQ7qWPNtoTNGWR278j7an7smQ2QUio1xR9
aWl2HHsv6CZHCj1AMgb8iOKPAvrijfTwvkYVM1b2X7PXAQJw+LzQVbOCBwNSRLlK
B3uys9vaF/QdV5kGfIwpBfcCfmWcytf0DWvTAIY8gqhTUrECf6Y5SRDvfzuw+RlH
EtoiVXcOMk+MPF6qMERgEayj9MHKyzMgANfvo9R5dUUAFO0Kbceo5GJ9wf5C8d2L
uYfNI8tOm3xHALEXOsJ/8SQRs87rADqaDnW7+DNmblSbS41yozN74bTDdQnsYOd+
amPiqMe8YM2cBXSlX8JMUqXCHmDz1yPAMflICkfL2XJ5xokR/8MvvXy6EULePOEw
E5MFiLfjh9JwVtA4eoXBqlCKd4MtT86Dl2dO3DzfW8MWZ8MvzXAWuYV83XDM/0pr
NdYkMFyCPFqLmD+6267chk9NpIKAuwwMMughEw02dSnEJfnf3SE3uP3ZBg+nnktA
0SEOJV94NE9H0WC6c9Pssbpvcc0HyHXfZb1mA5Ra3HJRwOd/PTyc+NQHN7xWZhMe
iqB7EsesDSPv8eSAeHUaCJ+thCsGSC/qbzl8YJh+p2j06hEW3s/Z5HTPhu35Y99X
KY5fT7liyl1ASjLDjZolZ2/0x3wBmj7rVP7C7HUQfSMYqlO8+MHRr0UM0MNh6vaH
ay3yxtXgEwDLi7xjvVxq9qJqB9YYwpdtdd3Mt8J4r565mSj4F656pzbnn/NIaj9l
u8nj7CNy0o5sDynhYpUlZ+l8kH0HYtE/yPRb+ThxtK2tpvtyK5g36swWDz8PDflQ
feCCAAzU6sDe8O3Zic/1ZINJ3Tdv1tzhs6OHx9Wi1pmng9W9ZWodar36DOf266+R
AelLeEhu3XMmDNy3HVNJuvIwdFloaIUybFJH1F3KGybesNXAAoymhCACwddzrw0e
S4zjMI7aKKq/6BUaNJ97SSIQOExN3rXiIzgdnenIBRrrjlR7sI+QTTUe58s28vcJ
oF+5Z4A+FPIbHo7dMzNh1AR6/vKNPVqZHASpDhylLCEVjk1yPwJ22E41MFYHwJJ/
DyhUTsX10lsvxPAoJkQ48njR0fQ3WrdAbgGqBP4ALI2rqKjmPhe1mlGkNBNt6/aa
djgvmrpP2IA5psoeSdWwsRU52sPuNJl7KGb2b2+z2egFwyqedLj3c0vzoTUxHhoF
jMl2ZqHVaHW5C/qqHWuDe0wnlbZc81ps0/eQkdBz2s9eOJ/r9MyAJqDdxQs+cz0Z
oU2C+vul3aVSQr253nIhv1WazhKWfFz/I9UFPbrmf0PYxqdJyVzufn9Aw8sVGNEB
hAmhZqdX+Xz1hO+y3+hcR2ITqYte6kxuV8VpGVA/qYeCK5IhA9UYmTU+JffXznm+
O+b564/ZADSbcQpzYlBde3uCmn3tDTIlIw1inhYu84wa+p4r5x0NCP9cUGcH40iI
IOZ9LTVnmnQDcR5vUnCTZxZ3Ls816FknU71i1kC+lw8pEB7dFUqMkbQJOQVr2xsO
aNjndjFC6Z0VMpHt/Dshn1UbrX4EMdwu80/7pAxZXHxZWeJMYuhAucWzVcm4HXj6
1n5UH+9X4ngptQDtb1bBWhJYgmRuJXu/neVseu68hHLsuC98IrgiKmDe6WZ8yHHq
KoTaQbNKsm/iHhrtR4LbS8t/uD8DJJXDkFVAUFqd/i7j3Pxo6yfXvoTQiS/3Aj1y
Z0iO/1bQFtdpE9olq5FsO1s2pmJw67V9c/70OAVav10f0uIdsFPbQcO0G4lI+Uqh
T+RxTQ15HU06hnXYf9kENCW7x+Wkd1IXJrBiJwr9BxbZBrqpN/wZ4u5e9ekIDI/K
JC+qCjmuJ78nfULr4yF3KNUB5haZQYwKaxpoeGvYZJWtCGDi6JZiIGxX8s61EiLP
UgoKmFXHWHFKm+vAInUG0S5Rcz7nYPQraQQvq8IC4BvS8Lo9InTfih9a2H9u7yFI
eVAmFAP2SguH7x0NnYioJEUFLVsUCPoSerMNtfC+s31toyj+WAFeBms3hZ6Xf9ru
eWteUpLwsNGgYaEfz9kCgvQGjGTyGHHZG6nJi2iGpH4DagMOCCMlZhsoEecCP9b8
AZ1q1CjC6UEzGcQfuvXpIA1UIlDIYkMoQVIRRnNVQ04bJy92zqUTohk5xk8RhOPD
9LcDB2s/8yTkConmVrLeugq8baR57GFowBbmpOFJnyL3wRAQxO6KEe34+yZ1j3+L
wsmnxT9tOEdQdhbA4JA4qD+q8irtydla+lt3swsBa9C+5Vrfz8s+uOPYHr/N4ERz
ii45hulup/3/RVrK5dhW2sTnffhI3ieHzZVAgMwIhqj4bY0ypKC74rLd7p1s0KZa
yz4OwU2BaOC3Xfzlq1yEBpWRpvgy1V1V5hrCXGaxU3WFV6Fs84lwC4OFxkmH4Grg
hII0Odn5ZLSWfrvw0RMzUYHPCYzkrHj9DX6qgWV8XQctW1Fu6csSB/LOYKic284j
tmIFsnObKC91PuWKf6V6sIHN/S8s7JTCJbJLurr6qRO3Kj9Yl7MqNHnDRh4ebZqb
uAui8Cf4CVFZQkGEp52QjMegfdim4GfSMtoah8e24Kvq8fcgwgtA0vAzV3xZVf7Q
26I7RL4/OH0gM6e+c2vzd7DCvYwdJdgOfpo03rjJd/8yt1nJSC8/F+jawq+YQarD
/vA9Zv8CuYBsUzZMPtc1DIjqhJNrk7rvdE+7WvAwXZQOYUs7EvyQ4aZrOK0pQAVc
fO+J6Ah3MOin9kNp7i5OXxSbDbLUw4q17MuobM8Rfqv02nUXC1eT3ljDxAxpFEvr
UyTWJSOXZ9Aza96pjZjvzMkloprhfpcjuFIVO9sPJjQruXXOjdYRQVSSeIZyieT4
SaNBu1JLpQoFVSq3vwzAebZubKDuftJuVvYf8o13KcVRDdE9qZE5ap/CmQaDUWlq
8KQJLfAqUd8DbSd9k+m+1Q3teZOTv5j5+CDRed1oyU/RX5/AytLuAjAVabjm7u9i
b4ZDlNYHTScl8/rbBgoRDJ/z5qzkux9nTkdN03lc2S7Ia2tfturgH+hTkC1TIk1k
tioO1MunkTmwR47xu+zwix+38Rnnlm1ZJgkKSxvyRE6tz70m+lae3IcfjvUKrlGj
Bm3JaZDF8RVKelvBzIgwb8/6FyUKdT/aI2AOKCkonwEkfwYSNG0Y3TvkTaN+iPyo
jDkkBCD16JaEK8h6TPlonlUDo2iLqbFKfr3r0U/3Uk0q0dgWSoRRcZ/wAR/SkNa3
KH+yJd3RyFqQAMVg1E+EM7VMZ4a0cgqdJr/jp4aMobDEQtU9JEranP4TE7j0F66U
ZD+bbdYehp4Y3jHYkyZ2tI8nVx3wEwCTHJCLHG+/sqaqwrwa0azLyCRkOFtGmJKc
VsDnH4wJdiMV0SADrkZMpbeBunX4m2ZnQ9Gt0321PkiHW9GqFqDAXg1ngJqfPxH9
5j2XsM5KnAQYirkJGIovEK786GzSpUIqDBadFos1mQ7N5uXXZ+Xu4mvLhzgklz2b
glRbs4F/HN8LIZ8PhoNosmj/QuaY+HyoEY27S65oJYpwRR7+sucmTJYb+bUe4tU3
0egfWFfArLqvBCEi5r+e7qK8oNGhAZxYqjREuxQwQnV0A/UWtFFyrKIBHS4zgO6N
ZZ9Pl0dttn58Qqg/G30Y45TIcUURFGHRBv72LJqRFwb8Q1Vi3q+W5URYjoK714+n
YalvxQclWNN1qejAT1Q7gmBQ4Pegrg2mmBQAoY7xnQRKc0xaXkh6r+yKWmFyC+Nu
8Bsvb5PpuOraeUC41Bhj2HZcX+/7UsfipSy53CgXyl2baye/ZezJ/zoEvX6kZVSb
hHUBQcveROMOWqXyiVP289dsusmA1Ez5CiV51/1pExxQpHDpYSQrMd3GZ90P99oW
sUOHhAs+hknh0I/2lRwCcQuKw4KqOnJI7hOBZt900FswG2STxiEf7bfvSb1TGjd3
puXuNY9y3qTj+D1e2VnWs8VZJKQXh70OoGCrsBy6mLIkI7Y5DXGvu4PzZXUcaW38
TkU25FHgTAfnI8EK3i1dn/lRuoP0oHVHcw+s7JSFgw9gt2KrW2Wv79Ua8f9ZjA9U
IEEaFRMtVJU6h5gm4GI8TY3I0NbKk/9y/esEq4aajLVeZvwg21QKKZBJrniUiHHV
KaafLPszbp5YGlfGPJmUx9+hlQXhXqDhM2evtSinq4SAuebgmjZayZCrSZg6bPsw
f0fefHvIXfvaAPskl2RjBuzORg9m7uk4fc20p1zLX4mB2Zgs6TNs3zhh3FEKj+4z
ux7+wsuFdwzXxg96cHbI+nHuSHkAZ8SKiFgvMvEFmqS/k0r1ZTSGrwgphs0cHI5F
7fBDunG2GOTYLQiyB/oQIvUjFucpHynIAN7rGRPPDYSRyInTmOizuUNNp1EklQV5
2ciouW6/y4kQB20H4oyKYIvFWyHW5JwI7pKK2yhfYETvgXk3rPDbMXhPRkMY1uXS
4zzhVv8OrgClNOCyNxYg9i2T2qWE25ik9D2OBzHMnIDZ5SttV6/QHu680ESpnMAS
3Rq6XzEY9y5AN+kT3c0X+QWw22q3CzUyN6/a+Ft2WpenCPDP3a4GR6D28OKFW1a5
JZ0BpiWNaFvu8EGUCvGX7/LGzn2LTUzJnfzVkJLWxA/V95EuXPVMyd973mUx4g8m
oHb5Qf2IuFPxd67y+q3qy1PHG2IRKFYFFf+JXVlG30HWkXfdT/9pw29Crk2UVPKZ
zJOMTZNE1cEr/nDnJ9fv7t6VT6TcWUlBCVE0jeP17mciDeLI8KAYYrio17kojqzq
WEhCX4a3IWlQ+0y2JI/gTua6ugSsRkVQ3lVCboWC0uWwJ9Cnxx2l803eVn6Tjdtb
fItpD5u+MSnM9MKFwOB14h/h6MyXdSOd4eZZcuencGHJTdsvw6Yq20eqJHLtbhHq
LALibym7Xy4Xq4ZResgQ8c+9HiRexLBQHI/wuqlHldc6J7fmZ+03wv8jJKSrTckf
mtKLqvQVMWk/6+xLkdGJYKYkdu8IXCzjeSVk4Zt7vBVs+v781iRu2QwuR1OHze4m
sRSC6QXtNf7m6GnH+94RgoWhv2a2jPs/aMskQ+OOsX6cyxQPd2FZ9oHbQrUpQ+j+
pixikkxZTcArfh9p4s11ZWFJwl6j3Mz0l9zWHHh/1wJoXQIDJOHg75PW2ytQiU+n
FjAKDmlpub+KW6HbN8J5ae1JydFwGmZwBYb8Z+NnWeZ4KufZnqrh5NCEMXQ8fumB
Fxu3wpX3J8D0RosT5eWwcCchDpGO89oDZWXXzUqqwJ6/IQe5u/Mp7YGuEIZXXKEV
diWsnCnLE7E448Vgk5cpCq9syiEK+5vxLYRSl7mtgv2sPcTHvHYYZcheuLmaVoUE
6gHzXT1IXJeULefIIpAGgn1gKdROkay6IuoEpKxf2g50WIGUA5wHBSHSaiBY1Gqx
7fGPw7dxcBIfCQ+uMqAmQwA2EYvP0gv4kjGfL2jsZQV9txnRKXcRJTXYpVeKhSCu
GdMz3AwE0LWbiW4BciHlvkgZnwHure3qNj5J8eIhDQVpwYxTi7q56rBQJaoLBMbJ
E17WpIgBMvQn/3V70v08WdRWwQHBKLaOw+0shjrR/wC1Z/Bq/egYtNkpEq651/Z0
7uyNxwCy+jXw/BHQ/yQQpfeW59TXy2Dihou/1POoKBGgpuXN/6EPdjkIbQ9B0Txl
GIvSAeFOlheBcanegClA7xtIGpWEVGc6zHLPbpEX5LvIScAoGd5Df24Yqohm2MQR
r/SHcDjFSjniunAEddXWypzfYCimyVkKOLzKE/Dc7R+MufdpeBa2SXZvwG5GwHy8
zSm2h+WJY+oFdAK9GbcSwu6cqNPpFHxXq87tCRIoPOJ72PM7qkoPZbXHXBOj5DKT
jQIfl9XSSR8RcTyJ23TTy863V5XupjXY7vkk5+FVtEe0+WWOdlToWyzzRfIUHFPz
wtmGia4z1h84LTvhX4HLybX84rBjtLQhmphrsosMNbf/tsjZpGA3ddojgONmqm2D
HTi30TOiXk1lB5DO9ukmHeJbkxOId8E5MvZeM/dKQUGz9svQtaYmktC/DO0q1NPf
k2QbuA58i0gbBYbDOaTk7Da+npp9VgfaVg6vVawZYCcvUbFTM8EaHvBkAyY5YqJj
9jBWD8739SkMa3eIXzjugBR8D2TZ7aJyZESvAxW7OTDH5Qpf2yXxdF+VJO51EExD
B9DmwEPJfatf65exS7e+HQ+OBUm7MzodIyk6xlbVb0frCvAfOaMOPwAK0fHxczyG
utThuu7l3AWgSp3F3we/LDr9Yg3qW2xSaHgBfPmjZRZ57+1ah4ct+N/2/60g/QsF
NK2UepwLrK/GGEQMI7rnuQkxdLwqAmzQPfdRb3KndxHEFjKFcU4P2PYls6nU7x4k
HJTXX3H/PjSIJQtF2yynvY33toJzNM/BD3dFHwxLSxjJGnRg40qGto7E/BZN/W3P
T8QHFfmtt4IVGFJVHU7+EP4VTOJcjvzlkKi2rgXgehjb5JtZVfelKxOUiA2xeVdA
OHdprJWKAA7lGKd5cLyPHbbTXO4z275aFGdd5jQlwCtybH/BoE2pFXN/qyTTWLx5
NjLmwJ0FWgWcN7f0TausBryuNsBg2/mzQ0Kp0lXobeaK1UQLVPX/3yULiPnwgsHY
ZoZN+Xcp36yJO4Q/kLeM0btxTD9/kHx1d18CFamGC3W2y8277/6nLFq9W7PkGKZj
1XT/Cjp31DEs6wkJGwRgrJw6Pd8emPk9VJ+3hckfnaUNy+clovg/5nrkjLwJveu+
CSphBZ7TjpXwnU/psl9X68wJVj32tFoAH1Jn+7eGAYYTSp44uWB4Uk1pu0O3Vfqo
4Mm3agx8OYYyaVJ17L+9PrMqR8WSPAXAcje9ZgZLlgG2+hV3lgUgB4hwd/xL1EP4
xVd9VI2uHDHjAjpI/nJ1DcQHHl7r/3ileCaqjpy679cak4Sq49DnQDM2hrXaVl1o
MpZBVexGG1Zrdp4qxrec0L5b+Tscz0rzJWLqKqsmDnYhGs0FNAnapB250wzh8nic
PxTK0WHKUe62y7bbaHxJYdWSLPcSggMrvov85ZmEdm7jHYbMhJ+2aj/ihGTF/oSL
McA68vxWT2EZ3TiaJH+LbWOXt4bt8gVEoGGQ3MLILY61GV/Cpj3gynYQd91lN+T4
J2nFhEI3UNwmX4rf2TvktDx5vhLl0IlGmXtEVNhaZdpanauRw6y4kJTOiIm7EQvz
lgwMER9diyvSv0uQx5nNmyjfSqxRIpU5sG+8tZES6zOTi5F0lGqjKnvNGZK0D/0k
ttrt2XAwMPY1AzOpQFrRUObSFdMNvcrQVr/6T+DsqnUz4qVYbeSvfUSZCiU+Xe8v
xE8cvAoMRyqVQCsJdjPS58K2z5ET6OPK1nXa42O0E2uW9u0wfBwsOTFnEKYyjw/w
l15QYe3MYOjnwDnZdFeq1HV6C9lXfM0RlslGypef2idWxfWH4MnawExuyHY9dlhU
grS2C0ZQe4yFVPXwA0YXBimG8c/qq1jOO1IjNK8KnjIx4+XKgihn/Uy95SRQnZQ9
IMvYvB70k4XbFD4BWFxY9TmVZRvbFA1PqmmJXccbGnoWFE5PFHxNe6ERsWOJBaRT
QZdMSTWEEMvBQmFqM70u+5rpliBQJGvBs0sIZURJTGGK1don6z+HUm5IlnFyCvmm
yBC5RayOlCrMXUJdVyKw0+Ebg/jYkCBJhsKHmHRdu9IqtScZduGnXz9ARlSbdJ9s
90+utS0nMdXYT+2TDRv35Jp0h7FGDIc9pklHcs0m55D4FRgguUYP9+oOiIxATdzI
YcJidWI6QmtfhSCKtfRpWlZCV7qRf02t0LFFeKAeBGhROgIf+wF7PtoocanVV80r
OT9GNtYlq2duW6s5yYoPJt+S0LUAZGFXY6jjZr2tT/JoxL5EcnKBm7zWh1aduUE2
gmk5hsQMRzeIQsQWTY0yIYrcY6RwQO7kAPbpx+z400JdwecYSgvJ+EUnq+ZvkpDJ
gAy5ByateWYng0ndY9bV4fQ0DfLGRjNVj5H6910ZGUoq5qjQwON+ssqqCPH+UBak
iQtMQtae52RSg1ZVbd2A3HIYZvByxLhYYuauBgvEd1Vkof+Rd2XdluXPRdYlzfRk
eVAH5bwRDysXWhA1dKD1sAlueiNEbbL+YNEDMbsAY1SJAe0GccO+UYP0Kkxrsod2
sOoIEX6rBQSTNxKtPLvnbwIOdh/Ppk6QP1CeYO2d8pGRIEFYOKdEpN92DW42ZGLH
Y5bfd0rV9wCDcfq61ZDAL4Qfn0ODTUCg1O4Q1rSXi/Z3f3F58FRJ3D7lfpyCqnlQ
gzM0ZZAv6WEOJlnwxPAj9cdnfzefCcZD8pFkGFxxDlbcVEfiWrWxXQQwH3cUBifE
eHeFJCMBEMtjOenVXRS5YF17ECt4L1Sq+nO4P4JCuwso3XGGiDQ9mCWHuMbXv4EX
vYAmiD3RoKkA63jKDYHCqhvH8tKuc6d5KQSXgQXpWn5Dm/UmafdnOg2iNx9g4Mhc
hUA8e2LI5zTlqn5fu83PMFm87YzL2H0bs94rag7cACWqZLGJlWLwGBMhsXD4lafk
y2mzL1PAGp//c1gjM1CBZnURsPhNCTPmtkq8pfkQYxHCP9B5JCCGsKgSAbhj8ImH
zjwLOsDuJNYiCL56hsRho1OZMsl8E0AI1w0oX6BTq08KLuTuTOqCHz5FvNCGusjw
yTVusFUrSXqvDFf84z7ZR7qM/Sb50igxFnPe4ZuQM6SX5NcPsZsX9kk003eniadZ
nw3uA6YLA0yumJk6QOagvoMWyQfTs5W7VdZxMPSz8HWXSagkpX9LAvUsjp6NDbN0
jLzeae2PxZBhWoHCZzu8rF+Be27Z3Gm5o/f79WLf4xcrIMlDiZ/jauzPjWleCVdE
l/ACyIRHzghl66a1vT4HqFLIEZryg1hxsx70Ps9xyakGl6IgZesStad4SWgPkBqD
H+q2ppc+8DCTa0tkaEDhXCVzW03WtHkcxlWhQZKPcT50x18buCShOewsLrnXI32H
G7JwxWmfPelR2DziPYlV+ueoWo+YXS3Fw08y/7uwI5FsKckutfBvBlerYYIlYsYe
Xxdyfvu43M3utf7Wifmh3KWllOTXIwq/aKgQgYAt1dqrCcUWurdIz98PbhUW3xPK
Mi/FdaJZUULNBRBZD7cGMO0eqca46rfzPyNS3297oJ0dWm7uJ3SKxEMirFTxFP50
KKrgZcqTfsaEAuABDJ5Ugboo810FAJjvt2LAe4qqcoSxdFgGl2X7txV1iLF/RD+o
RHTrOgReS0uJcBseAPYXwOWxN175bnsbVWlVwcCnLhx5Y1IxRjAItFUMwH54x53K
L0sGOCkFgdYXKIvneQ6FWePg7ucdtsDLJtmKT7zrSXt9pgmnxgRt5Fw9mPk7+jhp
PFzkGbGIke8px0OpH9506n2cK/Mmty/kTAQl3ag0CBTq5UPfXKWvSj/dOiPzdn6w
4BzLtBu1/GEvTpcJRPw4cL9mfSlJdr20qYQz9z2SaCNpoBczCjW57gO29LzyHBj1
5nDBsRvJeEwSfu0jxY1DM3rpVpIPEDK3js81ISI7L+1sMVq9FrTdRwCXgTb6GBAu
v0MOcut47zX+J6mN3uZ3F++wfcJ2w8Yxd9n472erU+XtGKlibD6vSSDD+nVR8Ztq
HrSRD1UHw1swRCsLAjwyyjFKfMOCc5ie52pq0mtWj27Zodg1yNVu8nDMfS4gXUDJ
woi+jijTvJSiopMIcGCZbolsBubCpZNPAQow4Yh2Ec2hKQ+sb2ruJ8zQzHaT90SV
cIqTHZMz0pVceJs2EGSfhoc297tcOlbKTcG1I2YFd7mE5hsxv7z0cPFDoTi58Ax+
JOnsVLd1LNtxINB3PqFifPSz/UrayLEpY9RatD+qX+3mRNqVVXmiIv8OtgSNMku1
5Rp9RT93eOx2zgCWDEUJeHtcvaJuNV2SCCH0yr2PrLA3bn3SvcHlgiPqNuqwBC6s
iLvGdki++7MDG1prhoD7zBazkbmMYe9wX2PH980/ZPquHKergCS2FjHUSuXXNM5N
PYMNJTKf79MNZNzsF3AdL0oXHgJal/lPVlmHzw7qy4oazoXfpAIzgrBfqINGThvD
e/sY+aVKz2x33q3ZVVGn9AqjgD9ZeQmyumG4ISSOYbN1d3lIeQBa72zIcZa6MMU4
Rp0G3dM3SX99ZJoLZsfXUErYLRphGYK3p1Z9a93VlpUwxBYGvmcBfs5Fdr0m6Eao
7KajYHWqZuf1KCTPnosZ3eK0hMu+HdKeVj3mZajNe7VBSdWaQDCmNQHC8K5DUcRG
eRI9d41OVBCAXCWCjgP+eOekl+HqLDRAn40IZ9ATx/2/WyLAa0PzuHZ7wdCaR+d5
DhB08mdtRI1enlzTOhiudr7Wofe6/EoLr6xz3EJi7SMveg0GAT+EiItc6Jg7Cw4H
dLWusP4VZBVS2n+5PhgGOePiXLxKk9r6bzgZRlljuAHBY4YEF0SIDQk4zxx3+xMF
LaktR/n5N678M6a/CdEeK/Cf/RSyeNs2mefuxzdPzUtjBLHUQpqtXm63XsjgzNAQ
YcR/LaVGHWn2CXCwNi/+Puejg8FXO+5rldbAJZYXkFH1Zltn+xWIu9lEZBFj0Uqi
TsSfFfgi6iWHhKdECEXH6gtjqd+cC8u6m9T6oyKJe28/P/vBxIRFElCFSi1JLzF3
TMS+i5AlBYaE58eX8XpbaiP0UILIWaWkjJ+if4bpOlABgxojHWmP1N53yFxUt+LL
fgJkSKyKO9YUyrxYuy18YdQAwFisbn57sj07oxcXpCCHgjpJA7M1lVjzD+9YCfFO
scOiLXlDt/0Ih5jlGysFNMN/5PgGlFo2+Q7CROWG5y0/7RTgO+vwGsNIiqiIDS47
FH+F3YIgznWHRYvScgUz/h0JldzYA3cGTeSN5g67ow5QyJF6iMjuDvFRw7kBFBF9
PTkTxRnV7nNz212UPq2NDHUdjf1Tn2PivDstcvDnRgn/67B9zctLSI1O4HcLqaO3
eUIXgIysgGylj0/5ers2iHnKpQZH3NOmkxVo7RMPwlfxhQFGmxSgAl1OAQBGqnmy
P6qNYLgG3UPqsE3Sv1D3AgWjENVAWc6c+lBXQ+vfYqXFExDyWvm1nAK0WMQbFp2m
dBQhx6OQdrYVe334I0ATQkG6zm4jsAPiMqTVpRwdP5eZmgLoov01VEt81YdeMzvV
PXsGHvrE8OQFGP/V3tFjIr+gUi2Hp7RwxQfTHo7sx6AXxW/QZCzGB8YKBRTPNcX7
hVfwZK748C9VZ6SyuW88Hpe2/SVZQONNPbOPI5tE/aiiNiXa23A31jtUgBisYA6A
3dr/EDsRxIH9HBTT0Vu0FK4Ig2XNHRAYnuWbnH7Q9fjTgO3BNsaETr7fZ/yIssXb
BXBvB0b6OeertwxD/E4EPlnhr0p3gvz4ex/WW+2bSv/pcufE7PEgUNbIM42EgbDH
zikd94cFQXYHAwRmjcvltwaRIUhATGHlUXmm/0f2XRTTibjvL8F0mgDJ5K1Gf+CY
BDhN11yErdSEa/XJEOWntzcW0FoL5nCtSMtORdfIgWCZ9ApJ5lP+dJJ6GTxNJxhq
rG49LmyyZ9nLRbNlO1VC9B9VqLTTCHc+YusxoFh91UhjRmwcFw0BnHGf9Uippezc
3e47g1qa8katmouPnhxezxC+2JMLeLW2+XJmT3nJ5f5HMlLMVOFCffUa2UOYYA+a
ESouYWsXG9Fd0mfyoVx684BrsqozUYOuLiukpx+YK+sULntBbpeAR6MNWaIEhRrq
u1I8+lWFfpId/xeiVp6yOWyuUdeGkglmvVVxuf0NT+Rx+ZM4eT+oZYtx/tlk/Txs
MYAQTeGC257LtQuD7ePfUAJcSyWL3x/11V+mb1jmasZ+fURni72WL9O9zJFeXT+g
6LYKDxE2sRNXq8S0a0wHbuiAG1gtqFu1w19PsyOkIQ/cX5wPaATt2w03Vv4Ov+ss
KhNOBw6vPW0XPJoUfq+huiCMpkc7jn3aIoF+pSrP78J11Ifg0is62jaIgP2CSUuZ
3IUfSDhAV1nhhDxCHLpwevbkCdAz/WwSzXhx7V0MQRulCZ9LJh04sIoy+ZWs2LRg
molnhhhhHlNBAyPDsJjFf9QJ6gTqd7NEOFn526R0tc/sTkbczcF8fnx3cxtqNLS3
4WGkwTK9dznyYr39dtUAvDnHsgnk93itl/3Aq7gimrwqZe9EroTLSzLmlosODNLI
ofp6SZCHQEWz20DWbeVDG8Vr3UcCgHR2+9qBxeN8wTdqtTCsCmZZZIaHLglRi08z
EoCt4Q1RDCOKsEw/A850oBAjkAavi9IVajEBx6Fvq2RZcYMQb7qhuKXH+eyOhTM+
F4a246DHJ5QWooA8Jyh36hItSxJ7QlUx9x7nwa+c9/bMxIobAvw9EcT6AKwG4nH0
ujJxwwpRaTwSuAv9Qq5h34l8ekB+taedLYz4l3JZDldyukxLhPSESKd/TmIYo1jl
CgKo6Vj0+/O8jt3bzyf3vftJzKIlCJPwAIY2CtUYJQmT9WYNlsDqSuugWDTIfxlu
bZ8MpGI95uY8j/AZghoJT+wF0NTmukXHT2tMlJ2STxjTmWDjmwHjDNqyL6DH3tOK
9vJZX6YEspJWKB/jo6bwqRaxOFZ5e5ZB0Hs1PUf4LRGT3JYCuMq3gA87ldaIybyS
oDlXyvJLPbsEWQoWSl2Dp3v0AW43fTQjDK74ZrdRenwVhtGa+zqsJ3nhZ/8vcqjg
7t3Kvd0Dp8VBXef8c29c0oen/rX2WuJ/Ky5RFiSMfwBTiYlMLoJ26jSNCo7xUxz/
wpvNIs5uxb5zCmgiWkwTh6QtKM+n2f9x2cO4CDFVVlwxyeyMJ35LKZnA3AUar9C1
RhOuGfXnIQlIYQQHBSqa4bU+3v12iIvS4n0mlMFAVML6paJ+F6nOGCgU+tWLXb9h
FqnnxPiOZtOEBD536zfs5ZD/MN8iMgusakWbqKHve6Nvi/wgFy8Pk/p0mnkEfoaF
+9NQMjb3Qey+5shRTNLXeUSlRt8zcrFZIi8n3WhRas5tF5NrwABrdZCwPBOtYTZ1
uMQojce8EV8t7ZQfzQ0hAbjllXtBOucXY/YokUCo33ip99jToRa9RrR0D+S62S8u
fYmi/7LTZZ8IB47HXrKaw99SKt3EnCxSl+crrC4FDLl+yi8B0ujuvqjjV7lebaF0
dBMKu5fTwVF48cqFoUA0IyKu7RV3FxMgkkm46eRm/kMwZNKeGSOmBN+ZqIKGyxhe
QF0gf0+5IsHWPikkHyMl9pMGhbdSnoU3xhVmR8P+7s2ZF3imVl7qfcWpRmw27inA
iLmFNMIH0PNtZ7dBGiERFg0PwO1pYbLuxDuWUhX4eQOTtJ1+BV2FQ/SFTjdyTg20
wEYSa59+OHiniyyPZsS9fnxjTFrevvpwiTB78zabywk73jByloNMqRq0XzsMXhIj
PvqL0Qt7LVLz3iKHRNAgppxl0JIzNubsuMt3Oz3/pRHo1NqqlsTFEzGr6Tf5NPKP
zMrUqnkqtfIezkRDKN1FjJjvejgj4mIUv0y7HIFzTo/HL8kHU90ZCQeq9tut24Tm
OjNOzKQRaamkEfroRw8Q1XVVWXEMh35MQMobqDikWq5ifBmqpEZzqNs2m3uV4Yb/
ayKppG2EO6Z8ylqdeozlzst+T/nSxHPUBH9ANLWaQ5nHNlByDytTXXHTZ2A3YK1l
5EvpnVfyGR5uyv0W7Je9VURhWQpHC0QiC7VuR8qlDPHsfKv+c70ZzJemNlKok4if
0QhTPq5DaMQxcYcbg8nn7F0SfYQD6pGarU1xABpB7POvbPrCoTxwDqX9Ouoepkr5
k6T7jsJmxa0OYz7kI8hDJpW5g3obT+sE7lOeUwL+hVggVRsDstjb2XNjOl+BDStQ
dHr49riyFDhcIQz96cMDdnLxjRlgMOWCb1Y1AQfGNQfS4JHJ+qxGoOx0zGJdyj/W
yNxXlj0t9xPW7XwXDSgdg8LSDn8+44p4X0rK8qMmgM8PLi+m8w8aBF9ebq2BI5Bl
JSsMwF1HgT9pHTylY2htioB8jy3L7VGYwaViyThgpF2Ex56lIpzggpwRddGHZaYw
4KzJAXPpm+0XcRlDfUt8y45ehDR+QTAldX+vW/XVyViTL7dWa/T4iRUJ6T80rWaO
nFeY5dtEZ0D9Nrswbe0ok0hO8x6CvDqVh3R7H30zEm5XNSsiUQ6k0lDDNUd0uvXZ
muVsTcKDBXoAjLP0+DTI9caUBBi9sQp2h5/ZQE+kExx1+A3G8FFBdywkhLvIEtAe
y9kE2tQA7FFz7rivSUMMjxtSW6/jOkYMBP9mfNpibFdSuyybMOzxeLK+eqVvgOZH
HV03a0b+pg0kmvLUmeav37qzG3x6wqON/qUT1KMyUQhpE9SSQSzZxLgFqGAgbd9M
Br+zzBOtNBy2RXMPV5byitH7OmbAgCBpKchVnaq1UYb+2C6uyTLPU2OXpdrVr490
MfYP93WHe0gw3IIOoVLWI6qyThF/GaPJoZSm1OnOy2Mf90KGs2pyIeo2qCNDpAWK
8eaEm0s4CQjsNT6hpiNRdMfmtGS8UJQThFMte6HX39kePJLxKBNiTdda2dbdP0R4
vAXDi+86U2Rk8UXhuM8+K8J4Vrr7jXuq9CSmlY+LSiSCPa3zJxBYGN+NWe227A1Q
E4JRd5eCpLUkW9Ny6MfHHd+/l3Hj0vkzXS2ZZ5B+knnrG+tqcf0LCmNpo8L6o6Li
mHygiYrc77GKZmHnB5yh6U2svochcCE9AA5AAbO2SSN45joqzwtgQ68BEEXfg9/p
L8PTNazglk7ayrbJQRbHQqZyqnxeajAOkDQdKi0N0Xvxl3Ui0hNygloPkEFCiHRF
a53DY9sXgoiKVrEcWqIapgqNgd8iF413xkBH3cYu8tiwNRAGi2QaQ7znuFx0OmwC
lnfNb/oblg8OCLhfPcmGaVJzu6DtJw5AijBzQsoEJJjh53TU8wAlrpKrsgyaKfvb
RS5LSoe5gz2aC9LiTm9UO8rLOOewEqpCyA0fKHrfaWjs8GQJV4sNr9HGc8AtTJR2
KcQvh0qv6Oe9QP1zHI2F81UpXkfEldsymgtnQ1O+6nvPRO0WhgVTOhCHSqPrJGMS
l+sDWkdyxz6xkS163xtSHzjY6DHsNyGbtmP6uiI4SmuGMlkzdljjJ5T8bKQ6vYdV
r+wJxJenwzp5+FQEfY0flruS0oKEZgXXzt+JPE/LqNmKeluWKLNE26JzirjiJiWD
WZu7emqez4ZkpkzPjLf5SyUB5baz5iJhVDWDdUwaDD7uQEPEMLYva6+w54E9Ecd0
Z7h1/zZRJgq4Qed89kNTq9d0QPLfSzApwpdkDR1/GXVJhnQdtTwrwl1s2Oixc3Mk
20J005uAnzfUFShFZdy6fk17cJa3yD9JNIoVS/nCwhxAJ4N/mzafnoNZAOJkfYxP
ptcyjI1ojbhMegnYbnaPiIXGms2YlmK6CiiAMUIMCSvzQRQ0VByBA25SNfAGoHth
dGLeXpKVZx2KdW1IEMiNS0Mb0n5yVvHZgTsbYnoaoD/GwUcJ5gns6caXOR1TBp+b
drZptNJv6rlcueOCNcC/C0Vx8LnobU7md3E1N0lzrr8W6Oq97nQwKjVIyqIUFKuU
pnBkRT+O/kc4IvrdEkl6rshVTdnDTBG/Kqm/TqXq4p6eFcj70bqrtBehYahAATdP
/R07pOU3cHpnzMBIrH1g1ymFIeSp37uR0rfhddSn2+MdK7uj11nZwU69TfLfuX5h
FnkiWloRnIJ0XluXERaGeTLA/QDv20nCfYgydQ/deigkZEotcTL5lLmOYkb25Bwm
RN40fwvtMRbUB6gQq8b2xUfPq2OADR1Ssi1BKLsGHgZmlFENxOcs2JBJk5Qw86W5
xwJLESo+HcU6yQ1hCYTjE4z/2V9w9KRVt/Haey3U8P0bzCLmoKIj+GSFVUF1DiNo
3l8IPbt5dJ84At0VEcMfhjp1S0joDpnlcmyTY62OjZWUrGoH8XWLvPelLAIXlcI0
vAQUDv4vZRdq3iszLMq7191Qmja3bWxPbgzoEgipxP4UcgAqby28TXTT2HPy6mzr
PgvrsW8tyIOgBzjkfA3AhtWg0eAppPzG2zeIFiU2MzU1wVry6QVGafqivuJG5RfT
9+FsHrtsiqzyFtdTO4pnd4b6hgzdawTN/lECz+/4D/jjxPwuHfg7vs9/a0xce2FN
j95p9rHCCX2944pbzSilyuIBXxhrhvPC6Khl+F4Fl4UqeH1a9H7RzfjaI2hmHvJ/
ZxTZ0IxcOA2yN3d2qi5IWzpv/azkWhC7z8oKvnEwQkx8R91Mug2YmJLdJrzqiH91
xkUBnWuWf3j9hQVECuL8zFHZOMwpSpagNG4gIacLUZDLa+gxcy4dSYfnWn1JQ4PW
9jM9rbjTFFKRlTcJR/4XzMRaYl+Ls1S/NMxgCNpX2Xvj7yWYK7izni5UgJJz4TuS
IP+0qrdNT39lyqCic1TgYpSYPwRVk5lfYJDzeCXbIRjNUK9ahnmhG9FrMzIHT5u2
u4/kPLLI1jOp6EVVy+sdUxxySNBnzhM9ICppONcGNK4A8PuxM+sQk49LizpvvZhd
iF+dkYBkKNOG7/Xn7eY/IiSifYammgKONZgroX30EN6iETgusUcypBtSG5J8PgMf
htcEXUGWhyxH0PYQTUXVCaCrSkunP+yagK5/0/eYCoh7NzW9czhVW6lMFcz3Qs1w
jHY0SbTafJ7Thw/gUyTtr8qhxAE7aQ8ss3ViEvu/jvsqNxyf3LNF7iZEUwbuPdu0
MQTSyDwdiQsGB9VRPGqJ/+6x7oxdOuUSWloEo2EOsCAH1UslKQcNC1fsKCPzJIkt
0ox18yCthqoUqGl+h5BGh+jeLQgu3nRUcTomWrhOaFcMF5G7YK2pMmiNgAeiIo5i
Ng7RIlnvVJzqJSRokJX6vMUdqq87pNK8wt5PArA5tiYmCUf1rovo/FXtMd46SXYU
Af0g8HfreZdPHintFb4edjL4ZO6UqGVQtjSm/eo6GDnQPP8XHyCNdarEuyMLR51I
tVtwGKso37/l9nK5UpB1+iw+zCN9krUrSOYW3QTmhspy7pHKIKOIw1MCJFnuvE3b
UqfK7tfXECfBEEzdrLpqrySjxH+nVvoU3IozGcwghA+2ZDjfm7EvdPZi1h35Axol
sOT7PG0ZrPz56Nk8lK08Z/EZ/QG44TjY8FS3aYZ6fZL3Rt2LGf1+WFHzv79awUlo
NHRmmL+NvfjN2ld9nfcPqhYTqFcxLv4bQlZ/CIJbVOZ5PVx+VxuJoc36xyJcZj9d
9yFLqaB2VOGLPocy+42Cxj0AeH5mBm71XHm8WfgGCUNWC35f+cs0oMb6FWcQ25ZV
YRBLCId14f0aJBpV/Kwd9cVDyf7YcytFN2jVbA/WCjDUNfWEq0CbNfzeihMayFnm
NOl+1Kh6A9Ui+rQ8PzVnf0ZOJswWpR4FZ8AFchb1l+qphe4ueK/EiIRiqlGrJF7V
CHunpGMlyu7gH67SvuMug+4C8/20N+yNtTGT5pgiw92+3+6PP+xUGtmbWLb8tPkQ
f6ce2kDz4WTh6v8Jroco0nn2cEDp+izlL4u6wO6vvXGBnpf/DBsAEeCcjBsFl3e/
oZfnCITUNqVSwvUODCI3zgxEC257Xn29GeMipDHjVhyjXAT5ETrQc7NXnNNAvQtU
c2J6uFzf1kqE6529aCSoFQi4i7J6u5Zq0OrWDIUy9J9bEbBgtg3NpuziBk+BRcmM
JoAHO8AXsJesUK+rQp1hIFBpnlzhZ1M1SfnCZMteprxPrNo48oN7pes8iQEBkdSC
vUQvNDBBUZJ5VtGIn6Xn30XvBZhvKl3O4eLNX6X3NrIq1UMn19wFuG/TVm1LxO8w
xNJMkuaTZ7wUR7gd5SavkuXORna0nDwDalVwE1KfUFvgXBJD4P3HpWx/7zKWysfE
WmswdbIdGZoU7c4p8cZZpuNI+OYVohkM6Iqh5dKwNYhZzkAEcuWDgyGlPIaEY6Md
I5AOvsulaYoZnfFx38qGIvHt6ZYoXlPj6297Qh6W6o39Neerf+5bpjMJf2r2576m
hELebOdyyRTEL8pQRrCJZIPoHnoNgGAWPja5InRpGaW1RGOAgsJxM51i8Q8/wWJA
BGBVgkgQ6cORAtdG4AiA1AWoOzV8wI17hNm2HH6bFkaCjnUR8d0ie/WwV5KaSnEZ
eSPtHBXE+PJgwuzpKM7E0Lxy6ITwfL/52n4yhwRTfMZOIhClljr5vVix5ueq4dKb
zPkJuRH0kzuid7febr1Pu6JylL6wNVpBtNNrQFYlm63R6vysl7dRaZA75gySLCoZ
cb3OowaQIywfSXENhQWNAwWr56vp1UV9Eg52vWEibr5N5mYOPKDWUpTmlxEV/ESO
xylBQpgJt4xg37frrfECK0Q6YCUYE3ip/EJ8ALHDFPygbFNCHyDKQzhYdb4cvK0g
Vt33afoecjNLlxZAeCLki5D0EcqECO2ekJKSKj2ybP59ILR5NW2jNoz280ckKr5z
cph+RgA/CwrFxYzukkcwWeXzl9pkY17ocktDeW0paCkw1mlanWojioYG6sRjilKl
7O6fV7E49wkOK0/amr1O+IjJQ3fTmTFsoLyaS7NBkBpucYlvHzB9o+H2wj6Q9E9B
VAz9u1q/b4wjbkE9uA+jezCTQbhQTnlm8pWNeQt4V5eesK/2oimHJJeInQwvUH49
Dd2HNG/xBeLLnn6C3L0z1T8KKoYlfrkk2u6vL/oAdkbJdE8km9RUbqnPVs15FoPy
p4X60+wVr4I0fZTGa8kxDSJa9s7wNcO1DMplg3uyhDTy7xFNvw2ZZF3phaL3wJyQ
GkG1xqVeXQPnLKGwwoHRIL2s4+DDq8ebvik8+6IKZxW1ETHpWRZrOSlcEig5Pt+y
u0WI+0xc3Mi75YwX17e0p7h4s+1LSEeGahbu8zZQQncGcgTKButMThXcPkEZKfvs
4fGIazQH+E8nSrQT4X/z/enpod1Og2iuvt5gVYPG/AtSpQFeWk036YF7WVDfc5fd
AMESic87w9evubx/7fyj/An+98za2S07IppYYiw0c8RC7ufcNGUat29ObAvA0wJm
c9L6qx/mVAod+AJxSECyAZ6sLrwaRASVuElVFGccy6yI0XrNNugBU8ibW9MXhdI3
w1Q8rj4bTE2nqfRla5ml1517R5tlikntlpDW9GBT9uGiFUQimxc51lpB3J+z6Jcn
Rje2ancVIiGEn0mwryEySJcfEjD9nwgjUUjRAghvR2l5hF/1o4RoQ21el6m88czO
2hEHTPXlTd4d8TpJdnJugWYo6sVIRwAWYRq9SzBhyI9JJ++fSQ+EZtTzD+s093G+
3v5hyBJSX+Ox+wJ233UCRuNtOO49Zp2v0u/G56OmyObObRcGZWuY+s0sQ5p5+tAC
UO6Xh4n5MYmdmC4BVkQYWVEQSNbbbErt4cldtI2/CiIs88+PIauILJ5nHSBsA/bO
NR1OcZa2WYOIGJoPMfXzX3IDuCRaWUxGAQ9dRE4fy+xTuTLq1pr6pZRuCYie4NDL
vx7q5zQk0O730wh87xOV/erb/faUH90+6spGbJf2B67r760YSau57aUZm7D7gBUO
Hve78F9PmCQ/WA8DnPcPRDLlcPjjSpsQrOVJPVWkcZQwaZG2+6IRI1AReZw3F7Ep
8y6GtWu8tChBo/rxmdB7u5W793dpfxA8AnvIwSuyNbxEEAftSzyyiMMZT2yPg2tD
zHrInpireEa3AOjApWYd7Xnoqt2bN6aiJLJVu+520EfHQLTa4yPqmvXwlU7vuuVx
8F29IsARsTeCCa6CJQ4Iz9hkgaC6NlWxskI14CLElqpOknohwkIR/w+1/y+iPFC6
wdvFQUv9sNXnHcxX7e9hRKaTEp/5Zh32+beW9iiHOs4uEM3Ln0S93iRIx/yLxNST
2lteIr3uMJfCkOwF2ecbhxR9q2uvM9WNCvL2Q1oHNPYbqp/SMKjXT6L7iNyZWY0e
vt5pzOXue2vhWKrjY9bHn6MU20d0Pb6GAvvr23cov2yYbs9RlGFhFgOzqcWysial
6jWfo72JWM907/8FxrWWdMhv8K604poGOtiYCbRS357Rq2EVd/tW/OslBMtR5iHl
hoc4PyrjVUVpotFGnpLu2EHdZxl5kcBCXNBdQnlbR2+zoOfRY3b9lbDrVWTfDg2f
ZzHzwrx52Tjh8tJAJo94g2K/KfL26Zn4h0e9sGp8HTP7pMZ/CiZ3y1XlU/0rhVeF
BLRJmBmErFFJPeiAtfdD9Ze/QPaAcEO8ydR0agZssvjACrFIF0uLmX2JJhC9+6st
/G9KmjsvtJgAEJokFNgTSreXBYz+nmmKrY4glK+VwKtNzUJYOc1Fkw1LshtPxI3o
X8wgHwXzjeB1lr7ANUEuVEIXRuWVEgWUndU5L1FLUImfREYAdMSqiawHatZhjvWT
i/Q343+WbJwiSRXtPFEohjTqdPde7Hcr9GStytNCip7Kr0gnpBF32SCMaZ2KEeei
+CD0j79bfimNRwNvzbw3+VukzOFGW7SzchKNxTvD2PWcQMQklyEMk3FIQ4CTAyAv
iOTYA4gVmNgedOMX9o+ab6D237im4uG9WnlHJTlo2gR7PY/6QqstADKxAweux98y
GRrxdWNfHq58joNSCWEvzSHXHdBtmi3QPkzsOFAUx1bT+Ll/1wsxKmV5P1gDKrk4
o3+bTxFCxZLhatKLZHxTKwp0Ka/rZyyfkb1SecJRMaaYGdrTGN4QUvTCLM/PsFur
GvgnOohPLBXfBNQ1Wrll2bTnECH5bupdHONSnNoiNh1j/skzSdOq9Fx+UqdpebcC
vuM9qbzmDTFCN/FhNZLKrwvS6SN9Ou7sYPetDiiayyazI5VK3nxWuKDIjsDplNqf
nFQ3ZteJl3BP03ugiRXqkh9PidPZCBV+npINqJVcaUCikXZhj4n38KD1PVDXxj0C
4AlqGNkxa7qI3OHVdiE+yRCOoKqFhFw9XsMKrxOJ9V7NWoKN++bX3kv8r0dCNm78
9BoFrUWn/p7tC83qWtk+cSzgTyfpn0foo0bKbyShZvm4T7RdeLvZFtt8STS8UmTc
+wDTwdtP2pCZYX/duiYcvcy3wvtdUrCqWwy+v3sTQPviPOKH7911gdrkmu/fqiE2
pmC0jXgx3mJoBN0cx/sW2UmThG6YNFt7WuihvmlOw6lmbRs4308Wl8VHoGR7cKVS
b46y6cp+ZPzXYXyHbF9LTnlgZBvDyj0MZ8sBErBljH+2mfFS1F4nlYvD5r+OEPqF
HW1Otz0jbOadaptWT4BvNFv8GR5b06w9pT7OzdacV4xz7bNMqBuYxKBzUMbGRRyd
AP4P7Hs6yVkOWKdHP+20gP9eaWzl74xauDtE6asbcA9Z38PFwbcG5afraO5q6tYu
ASRSbhZtyGhFrhvCog7zHq59eEeFJWXCQThpkikHybOHtgNU6ZgxiO2FcmpYNO8Z
+88sRNPvExHKKxb3+DGjURMdw6ULueROGUlxU77+g1zpoHiGISaEEEmO2c/8PFv3
PB8dNC5RgZStRNc+HGS+756PTHu8pn+U9ZcWyK8yYAKX6GuqKU+DwnofRm49TEbJ
CCvVNj9aYSIhN+VKayfcZlPzpFtIczS6Ail+MoG6iTbpfR+x9F5ocfSfm1Incw6Q
JPVAuklNHYVtBMJHIMZZ6F/KXVsQQhbFp/+8WyH+lQaKTojkfQe+shKrQyGjaxIT
pjvGrF4BjHFobOEkNo1Owyiz/Aj67uB5bEEy2+UleFSYo091KYCeF8QNbzut/IaR
Bhd2+Q2UTgRqnzyFigLENluJNkBZkVQVUKciiS726vkuLLVAprIQWawzpywdOTZ1
MlqkPG+eCntBiFtG0T7dRzHvc2wHP1tIPxUteHkqJfg6Mk1IdppDkwnj3HKOpwrH
EUPMLJMFMuw9I+4RjvlPnJ+Et8FMOrydV9e2axaAbCKI3DdGpRJrQIaVUhH1GaKC
mlUY46DXKZAwIlf6FQd3y15a96kq0l+wyvH1IhLly1KpuoU7SPgYgGto6jNO3cKj
mIimyq4CUFWrNXz2Y8/3VGgyKUcsAicJvrhz06fdcmJk9GSBO+9XBeQkHQPjS64N
UPMOBUFoI/lIHAD81ozNMCvclpYrpTdUtnsffVM29wgufKC4IpzoOMsppuT5DM73
NvqGrkiCRNZNnD94iiB15D3hvxAxZE7yT4Fty3lLO44cKwZ1RxZwPPQRtXxi8YEo
cvZ2XE8gwgBd8pbjyEvkQcwl1RmDKjUr6CxQ3hlxT7nn/RoiYfIXer0FNX2awS61
KQ8Na6tOfFbL0SG7iicGYK5wpwR7oI9sL/+BUMyu0lUxe2SgFSKRj+1tPt2LLoX1
q1TZtORyQc7+wVBdgvq6BhH+b8Ne2jQWvNRjqCKzuaWLpHPk4/dUxxWHvdcNKmW0
VOb9bH33zr3lsmOONL3UmFabeu9P1ilrijzcn2qNDq58hr46vhzn1KzNhmUJGnC1
bYfsWcFmw41S6rcqeuWnJH4XsfAMyNem17Yfjqb14OW46kGmyK7+2k13KlieYmZn
l2pkfTbSNsJvrUn7dCeppzQB6FMUgbCORvRlclbY3qe3Hhk4OQvaNH3cA2fAR2y9
K15hgJBrdKG0byuGvHxxeAU0Swv21dS1Go51nv33ax+fPBm5jM9O+GTRo/gSY5ai
3yaiu+YGySziJNWxoqcccScH1WK3T0uzI49UxlLcwblv3rqJnS0imL3z6snn7ABW
6/3JEWOQlV3s9bPMg50rnErJeoTLfqNLmu9eFEEdJiS+92cVUdbiQkzVh4zQLU3f
pbAmiMMd4F/TEsl6CEOd2aJyBef+9hfcwB1rUPp8+v0wO+ZBPZ0GjkU8CnrAo4S3
yQ/aKqN/ETMJg4TimY9t9l/KtKBeWthvFx+yQKAMfx8JkJb3zeewg7IVwSbWJoZA
/WykddrOehVBEAxGIueB36geNeJcv4BOAjUGxrFtV+UcYIzNNN4WUTf5bX7TY92b
yRJa5ez0hUuSpojQ8HD4UiLp+3xLCvA1hcMmKRVfL4jNmwze+sckZH1xkrmU3Ddf
HqM2/4qI5oJAWQiDNztYX0OygzEuRIngRCpqQ9WP4Bz5vAyc6xWP3ouBXItkkVwV
2DNoDGbM/Z2prf6fyXmAqiDVQwHltWd+kn1CFF/J5QnQHt6Q/u+mslmM0A+DhYVk
c6AvoCTuR1FY9xVsGb5UhyPParMYUqwVdgRBkKY5X6l6xvnI3eH4QtIWXVgNFps7
5xmkI53q24hWH2ErKU3p8nNL6jlf0zWQDc60V0qtBinAqXMVAjSj9DK4uWyvepzN
ZOh0jZa/+cttwKX4qxjs0FoJuBRoUTQL9SOScU56VwL0fjSBYE2+locXuuyeMIln
CmLzxjOnqWAzS2HtnSljKN8pznAJn7PmDxBAfi8KAgBB0QzVxOyc+RsYBB7iHpTF
HcH+XVDQX5/ggXWe1WksleLtZ+lUl3DmB7jGmefDvEyfFy6ix+qpFvr/CtD0XaZa
LJGpvpYT9ShG26GCmSRWsjYs6VyXPvwyMGE4iQjeSKLbEJEcdjCRS4H2CrljfGZx
ZSUVBIhjxS+Ns7/jsfhB0bhM9MvZ0RelkppVHCsoOpyc9EQxGu9oOU5lnsbnHyVf
jNrD0EUEi15TgXfqIxe0Z5I55QLXOx08IW25ZHSSgl361W038rp7Pel+rsigKjw+
BJiKJC1uQbLApm/aLbGNG/JjAFXdbftEUmG4iKY4vufzF+45/L35xOwqqIPzzARA
frcSWKqA0raGLGYzJc1EPPEJZg3ip1B3RXHHVxhuokoqte1kLbgYNViau9zv5pLJ
cOW4M4FLuK5Dsw5GtvuwM0dIbmkeyGAtYlMoWN9FBISrY1e3vzisJFbd95kzv2NR
i0fDPNC83lGzr/2aa8OHdQK8YUGbi0gCf1wsuP3A1WVsTXRTR4a3yveLGxm3Xotg
mYHLfLQAQnFYxYb0b1Ctw+TBZ1YsiehxSA6z0DdPOMLErk32sst4EWbWX4KdrWgu
GQHdlJR1+YyNsiTW1248IZDN/ITkb66p/PC8hgI7ZkLRh5KOI29yrD3ZFKmDyRWE
Sef531Nb4bqHj0BbjCVIXxiGwVJDZcc7P8Qd/w1Bq5FY/AcGm09FG0O9Z0+qiguD
PT0u62XzZUC6S4myMqSPkK4LiIp9R+TUBCkWEaAOEa0YBDypUXdosgZwQCn5/XGo
qodGkV1m+MqqApd5Zlb3+2GZWFzo287Q+xiaUWnXws32MQHTda9Fm5bP+5JzlVeh
PDNi45eCSwpYaTRSn8x+aUac5gQtPvr+a8S/K8pOyx5PopiTTwEhkoK95FgM8opt
ALBqVFZYzxAtaMy4+otNDyjWT32tEebR9FFCVzb77BE9iEMkXvgvIFYDVPZWTyx3
LP1GzXwAoDnlUhOQtY+ERMpdM84tFCUEOZJ08yH51i7Jutc8tsZjtY4bLYT38jFo
+qXVUSfnknHqtsvfWfYMttJtLeBnCs0wCdPV3beSE2Pyalc9aYpZy7csFJHxc43M
5aLtEuUp5kuoXyqz7po6WFVbROMksxfyPsE8hHjpZfO0dT98q+lWPxLeCicdVJd1
0FnNjdaGQ4fF4DSOJoRBrbrOpzNHyUoUroil1DgFtsvZm88oF2JhIsGcZc1e6+ry
07yrcbWoDOelJIVSEld8thUDw9xHlZNdvdvhjGf4Az3SWEtJ+A22kj0pw5r8XrA0
2de5IZJl/zhLOleempp3nj07jQFJzgr7D9R7PzFoLvAkrJrljsZ3Pc0UTGI+WhE8
J20QTdxyF88nv5sOdjv8yvjwgvvygF3CwzMuRpkEMMQ9L6+H8q5oL33kW3UlzfUR
vGWGTRQ/D/3eO73kE7e2sjw2CC/21WjAPlklTnHBEFsI58iPBDNMtNfZTc3vm538
jJGjv/R+Zk2yfiGfsBjUXuJ6ysN7FlFfAp7Rjk/0FPXbsmBoKGvn9AzsuBV0YKUx
6EQu4Ix1ybkchy0Xa5AJRlOLY8E2L8smVzc54UPyFDIkHwO0eUzSykC/7OzLQnsV
drGU4GyiKcxmfUn8Ly8d34HnIal0zsX21dkDRV3Mx2js6hMGbK3mlIs0kN8UyFz3
HjFvWgF0uhN8dhPVhFUokgw271KNBgvqh7tKoGkPdZohcfux0cx2G8Rq6PiwIvI0
C7m5CgjrqOjZSavQa0YjMB/s2PCgThhI9Ur+6laU3l6yoUbmKl6lz/fBj1LZZQjv
wk90p9M73SOupNGTPZlRX5ra6ahW5biy+d22TS5tCpdWifxeyh5so15m+wlHqTjB
wOJDH0EJ9aHYLyy06cwxdHpQHylrUAThOF79ltleLANQ4qZyShupiQAzP8sbH+nH
PXcgbvX7Jpr7LbswS9U//9LjRZuVOusETit+LiVNKCYqF29LL6VNpOqBvpf4kmZs
UhtdZwojGD/zDXLJ3hIqtaLhowHGA0QpBuHekSW9OBZ7Ttw9FhzVQaFm5hAFjJLp
P6h5GQ6y4qufVylhJYkFv5sb/0z/7sksWzZCfz7Z//Nm1C6m/MJKFWvRCfF4aYet
UftLvfE2LwUztVHJSyX/X4AEtyOh6iYNAz97nFISrQW9BW9HhMwkMmMLzts0v71p
tCxgb6U+UTcwybaaGzkMRtwMWSs0VD1F/6SwGNyuBrfkB5GKUotmpKnyEdUs5+5Y
MdRSiOGHVibKMW6nRQlVdPOzl00ujqHvqyaxhBwX2a+k02Ztwc3Z+ziJC0FFtUDQ
ZDBrJ1I+ZQGzRmyyBOswJt2Nv4V1N9MZWHUSZ/zrMfi98/torH7y5LPc9Yp7LFZn
C2VFPoSW38ZsXThPwLsKLlc9qdZDj5x7Pv9pYUxurbSTqFX42q5MADeykoV0kUQX
1/45qcGd22BspEmdGbWHQHTmzzRnQjtzZvWRslNTBU+qvLRmSnJND70jh0tPxq+E
Adu8P7haLkJJkoQlVV06s4I/WJspZS7MfCAMZSjVrwStySR7R4q9tNWceK6SS+v9
agIRxDCZv9RQOd213dzch3iMylvSqBhm482bKYR5AgOrYvsHEI27WumLUPi+fmR5
Zq9IZKLwkNLvoUe0Il2XCmJAp1rxhANBJjQQ/+r+v3i6YHxEpHgIcYDL0WSecxyh
8/la+BeltXBRBtUJhlK0B5J11FO4GaSD1oZH9fMTfls1GYXjXHiOah+RWuSq3A++
t7KK2/NbfZ2b7rrWcxjewS/2xfIhACYB27tRiRqChjpOvcYU09l7qctPjKh6NPC/
MKf7gdFd2sCB2iGYp7kgEsY7JCtj4dUxTnhixDLthX9bNzI4S7M/8HpsKj87wkxo
oU7bnIGMjjYWEHUx7pxn1HbchLF3e3H4OYE4P9zf1q5LphumIRHO1+kjrRYUORxQ
KQmBbvbNcHJ57BTrGudvDuv/o+46MvO+ODm8dhpcf23stqo74SvmEtydQ+gz9Rev
hFCT+yDdf6fbbqMB9h1pgoHDANbD/DyIJuBNzxiZCrLiHu4yO7iGDwQc46hA9m6+
htO+6Rlx9vSozOqPY6Ei+9CD71NRyPTVDcLAm0qVP6kNq8aUa6wYqU4UeY+YiYi5
z0AOHVCp3B4xYUOnUUy7IK2f5vl2hUho6lYRqgx2YGMSz1ztv1vAS0c6nSyk0aFz
A1yHcJrokDj282dLYnheSiHR+Dnexw9V2qalWxxxJEziuMTV+Gi72k1+bYShjBUk
sbovCQ8+V0ecJtnlJKB3gubeyzQ8UNPQHKAWWclAfSEMwp//FQ+/ClXJlEqtbfQP
DDZe+fGXWxWacY2FjcaXMmR8oEwVAFOju2iCC4odSKErupaM+fkEjYa0nRejdk+y
OyeN7Tup00Y9aNvKpCU60wWNtcdGIBYiFilerN1O+FvPR3IMXtMpB72QdAefKMOf
fGdVTeu7VYWR+L37o3655No95DsFySVVZkhU5dzj+Z8Xa2lZajY04DjOZYQTLxHa
MJDjtk61fwVlCNhR53da4UNoQIsIlVlojuShUF166jItDvaPiqlHKtz9v8AnD+2X
tspbRAnVIiJ3JgtStiS8ABWww3e8bFbWzY0mq/Z6YHypDXAZyznu7u/PqRVnK4MT
Qi6zpxgrb1Iq9mtfmCQbJd57RLCT2eshsXEJ//1dqxqzDduxhZ5C0osysW4RyIx6
IfHM7hsb6uyy4PsPJn/idPJ1TJ5/JJx8PpZeY2/26SS8hdUakE1RlQrAzVlNIat/
WdD71BSPu9mzUYvqIoVQKQ31U02HbDcaDzDSg5AmU3Hf1TB+acuVaeVCofPXP7Qq
Y3TCYL4HNrL5IgzxNg/BMHUXT/cfaL/0MgfIXvFW1cCXv/GccaaGu11c2cERhFVw
aWxqv20Go/lSOSWIr+N6iOppZkQKm8NdatCOYPk4IzgxbGfa3hssP6le0XpYKdd7
5KrfdgVgY5r0yDgh3VZ1bWzdANXCUNhNu40yNel9Mo04i7W/XUxaFz7kF6/mJ362
jE6Wows1UgRPC61qqWRYt/t+yQjbDtaCv6rm40URHsUdassppmTkgnVe5wnHTUkR
DuB/UxbUztqiEL30lNeDBOOISjabgS1CYLEfGHvGuqpY3qWIzSfp3VUrpIIt8e7u
/XQPTUC/Ep6mhBGaHqs1zHq703s4Z8Bs+IcacK/RW/N6PdspxW9HujrKDaYIMIrL
hUs+kHPGsBV3zc/g/kDyIOx3bgXbIVDyI42nIqfZGMAfuwKgbqX0SHYIuKpTgTeA
4vFVX2KeUSDcgCl6thCQYeSelu77pF4fWNCORbqk5VJ916zgPrytZy6zmFYlAQmq
FgEgbGY2Xa+znVlUdlV9g2PiSDHwcfyV8/QBuMC4PREDwArOVRhU/ogzaxkUPkJB
l41dTKbIYXfi+rbhoZSEV59BWlEv3DsHurjVybaHdq/Ns6D7LNlWeFTUSsrWLVyd
s87TyZ3Zwn1G+AviJ7yv2fNfILbb9NR+dq4zcDUETmY6e5GUw2RMgTZ6LzriMqaF
GrLVFPvNapH8bIKtlt9GPQsTKq5RWKNUq/sW4BzT3QK52fU52lvdo3jeYBEkUaA6
/TGy/ODoD0WPNVRREvq9uydg7JUtiazT5nnAyhQvUQ04p//CDvylok+uZ3hf22Hu
rnHZRaPA8urvqyD1sBFBSpnbxOKqr/iRCzUTWA6YePNAuHOd7k9W9josiXoqQqi0
3HCJFx0mihkr6l3riKUrzGHQMFPeTdR91M6SASmw0F8TXWGvzZgTCscyoXm/56Ur
RqzF/+oY/6nZnmP3x1fpJbSheQuIzR0P9drZonEamEzoXDsDqphLRIqc5vwW65vr
qF4VdXbbi2LiFkxKQCdly1Oh2bNDjnWtMqM6q0Z9N0dn8O8bQmLYlMnGAnrhwx21
MOI/0rht9RMtg83g7ThEwJXfThWq7NmF5EEHXfSKG9q5s+pk78+aYrY7xMPfK/R1
RB1UghoU+u18szSCMneKwSwwee3KbAh5R0cgNN5JzoQM+iIKw3tBUX6X4C9kY6ld
X1OsQFUfhqv5b7PZamo2/HPhwvv4vmB2jdYtnTYwZCS5Vij7KGzt0hsGJIKmwOny
1qNiFUSUIJIZE2yFU/Qa+ToSj6RHavByflMJUYlX8fEfOV7IqLXBMd6ajRMr0yLU
SFWCSh6Q8k7WTIvY7iRj5dQscNF2PVXyXuk/Lszwi18du8MIudeSbiwyem0EfqjU
NS1WJ+v1fuhZfASJzWbQOd/HYEgDvi/S3x5Y9j1hvS5FLXup1F//3WAARoOSQhYr
1qd2409XdPmvSBcUquHEAlddRKSrc7XwRbE6cDaWewtkSomiUkZlY5zIfPFhv9BE
7D0o53CLMYH0ixwPrqud0WhENkovkZ52cbT955r27z+D6roO7YSSFmItO2GZjIfa
t24qUm9Rqvr3uUV1M27Uih65NBHkz/JEgZJOXOWVBpgWhVlVAH98AMkiaxgzWdl/
1MH2BoM4bq707UJv6rJ8tgnLSmtwf5MJZ+fA+tJbYctIuN6EbWVcVaIKaym1OZEB
5tF62CcFGUOaCoFf2YMhSTi9M+uml2n2FtB0eh+NRaKsX3ZjTievnAs5lymYa+Ty
QoKxu5Pkxh/KT0/ermyJDZtzQ/gUgp8AyheboEaOLiaXvoqrcW7DOdbDT7vAZxyN
sYzxiuOG/WeO2ogyEPAGfikJT4QSpP/PW/Jn1HpwcI0yjydI5nb80N6bG/R/9TIO
K2bQ//xnpWyYRRcmDrM3E/39OAoYmXyRSIQc0muSedIybuTFa8ax8cAbojRRCZ37
FJK6ssa3lAI27iM31eWeaZ9xg/teXaeg0YnnciwMlYUkbwfgA5yenDcZDD/mcYPP
B8u92XarScQrLAcTggc3DVVOVyGpY62GSE2vCbdsI0e4I62av/K/GTqton5WK8f3
dms+Fj9Z8H3f8jc3xeF+8NH/0gi/2JneUBRLcjT/vd2lpAHpGXBvJG6x65ocs9c3
ifl2URO6MAszWOJII3CWeeP7vugzhHiPVFtc/HLidyEQ0UTYXqeiaEz9y4uTwgun
mfslFKJF5FHKqG42HmyThPLR4Vem7f1qofegbOsrwv6GONZWsB3n4CKbAZPkRqPC
zkYaZzFtGfIFfFjjiwB6IuCUslC9h05XJ3TrK1+BUSruwiMx0c9BhG2a9zBMoBas
hrv3Bx7awimBr11v8vWmV0nH9Wxxj3BUyUn2HK66uCxXJMnkIscqFHarODkIr0fc
t5m5ehLA/OCrIwdSaVhf1dBR2ev8Fr2sP7XuWRvcprpA5jduM+ADqEAE7XnEOuZT
b09U6aVe46qfmok+eqk13TBNS10+oG/v9hOo/SQmDcLQryUftAnWEAEyyRFLYKHv
IDbLgykZ62vJEOPNFXitVHBc2nnOqYPqueNU5vXvxiSLSWV2ko6F0TgA4eoZA+Dl
tplZ/nniMnO5nY46KIwI2kujC00xeucsWwM0yBzyQLLFoD2ocL5DB4Bv85fleU/K
RSefQGmjInHyoQl5nckv54es8MO6Uw+h4n/QdRRy9ia0aK/6Osvw0Zqyu8bkFVC2
xY8n9fGWCRcCoRqibZNaqS3FRIlfh2/wd1lEqkMkbYK3/CMRDnSMzHtVrkPYAM0y
nxUhHKizsH3FZHFn1tAu9EWeflz/6iQxKS2qMSeWpTD8jFdPV95xjREvSJevzRg2
nlaKLK2FPzBCuvhcYGyWcMNs5AL8m+0sQe7TPBh/xRIRqQy1Nq00jWBwml4k8l8/
//dt9qrmz9d7+eoJMHWRKfYxA6swfzTqJFz3AH8N63Z5S3FcVEAd6oz8wm0laW3v
7vxynkBQcWDD5vxlhTFm8Z0TrJC310aDgSWQePtf6FWVgcB2Bs2w0kwOpcIophe6
/Ea5svo0/xBGV5ps7vIUwie77Dn2CcXxB77EU96xRQYXliImfGscQ3Uq4yo+V2e0
81KeuzCssZ1lPlqI4D2Be9weQHeINEReyZB9FETH0RdzR49SpUtXSRM+Avx21AKH
5VDgIpOClLNkOChXEDCTAWRWMCgVs/QlDs7E5YcPYJaN5LQnoPZ5MIx31eH98OAb
vUh1zi8l7M5soapPDyyzOj7sTdVpJohyBZb+ST2XABvLpaz/GvqInh3Yhwr5q6ug
HfstMDWFWl8/I8RPwVZ0KYAsPO62aYJrzzvNr2YyxBJD8u58zYHWJm9kEhBSnCLi
t3mJI0j7yFBZ7Nk6UdZbJW/01ENkwSFAT5G9kCPfvhjZnFRb8zZx9rBE5POAGdu8
LArK5MlNsCpWleYwPWOYPt2hUFixkn/iXT8xfDi6gWPXJGghndmDU5idw163lKtN
jcu3/YrNPc/w+dU7ZgBMPFxbL8EHPnpjySuxVh/L1Gws2JBisX+JsFGsCOTFihtO
AATPUKkGTaikfqq0O5IbeXZLAdB3ItryUK7t+koEdwaoXq+h20H3/QsbQe/5HMkM
Z73wqiiSqoZwQNC0tTdCT3zm0i9/9ZjyJQc/UNAXaRdBi2IsuWkFm3RvDJIKOAaJ
Cxhs6FnNl8vFMcS7Qlr2ex3YiXn1sutO8IMVscR6TEgLoQ0F61eh9YN5emN/rLqt
rrqXGB2HW+aIQo3IGQXyBhxIEtCIAgkUl7WNCL0IBS9MpcbW9QhEP4pLl3CAgvUg
Yjd8Ub3YVzE6ZOoAyzfPQl2ZhSZsrbKAYIBRNdLv23+98DECioo0LVb5DOxAs6up
2IV7LUWrLgqc3zPPrqEiAY4exAbDozaBuwkFgrSSt0i6UzMjrlWkaLW2rFE59qV7
2mf0ca14WyPuFR7a7Jy0qkyVQZas5co+deHguyjKhS9FzvM+Z8bRcOsTqHvQVIoQ
6hv5EFJGqEVnoC6nBpJn4ShCfphvN/hOC9et7ehdyq5V1O70dR1I80ZH+rmEkNcS
jewIE4NbtkategpWjFLNFFe+fbH3Zp+ksSo8vtYSfOgACSVRnM7Vv+KpQMVBRyCl
epg8lx3bJaDEC2qZ6vzDsf533AMrD8FHNs1sIhqFstO9kmtdlnP450dMoXLJVzUb
XZumtQ4bUS7HmK0PWK7bEs/NCCoPVbT1khWhV/hSzAwu1mSBRuYt/eo+L5S5Bc7t
jqlCQaVhm6fUYjDfCT9+BarIIp0fgBn32FhFTkWSXperbprBI0+w6pZYiOq0gqUS
FvGBR/18rMTlrX+N3GY4k9jN4iyUVog5u+cf1p2uIq0xXiwDdlWKwzfd4SoJWY/6
5Fb8C/xXpwYSXgL3GFOq+cvWoELXDOSgKKR7cBKMrq7alUhftUccmgZ0fKn7TIZB
MYTwzkzbwEntz1VxlAs1LKgBi8uE2KhxvAIhaGX/HwcaEaW5LT+CPH9Qf/HrnOI+
0zLEarmY6WJbbS66QYIm0/jpJqSQB+yFsZCk84rQeZQ0JGf5M6Zw8jOv7Jb5ogJW
/nv06ieDxLKzeqiDHx6A1uP2GsdwWFG7oau8fhp5k2WY1da/fA/0TrD7aeIKxl33
tO6PLrDyesE+aCqlYFdcvMfOPDn9xMRKVsSxo8+CiMlKLT6jdBpm6gHbxVH2Hn4M
ePmibv/E9DeZtvNvEF6YhtnqbQ2Y0EkMP5VW1Us8lJ0LwBjAC+plorGD6qxuY9QQ
1Rbm2hZqASCuEo//jNxivT7Fz5YRGnOYA2Ax/ulzB+FBoqlPdVChwMWCFDU/AU/P
7exikj6vq0BxNwHxzmaVws5QiBDjkWhZ15bx82NQkXQbeN2CB5rz2/qp7aCXbiVT
PMAgVck3oBbnporYmrTwQxuTOLs41guDhpBgFVxNxGSXRwt40nQfp+pXLHhaCdk9
HJZ3o+U3Z7dNL71BvduFHCDyiLoyvqgJaVFlmbk2tLEVvmEN80UlWh6XL4e6ToYA
z2vS1MaDR8pB6LT4lUW46VfSLE3hiZ7MGjq/mbH3iGauB4z6KDc69VDe0fQeOQdF
eR+UJsmZ9PT/KqXYZC69W76D1smZPjCVj4zlM/HX0FO5TYKTkKCkDsIlfSVdQH76
SE9SYL5cQ+w4tqr6nJFTE5saufvXZWqciNPJA7+chnsj8NZVJiaC8rBAcZx7x09n
SHwP5kX0VyPyAb4l4ejKkxjuJcSuSNJ9+T4pXB71gfLiBJH6Wdr7U2+kanvn1J3h
k8HPOU+wSCkjaPXAPhn9qHd7DqP7G5E2fz2igTbrGucMyv8kmozdo6DkNbhhL85K
G4SUBcYXO7UI4vW5o5sYuo1qI+LLkUW6911VIxjy3YyatcpUiptvanC34Aboe7NW
gceeTEZMZ9sm3oJQlJ70ZmsongUEc9uIytK8RYQJOl080C0+ZFvmStHGCfit3WnH
T3kIsTo3cv3KZnlfQbbNDeIkbTTcKUq5/w7QbeNtloXckecw2W9/Hq7ESp9EGOmb
S2i8722z8hHeb5vpyd0L1QeiZTXcwSJSYCG8/E3GlwmNKOCKbzlzO6gnFTIMTXAs
3HjvooLxDpWwCdIBO2iVhLKXiTYNn2t3Vz2mQ2r1r+LlBa1MfXTCe2rjsYPEsvMu
u4ec+Rf5ySoVbnb28GlWiuIqi4eg5osO/UIbEnfVnBSNMZuTQImgsAsMojrDk3WC
3g0Ld6x53uIz3avJRUj1t67N9zVVFxyQJEjm5ZQApN9aUNKromRQvt8wkpQPYm1Y
dHwMjlNG2cZgFAhvBPH4kxsk9Wc7RnChX8mheTOjRELbA7ICZx/ngJPFgwKt0+vk
zXuDuBbnZqtiUR/urzSyDn215TfSGpDP3kuq15J5beuOvHNcOKPeP1+eUIfjhoSG
WPFYpNTLIccHhi9UVlvnO2OrU2rF5Y47S1MXo+ZfEM1HGKbrNWKbcYzDZe4IEzev
OSwtMUoiKS+xuMG1QArvV51tUgI6884cIKUGacUYEePBnPxQ90t3iHsBmru8cLtt
QdfP+TSG8/1uru2aj7VDyVkXkYamjIln0e2ejfCPe8DD2Md63Xenf6ZsyDhWHI/H
X7oU4YMPhBcAM5PWfBFb8vTrWxogGiJSOOb+OVeTNUIZAFTWVev0KNxD9bwZk5Oj
oYcZSP4vLgtNzawmuZX9b4Os+hW9oldPycV9BXqAKR/gxjfj6UA8BGWASQkTgaXn
BPUeM7xJab/UwIgNRhk86fYqRvdLcwo4Jf6fVj4mPKcmaAQEsyvn2yGHPP/XR7kF
X/CC+Nc66YLjqCdv5UTcaFvndMmoaYR0yDROJTEQ8RJXseiCRNAM2rDY8G7/FKzy
3h6XxGrBIrEPdxF2m40eIb+yMKuI/DEGxoynbuZXkWxtcpF299Oyq3NqPe9Xz3h9
8A6i3k0SVylg4CkWiRXIcM3p8r/gVsCyBizprBRPsXM5H55BKXcsRgmlp1H2G5AW
P8VELyJkJr18zazc7kIoN6sxHzRN2W5mai58IBzyeO8pI4XyXEOft+5W/sAR2H6q
z+uE6N8u7VE4o8z235SKwQM8U2NLiKCkjCdN/gwFlIfxQfTWsQIMTuPwaW2OBSM/
NIpXdZWwxwCqARs7+JrDBZ2m7ULWD8SIRZr8g72ITzHCCNY1wV3c7B1BBrON8VM8
jL2dXp3nyXQg6cYCGDKLF8dtqbMy7fp+bif43ZP5imDnvyQYhLsTFb+8LoOTc8DB
EmF+a0XCYxcHshJtZGfQjzz+M0cVn3/WvY2iIYXBIw50MEK7udKRUiGrQnYrfUvT
c2BmyEpLdZMFHWLLmkxH9k94FeZTfON0roXE7raI1mi8dtfYsxmZBGwloIZBLMUk
u7lg+NYlEk7B5ySz6qwVRW9bNUaRTHQc/guIF+JFsaWu8uDF1XZjE2avbovFwwV6
RmvcReqUU8VUpfsSevIghfOiip0elyEWtFta2yyKzPB6ce0ZhFeBEHeB9gzpItxS
heySR7M3/uIvChXlR4FC38fS/VeoQIVrYuQEwTtym8U1IS009ZdyyHwVUH4frmLv
1dvbkEDksRzWW4/rS2QC9b+N/I4gem3XxNZIfbiRJf8bUwlBYYHPzj4vLxhh/oQ+
M4jCb62nh3UzetDzB8jW8bDbpO6KWF142Ex/k8vH6jV8kXaiCbnqQ8z6ZcLqRx+N
AaymGrr2K7bWhOSoDEw4LJ0+wcc3rBYVs0GJddS5yabR8Z9c8yLHtUKpaIhp10z4
2buQcML+/WFI9Jo7GYX6JKf4CFGA6OhWcF87HjR5AbA8sB2M5KirwuyjZnCd27HY
7QxhUEPE36maXYj//XvjAmsxyYU4Qy0eji6o1H7N+irarWDRPL64Zeps2SO3mmL3
VYhgsi5H1vhZueblb1+gu43GPZiwfi44aB+8xnj4p6VbGiF+O0Hf5UR1I4+mNRRw
8sXIipDcdIVG3rTpEuNJhDUzNRhWir3OxOxPoKyJqUE39bch4DD6oHbwP3G+msu1
JGPoqnnV3Id6X6RG4qU0LBK5yOTyQQDHvbiISWYPSa1ATQWUsCAWncUStxtZ31A7
kA9w6krkJBIl7n8LUuwjC2jj+K7m3axkCa5b8Tb6UPN5BYpRy42/dEVpgJo737zn
8IouF6y2V6XU9aKz5HhlkFIsDTmwhW2F6GZI3exuk5HbSUwLeuDDqXDww9czodUb
bnhjWgdy/ZArBmwAia+yv76cxe//n+vuQcMvfsD4HT9pEc4WqPXWXYQpndIWWveo
tAtEimpnOk6zhUuh7/pq7jpTWA52duG5/qc2VSJ1poZ3ZzUguIp3C+rtvrzQ9cFe
zL2Ic7+Lz58t0+U8z1eVAbe67768Lh7uPukzk1rOHjPjQMRh7yUJ0zbsE6m6G4wA
zrwVoSzMjQ1dR3oe+KlPzobSHHtt1aHm7tFTVADIx4KxG1yO3QuSvZa6MliBMed6
8gsHJkCPr4f0dOgu8KWt1JcRfvjWNw6gp4vdlwSU3xtWXgg5TzPgxV+sRlGYCDel
6fh10LdHpsw7tjuUjXSO5xEENi+wmbp01b/z/CW+Y1veLqZNEjKAG72yrxqlJgGi
qhpUQ9Nf1nu2MlU1qsKc32GnxJXmn66Pg+9fCVQizISzYBCetkmHfMx5YQzHE/7D
bCzMXl6FOrR7i7Zv6o9m5hnBf94CY27V75QR1v6nSbr5Cse48ZxAoBE0FYseIZ5l
LrAs1WONyztRdyeolpjrMH9AR4QmTyXNoNUFExTNYluvD/6iELaB1IdfbS6VEX3g
bnY/TemawGxn10ie7YU3qJZE2uuI6rN4mMn5RP3JVQBoFYs8OgbGKJwGIXG/CWJD
/AhAkgoQfNjbYOoD3Cx+uqbjpN5sq6Q9rtkZmSDUvuvbWfG62EXKmemiqrvj5NGg
6fHMCwmwgCKWQJtbH1E8lErWCgQAH8VwqHbQs8EetAnX3mj8nwE5p9noKUnc7W0D
SCp/W1sGdB0D4uRramE6WE1yzj1s8s2tFvWmI1eky14MYBQLBGBCZOCLqUWme7p0
zosQQ8IyzdaC9nXcSyk0m04hwcQtK4ISt6CfM+sE0bNPyWycNiD3fbxxspSSPz6G
9RL+se7WgLkpfOzuf6P1Tzoe4FHYPRvVtPu8KfIoG/xJVczLwWtUubnQtQAbllz7
SNhFxFrZd2GvdoSrbjo9elp7ksUYpS//34r0ZRPfEZBNlbc/TfqzUU0+gGhuo2q4
C/CGA3V+9YeCmWDPBo1EaXQvQMrMVEqFRjVI6P4PqS7m5Fkzjix3bqrh8+Ooe/+B
dz3M1IbnVS/JnKCjIMo7z8JL4e8jcW0ttFHvdANTQiy6lEIjrXOHIqJPS8fFEX3z
FUPfCSusDEyN8P2YX0g9tC4+Pdo2PO9sfs1iF6lUzbLrZtvDmK73EKFPbRXqXTyd
JNnRihEI0XQgon5+rdosVtmCREsmk5rRyRJrxzuUR0mfDSGpisYIUIpZnBXWvQ49
6T6Z9OLDZh/Xf+lqpgyWlmBH6+Z/8IJv4hVch/abzkwPkCpcafq8V/l6uEnh3dIf
OPdkKSbJnunjSIZn1UWW9hHPEwhM3U3CTpQ3dK5CGP/b+xprxQcp+7jwCcHYGGfj
clfKVuyQWx9xeVMbzNuY1BNhAbRLyH68u4dO4q7sNIOd5go2V24F2DyKdrK5Y37M
CQExwIr2gTzHpQwHGQmy8UsRUbPDoSxQxKE6naDVGMLC3eU9acTRR5u/Hqe0pOjh
9DPAYmflZlB3PKqlCtOu5YiQkRbGoKkBopXi0u21tRc29Kr1fAC8iJsBQGs7UicA
byI0Y4arzdjvQ9RM5YbMBIHJ85xoOksmcKiTtoF3vJCueCgjkdiRvsTLKJuH6JKu
VDun+izsiSr3eVMMNh0qSzTUrFmNFhgH+1qzH/xFKnWFPhZMyKCl8SMCGrajWWne
DJhGw8xaCocwaegaq8dwz6fKYuHW0c32aDhgzaxP9ZVRJddrpsgfbyGk3z0cJ5xe
RQhlBbhqVgxTFuwhQPv2K3IeQjMKWMnWSDMjgmmQIPQKVEYP6NIM5BA/R3MC3k4y
nhLmc32OKywVOrHOs87QnxblSvEq6PjSkn+r2H5UXgHtx0eMJe+e7xuTrMwh56oc
lwWHkWuplsa/1HD0pjcR577fGYQ05ew+Un2YmKkpK/quSg6eZEE3C/DSeuotUGHV
a53EmMcUuPvEjtaxyZozDpjN02yoX9hXB+btNezHQEnrYN6GYz5QVdoRZpPOhB18
yyYJIq4DExYvfBTLUMSEgNIs1B7PWFUyoY4ZQLMelUhCOia8/WHduLj21pUjUkAh
Rlizftw3hzKgICK6GjYPtltQO8NjlCRy5yjnIUhHb487WnuDqOuRsik75zY8fjA4
rGHspwbmg4Fl3cz5qybLkONPIcxy/gP+zHiVFVQ7C7Lcy/dsiyQ4IAwVQy4EsNBs
ieng6SHh5cVrF0xqA3ESxZHaH0lCw5zop3vPnpjN0H1sUKzvtnnskdcWFSn4dmNV
4Dm6pUcXH9MKy2ta3/U7+VUU3Zp8gBSql/7wG27Tf9iwYMlg7DdbeB+V09DgStP6
aokEEDwjiJhOi1/9SBCllQpuyOBv41PCV9i2dS6jkv9mUANk6tEv8fUahB1rDrrW
pk+q7VTPPzIYxDRqaNeTaMML5hkw7Yn2ZqRHshoqCk2SPdufUe5haFx/WJBR/NKI
D2Dausq9HIXZemoZ8lbtDEjB2bJtgLy7k3IjUYWi4Om4d0VvcChPS30kvOZfqrHA
wmb7C+Wy0CcQQuKVxK88b3Jd44R6NL0R85nxqGHLMtxk1+1Co0FA0CDaCNfWg6pN
8ubGVV4H4gCZLyH/iKSp9rq7un9LhM3iD1jKseSgx0aKVOtaM3NtAOBaaU//B96J
4gCWihdmCdMi2Tj3nkWW4yN5mWW+D6voNkO0C6XGtAfL4Xu09iQ/yrvv3KfrT5EH
ELjbvIbQqw0zQZUTaIueW3YYd8njJpC9ao86CVP5UMpU0r78CeqtG01Jn5KPOi+k
GXnn6/4XokIPKpd1l4tLehdubiHLkROZNcwTJauOke/NkU9SyhXAdjIb9Hrzbeq+
NM70LVTxEInhX/i+Ik5PXtgZ2OpqtyzYM+TqWCJ7HXGPu7hNsQSLbf9F8OsbMIsF
RHGsZfoN4TT7GWdXV2UPXYfXcatVeBQ6KylvP6Sp64+V2LesVKlFyfTLLcjgPHeh
Cfom4KUKPHJ1rxeoTnu7+KFo6BOs7BlisKv9g3elLm6Tni9BDt1NGr/JWYztfH7P
ty8pIH/wCpxUYPmcLn1RGp1RVP8+HzTyA1XhyW23RYu4tJGbBnJb0SE7XT5PkVLc
naxylGsVRdY2nNEux10RdyP897fRQkR0AbT9PRnGdTc0nk7Si+qr+BIps06txoZ6
YD6TPnwUC1JzAxBZqwHgerC+uRt2W4gK3p5kVRp0zJUnpjgY23xqS+eEb2/9HjS0
EEFYhF9kJrdKx5v67VPYgKoF7br/xzpBoS4usFk/UPtBMY9iPJrHg6x7dMoDnu5g
/1x2+mlhTf9dDU0Jt0Kq5ZGkFKYQHw4tKay/Jj6mUZgBVrV3kt7QWfSwIGys/Fwl
tHnwRSFOZ/KOlkgITJzxyMtLMyEJAszDnefqRK8ZVlfRYbAEjYajHtYqoJWR9o6H
bg2sS06JdFpWS7zEGE19DoRser7XYR5C8evoqOxMsBR5tVchBwUi38PlfwMQJfLW
F9ROFLayxIQDl5Py8pyNMXkOjm8VcvrIFVnniZUlWv8DHIMwaILXnBqDVZven761
IHiMA1nwSpfDH2KWg9ZR71qctG1GQ/hNN9Vs1SSRZ5gOE29ah94Dyre8wksEMCuV
hdg+6xdQVeNoeLFnTSB6Jc2XsdxHwLv3UgHU+ii4dHqMv8KDUthAc98qaP1rRtb1
H2Vp9zyESrKXe+0dm0fVhLgc3YATUfuQo/xNMxTsDRgU8uPN1yXPCInVlKy7krkd
FzMwoIzMXxa2pgoQpAO3qoReVmR5VsqZ9QguKrS+3mMv+Y0r+30cO3lvn/lXpZJe
2yv5CqNqoXyb561wcIwaXuHR07ZGLER6Fc0bbYzBszGB44y4c+CFAHBYqNKEsSEg
FEqPKBqTun7+3Y7vgpklp4fSZvYrOcRg5MhRRK27lRR5nAidrVKueNq1ZX8m2mfl
AjtJORe6nZpo39lYapZwYcJjSbSjWYnQghS+KGRtLodQvARARMSvdM3YfDJ1yS+t
baHKieLwnEpU6v59ul8QEGObzTnYfbSppL5DAEkzv0VXQj5m89j9LiNt/JKdj2iB
i9ts4NU7x2AkqKcMyEdgV7dKdNOEDKMqncNeLYau0hF/eZFtFOBiwJ5TNd6UTlUv
D34/R8R8DU1riUT2Kfz8m/wn6/LZXCDCMgSQuOU9+UmCeS9H5L6/BVfklFFKd85j
AbgzmeNdnWFF8YsQKaZAnvUifs2LuW6llrTdVG8Y3EU7Mk9mL+2m8mTXwq8VHG8z
uRA7Ni74Zucnzb+B+Npf9j0J+Lp5TTPwmVwKO0DmP1R5tWyyPW14GtPfBSvc3fQV
ReQ8+FlZi5OJyfk7IH816i0GBXbSbTwMIaelzQRu7+pJoHuHqnEWnwmHXacujWpl
u47sBBIc+MJg+LDOa21hw2Q+a4ikRjS+djYNMFRW24QJmadH2jXNiMZcBp5oMRYB
/cBi7TFskHz2ZWqSACMuYDIZV9szjhAeQj7NY9Q0vjb0cfhTcE1mOfB3QrT5luTE
ObxrQV/UxceGvnY3qlTyRWWlWhbBiaRv5kYKN2OaUfHRK5rWE+Astw4TqZme9qEp
hH5M8jwPhQDX/O0lpI7Qd6FNVYtsM+y3voLfoCFLzZMU4PV/s9EZ+jLEeQJLXfEw
IAtKJ0yOq00nQieibvQKNLj9KUxY/1o3klyOEkjFTQeASrYaW+bY/easAhottLDY
6QBmnBXcY/ocC4P13K+byEHQ/0vui4P+FZ8FalFnsU39kCNhYxoxAwrVAZGxOFo+
GEILLtqm1S/7zpusrnanhTEEotynYlPdeXxQXy+b+cYDn+OZosRxUAAm9C245JM3
X9wp3O3CkPWL/KLBlmkGRPoM7bGSqVjouutNNzFo0otgfznRmCDE6hxWFL1F0R4z
z+s3hGgerM7FO8CRfQMn8DW+UWru2tadMA3kb3ujO98/WUGSfW8RtFNp/S+qWypL
w5rH3bJH9GRk1//8yMP+JSIrUwfOba7FdKoQmlA414Z7LU8cttRv5t3j/upZflm4
MDAyysi7Pya6alThrRwGkBOU/rzBtIKD0fvWRTV5EH06swQ6dnTu+TZ0QjvW9j9u
rsx4yD4wGOH01sYV5zs/EqcJKJu7/utviLycytZFhqItT/gDwkXRSp4VGlwRwW1F
dLn6jpBUo9lk3/qr2uEXbgLUb7XskQIGdjQYsPOEWhYQc18FsbwA3kHGRGvnAKps
hWwe2BQ8TQQI6KrRQcI+NuuVUisgBVse6AlUTqLSmMTc5HsnsVUrp1NDxqVvZDtE
zHrqtk2HEM5uZl0DWn0bczo8U9yv3Ja+aYCuSE4N1bx+VRfLEpCha1KIpEnrY0bb
3Kd5TcceA5tcXKUsFxVUhgguerLkmNWyy7dUYQ0U6cIuo8PC6Iuv71DgwHxeysEy
sMpUimjHYmbys93MchUVpc+A3fwxZwSg+rgykzD+yPOayo2mhsK7FW+3FpHpFmDq
9+pmHcjNM80/W2f0GK543VAN0PJo/fJM9YDtIH1ly6YGusrbtFDJUFWcdFK+gs7I
An4Fb0U69OMpi6GyY99hx773Yho5Baw8QlQdPnRckJ0tdlgRwGbYDImBPH01PaVi
iABIYWK5QRdLdvmkc04dRYTO3L83zlOfB2Q2Z8pfIa7PTWfCJUXSUeVWi8rf3WZQ
EtC8i5i4hY7hJCL0iMOFxdgkOCfRN26IZ+nf+YajWsjzO4FaFp0lvK01hqVMhzmY
+8jzEV/ke8zyJfKYNR42WKq13sa824Nw+KESh9gelGC86QnMFXjkXGRSl6qL3ycJ
qlKcKPw3BvZbUdty25RUDgqhNXurkxsx59oRZ3UtAXsFGOIILA4LowFOrAojzL0B
KF2VPg9TQUvDDkjN1/ty5w6qH7OPGccMoHXdKx+wdEzWyWzMN7rXv2cap/+7fbq4
1xz5gJBLfAu6vAX4eM/N+4yyqoThqhpue0Iq5XFn0rY9UywM+9yXEUfJ8JF/xIUS
GHZFvl56Jik2fxLht/Xrcj7QqGwgoJSCnIKmOJcyaFCFl5uM3nBzwAZZTVthfbDn
jBKqRm4/msVrpr+g1xIYNxoU9g44+u3hcrd38HRNJ2Z4kegQoyzP6QoGTy7Uqi6w
SEu3VwsQXdKl6Zxxyd4DPBJcUpQk1WDoyQIZMwoLF/fFOX0MGhoJQp1kqw/CwEQM
fi4hs9FBJFFlCY6ckFpfYQGbUDxEJ+9zGD8bSoESXs74z7BbYoqwNYGin9Kj4AjF
HouXoEk9JcSG/PH5Bhsy2n3XIU70CGhQDScgXBKi9FUdff1QX8GzCUq3IAm4fnYF
ZfphSelLWZXM5B9PLfD8fVeS7aj7+pVMT9I+DX0j6yuw8ML7OdXxybAaMAIN9MAH
SrKjWA9A7sHQy0sOb9wr7VAXdv70zbqOWDuopH8mCKWSOZ3y0oTAjcCfE5oWvNlu
PzQl5jvcojRWhF5ZBB6rBVGM1dRLSlwFSxORovclsPFePNVrzOvhq84iNSynA61b
ce4QMaNsovmq45BLge61HqSaFpck0IuYCljlIaz9oMtEvo8qFOXNGwSrhhGlJlSH
VgpvGltyUdNGjZFGheeB0NDyVPWFEX+0PE9YWVSdVoR+kn0ox+9qf/5hF5MTpl8b
IZqmu8Zz2TPK0KdRLHBq7Ag/3XbaWDx8uwnxOlh9W1Lf/Qma0psEtUKwdPMsqg9g
v1SFqARHtQuNdowXXWT5bbLkFdgPkNudGJUpB4mu14KzwFkaPe1Zl66kulIFt02S
dyP/y0k90ktewCCZyJYDkEnTBAP17RTkZ7YV2LG3FnnZ2kYhypMJV4L9EuueReau
+dQHFsU1EP011heuvgdTXwuiy2SrRalqHpHcU9hISs7Fb6MsgLlttd98rhw1VCRv
sVMEeEC81FPFzqkSPJISY1JxQDdPdasP+pen1F74I3vqbiQ2D8oei7fIWg3w4iTB
lb1SrDPAtzmiAC3OAl/VGY/DomN7XujANBt0dbBb1ZlIUK7GdG3vhq6sXGpufOos
piRkfZaYEsCOXj7qCYRURzVmOdERlkqFvKVkrueoAk7LgrFKbhKykheuPLZYNZju
kzHzgviAK/K5H+1x3XxcpLWnnoIyvNx3bF7FjM60Q85a1EATHp/NvR0ssVB4ipCY
pNb2dIkwxxuEzfrK2UCt6g6BpLA2IPxMI3svM20igUkwg060uZhQEx1kS/LkRhai
BflJ6MeGXPJWCYELtpBUdHK89dE5Yyjs1BfmDQghN5xQ4heFLfxmnWGL3nxGSBkE
kmGwG0aSc2kQIIscD8eGiXXTUv4WqulEWFi9PVC2eYZuSU/waU92lSODstuKZ6hS
1dN5byoXKMEr+bB85oM2eM/dOLO/szgcx9kyIfcNf0sxEPpltElIGwfuYFlE4Z2I
wlGb0KZJ/U6yFTBB73kDG4yZWzhuj+O3maBtqSade5rvLbqqx4Ib56Jp3+6BMR/o
UaQfV38E8R2GDfq6RdY7HYlwoVFJMNf7SKWDmf9XHLbJEy+hIalrKPv388XRsqwp
+BG33uaSs2+GsZYF999d4ZWMWWncSl0I+3U0VmSZ2b9vby0MtB7RKgt0sixfA5SR
iuBCpY65BWACr61tt5zZDKmFxtw8f+1Je4UxF/TK0nKmT0hCyhA3d3S7GNFQkURe
NSH25jUoM0x9BiR2dM+NpvnhgS0H3oS7uW06Ora0PhQimD4u/IxXTFFXvth6VPSY
CFAsJMT5dkORnOGUJxxLXHULAoR0I6diFUCpinB7DfpXxnitMTx5MTbExpj24r3m
bBlXtODs/6mXSSOTLgeaZ1HZcZRXv8FqHTHj7oUVEXgFonQb5QCy5ySxdmk+9rQ9
Ohai2qShnOQKHEQA/wIRYLAFKKH0oEvfTRSPn/yPV6fnsxz7FzpfYiXqKy2PvQa3
wJGbIJWhDP0m7zuvO1i6eWlyz7Xi6poGDCw4n6uptVo9k6gPLE+0UH5IOf6EdtJM
9V1QRUJtCiW7aQPViMo+JIENjp/F1h6NXciYspX0KE0ltYaarGVRAghWsiFzCBia
F015Xh6n/p5fXZTtbjkbqutv532KRDXUiCollkFGu3ujKh85wSSxH8r3Rsn5316I
RT98lZ4H50c9PFIRilTGrsmQR/4vxI3wTw17Om07d8cUOn4kaeMD1VT1OzY0qDKC
vQct5hH2nSR7NdVigiwQtQUwVf71YdMDvTxqxDFpkebMtzMGDWdP1zbE2Mo8Fst0
L9dJw8RS1x815p+78GiKn3ZWdLAAZ821M7o+EgVNCF8ZOJIT5F+iUsR+2LqavRjz
faMZAKbOwGdp1UncO7wY0ehtJoCNxukY2np5blK3snIw8YGeKs8Sx2r4aGdxd/dS
3I5LNk+cUcCSTJG/TxZdu1htj2wmNBCklPf7OlijMCPNRsPVSXfg1WnwL1cKC51C
neFVPcPV7/EzaK5ZD/xDI2ZE7QvyScZ0oQO2Utyg2fGe9uE3Q7qULo75q10ibwfF
RvNk/fZkEUN3VOV6c8U52jocjygDr1Ksjg55U0IF57vXrJVcZCRwFRJ3q/IPYqnK
Epdoi790a3Ad4SGg6XHrfCi00OAMQbJkcN/3l6n3kMCZN4HS4RCpohNCI6q2G43K
mosJhRRTlpw3H1eZ0R1kQD2ri92X6CLAWXLJCkrd6q6b8eigZjkUQ/t0wYgTTFKz
T3tXuLQhpy1z7WI1rnDL9MmezUWAHFuEg4rZQwcTLsffrp11Kw+ZbfR+loIy6VGf
7K1yAEP76Cpy2YfrpmtY5pzAlI1kk0XxS/f9rFO5jAiuFPOmKlKUcabA0tiZuWv3
p/p/252pnhLePuasKyp+sOrsHYKrFCDuvgI2uSNQ1s6ly8q/ydkWcTlBz4/WLTNg
kdSgYmOdeq4j7blA0gRj8iZCgR5m02zrBPZXZk2PejvllSpgJG7q3K6etrG3bzAL
MST/seDCTmUPb/mNJDdfvKUmuDRlIJEPe9Db8sPadsyl6RMIpvoC+QtKBDEY+yvU
zxmCihd5Kwy+eQ5xpfVMlKoI97+omt4TcNWB27jy5Qri7Jp/HYw07XgOL/m4jKAl
59sLKUntmZ7xoOUM7eVKLQjKDgewyaA9uys5BPVtJReNIH0LDGYxkchFNLojHUD0
q2XXQRviAWhUNXOZvOdZzfzyYVnXFCv6FpMdHM4z2XYcLwS/yc2ecFVcBVzETYZl
lcBDGSc6DUxJwva3uMNX/xFrn3HSNUfdwt1X2mZJDIQKyYDrmMKcWrXV27rsbByO
G32gXQLLQDSGPDjOMAXJBUK5zlAGDC/bkOyO98HYnPPAH+KcyVRMXgjByHsaZqv0
Gi6Fu4f7frmqK4N5s6tziPjV4u5ile1zeUBR0jRF/3SGA9Qqr9RPimSGJWZ6k2KF
TVSrVivOmSPn2+aiYOfxbteOYHxxyCYrMTJDOIuxf7P0AWUVxgKwhR2ZF72dVnCh
aRcJi68DYimBkg0iVjoapEn9xpulsZyuWUksmQWDRqWl+tHXQxtZwipP9sBPUQjr
hFMeLlVAeO5kzWnnkJxnud41VWwcoj5n9qO5Vs89Z1kx3V02TMQsebMHQ3e3auU7
C7chMKxOxox9fDgo86Yk01hrMtse/heDEDfW65s17TX5b3NX5OUwkJ0IWGSsm52o
i8oKF/Xw/dXpm7hYu6MPJo3K5UpqEhqc0UYQcbahi/9TJGREEYUNjqPL6ZuO8Ynk
tLCdYpeKXb6GAfyyseTkmYOWl6X881PpOrPig3BOsCaSdbnzyi0m5ZYLMMl6STuQ
gMo0mDOT/tiqGpEuDMFk4j0F+rBjCV0xjKBgbpy5d1iH6mAg+WZOkdyONgE23bCm
x/dtvi5kZGKxoIQ8lJtUObA57zSTiCt/35pR9jl8QSCTr+GSmg0X5KlEsF3299PE
6Udi6zcoi9TXOPeZ/OTy9rm9rw2qWypj9G9hN6jxl06Z+d4ZnjqVSVSW/Aa1H716
P89P5z4QfC5tkTqvqoVWb5AwkCslXcp4q7zqnsl4y3yOEHd2LstT4EnJwlqOW8G2
V4lr+NxtTOCDdcXyNLOZyQ5vlcX8KrojUHlEcEetzqXcSWG+XKQopYLWwIMRszmz
OOTXGBCOC0MNZSbEqTS9ba4GlhfhPNoNpHirie2zifklpt0+fYh+nzpzVvqKISMM
wGgY3Os6HtFs/IYNd9K3D+nRqX++GpUQ8cOPwseJ99jJQd8g7oth9QzZVLgILpzF
YwOLL9jqKYIoHJRasdfenSqa6SGhNDta2wtBCNNw3WL4cWG6WznzJU1xHQOYA5q4
31rc6mLKnAigxrE0/NJbI0bN/uZi+zqLFH8N0LTow//akbq9mugYrdBnLaJOF/YE
cNI99FrYuZEcWGKVWVbgSVoUTkuKVXKQfB7w268yowxsqIKmLVJXg8NITiMmfRRa
TpLA0s6xoAnlbEH55oTHypRAi4H1NMsMrOVcWpnE+Y8wOQwWDeAvYDbD3BgFtDcL
pPNY00DQiqWpkAD2GKrbnia/d1c3DNbi9SPwJ4lcvpEd6T3T0apACgmInyq1jza5
RcL8tibOkn7FWOXasaAYQ5up2q6gLcRnMo048h1doMRtnwwOJGoQlkgC+d/4/2Be
PAaAUTtygZ1oc8yYWwAf21VYN8aLJPcfaTcWJ2CTqMYeEDSWQy5zJ92lMGJ5oUBl
pTbKq4Pzgpe9jDPQC6NjoHs2mDrP+wIa1geNLdCbWsJQ8bWW6rMkKXIFiwIMrhUq
e9xwq3KO8b5BmR4LKbY36s22N1wqy4/G7hPSbNbkhp6HR9zHEiNinuFCoSIZsM9Z
Max+yRZ/qK3iAxLa4gTYY9qECZML9G3xmyMfwr5pfBwV8P0s2RTG9oJ3Ek7pGJdG
j8Z+HzZjFL1HivF79RCNsLyr512bhZVQdDZanhcq+Ngkm8ff6mgKSrVqZYjBhBXf
2NeaZbum6rWJ3Yj3Jk+PsfTppyXb8Ikhrt9cK0399KjyX85Xqrruk3s8LgstqQMF
nbVg9zpy/RRHXs6q2mLu9bpcEf/ptWUk5LXoSXrZ+8phAchc92BHMjH+1vYpJMSP
u2N+lavidVQZ9YUSy6mZm4Kbj51fVLDiYNPnARrnsr31Y1UaGdvndhOjfuqFW2fK
7gGEeO1o2gOrhDg2vDEr7K4e22ZNvx//7Jhv/XY6xx8RuCqfqW8631vDQqHCXjVl
ijAWxst3qaXQku/+2Yb5AgVb9/oCWZYPClVwna1Zv0PTIfC+0tQxgVGVUjGV3z3q
cm86GxLNF1b8Q6BBrh5xi7uE2ho+BehpTfXcQO/QxlYKjGgwghhnytaSaDy9z2Mt
GGsH4Sp2jztZ3ySQXwdT0riFnhXK6XR9RkvutzKLgE/0qYyT2G3BpdGcHBcaZZ6U
vKJFR2yb6FmUdyYi/kQeXHNKv6SYFIOdz2RCKcnyhgjnpZ6woOd/EwVyoPxUQUNf
+paV8//yzC4JhQtoIAx+5a/LteJZKWF9yDl5RyBbkMarI7GaqI0G/ewQWbMEXR6r
iFVyHrfsn3npJUv7aAXZUxnoZD9HioPuMWTi8ObbYA0lts2qKNnz3QNtCsD5X7pY
05qMrr/JW8kVXusSWliflTk3Pf2GcO504RKxAvJi0cfg49WcYI7XsTp5JP6R1f34
tuK7slYjZVxxT3PUIoE62a9Ol2HOwavhI436LlOpmAelgdRgZtdUspnGHsIC8xqt
N39+9D+w5bpD49Q0hwDXTttDshKdLXr/GuEg+RjiywmMA5ftfw2LGBOT6/fAtr2q
q1kFStZPrlB+Kq3q4RkpZKl1CdPdJy+g6PHP8BomqLeI0nsmxRqGt4fUVDbNStA/
abjbBVgwExUbVeoQe8TFMHGyb9gFOymGTkXD4WLaA4LkXfC0ey4R7pejspF2p2NI
vVmHXlsyr8autDI+JEQyalMMzp+Pi/wlmfbTXR5b932cFBSyec1wc7uBPJFeYvpy
CJtNVT0oXoFqvxV9xgg1hywi4MGx/8qVkr1oJzTWmBszTqG9a1st2LAhnR1Mh5mQ
d6FC6vosKjVfB2D1fFwaVsRjSP/zkvFs3Ogw5VruLRdbcdz/3RRSezfVLP1lVTZi
/tZum6aEVSnqt9Os0VJF6brP+3aCjH7yKAa5aPtTBa5ol/WQSLYieiGnF+VVBGpj
gBUIJdwBNXYftXX/zdVhKQIv280ifG0pTVCK7pPeLyZKdfoYs6UQSsGjtm26xc/7
AaMTOLr09OJj4EaBZ9n2oYPf8MBPj69LBkn6WFkSLHjJolZPinqEUm+s88b/9EfX
hcnOm06G8RDRMPpjMroBrYetY1Opg3kLT+z64CA1z490HxfagB6+fRYnqdXuJrRI
rVHmKRSR1CITypHiiyQzWkYkJq+fUoWwaJ4bZGF5bBlnzrL8ZZsvHeApnBolmAbV
UK/wRqmBQrOErI4ub3T83cp8C9xs8EGSjdvmLfVH8D7sTpV7PMcPBOlgJMwOhcQP
Hwrb3yR+MlLyL5l8ZKc7Zf/1T8a+qd7Y2DNS5egqjn+bfYGKrQP0bfyp8de7IAAe
n2f0NKzI+tUy60VjdvJ/jgCrljzy5eKwLzaKdwoZixkkeHLvf5kSYMNC58XoQfcl
3eOodtwFL1PWo4jqHtcaMrlFZ0QxqgFiiECVdH3o3h+S89Mli7/piUAdwYNUQuRQ
Okz/B6MvPeDy/QjIAYejImoJSOQJzOAjMU7fe3OZ+8SlJUce+vO947oCn6PV9Fl1
wFh75QzCIW27nutA6BSG+U4j9HEgJ5R8uUE5COMJcrDDAeQUp1qnwuzoA8Poh3RE
JRj2nachtf0uJ4yVtURiFBlMh2PkUe9SVgON63BkmZkXuFv9St5zQQmt5+0HIr5z
FMFZuZUUfHaMUKzyzEwxLe4CuC583dUL5slHqP1xFnnAIJW5j40m+Il+asFOBqj8
ZmRzNZxvnAFV6CNbjPV9KMCjLGBP4GZwvyBmdAq1TD54s0jqeFRmabd8gRBDAYqO
y79oVYDxPg35E1XyOx/ymd3jZ8iYT32hZP1h8oDKVgObe+TKOWqdrSi9mIYFvp7j
4r1RHOJURdNejMcSoD2CUajnSfp+RYpk6iqYe+8lUc3ki/R/rThU5LsSgfcq71Za
ySZB5FD4hYXLpAf+csYMZiF0o0ehML5cZQFLdXcDSU4WZF7xiFbfOZLobZYtH8w7
GNjr7SZLpR/XBk9gpR3CCE7czEYftHC++Vog3fjZ4CxmkDkVGTCOcv8HO3+W/xe2
Bpj81Ed0Af/M+VT1DvG6iAA3P4dwDKT5H8myqXXEb2SrOK1AjGUqoh/y0pqRPfpI
MhtL3F9MpBeWXJ0N6feHzPlu9aaYHz43Ug3kU0cbnx5rDj9R8JbcX4xpRkx7ibdu
90mMCKMI76i3MmwHHQguFaPyPJNJlh0aCxH5yn6BFA18DCjdkVhF+z2INAeQCGoK
BfDrVziwIL0fmm7whLWbxwZswM8/OOfwPZGUI5kTrYaWF0hs38ENpwRXKQNPeaCl
dob8IwWN9OEUQX3hTFG5jNcuQPDT35lFSwKZNRUeoyMweuVHbTwiWVWovEz5vv0J
xn83BJJKslaTrM/1EEPmGBN9LdKzaQG1WARx5sR+9KGNDK23qVlzfrLfAsqvCV/y
Mv4NC6a+UrxMH7mlMGO2Q5UNMgam4MmlBmSF/tREzVVoGJxAc5dw66NKK2PrvTF0
PzKrfq8UPPoJb3ib4jJiAUEf3l9qMpQpdYqTeduhnZ5t2Y6/dESPl15wj29SVWFN
42wz/H2Kyv1ns8vJ7MCDzyOH4rHtU7zUzo7DpBUZ1SPjez+h3DZVyqKW3WJe4SdD
CSOEXvQo9leB6sj6Z3gUIYieN01ShsDguaOeM8PrLJ3o5ta8BvH7W1k6T9MsWOKB
gsQrxaTvb6sePbTgIZtZoDoxq/+VK9GHtlRo+49IMshMjlqX8C0XT3sRkZgyg+21
188SPt+q48/iF+J6G4ATNFhIdKUSBcsD6nFQyHqRtzTc6LfMDtUd6a5shFBpq7Vc
v+VNtFaIzLCHNkKPH84aAujnVeZSa4nVt1t9uEIlcAG8PzG/HC6wQ6nhzhXA+E1h
rmrPXy8qu0PB0V31OWTKreV6cvNGkXphMjHlLry9ZyTeMJB7+1GnsXhsQ9GUw0SM
Mri2JmF51lvOJT06vYX8LVpjWsJB68ihlsRJ7AeztGn/ZYpLJpHPTFyGU2evszhD
WyB3afuB3QiZcMqDIc4IrSrAdiesGQG4ASXJtIX21i8m1jycw89jQl9ncnT7TZHp
z2xuwB7KljgD6Fzx9QjSd+LvHJU5gqEv/+u/keUG7wMge//t70zyuHW+T45IzQBq
GBD6H+0edYgrO1AUgMedIDbTEak1/BoLk19C4j3rVQ/9ROWuWvK0wCmVvOVrh9FR
8YqyD/030n/gf0bnO+9D0KR/PnznxagHM4KrUcUPlvrGSJ1XXFUoCUNF7eEIul5c
2bYw9luH30o+POyMYJsz3MCB7i6Ew4xCEPHeVwgPC0Tk2gxR9j2AQgZlcKeVw2c9
mPdOXfK29ZQcPHYA+yJ4n4q7OlRpX90BXqg3tLB88U+WommD/qaCo2I8/nE69dA7
rzyE8CsEGzBNqCVxEmGW4jxzW0G2puqJCj3P2N+NIzEso1m7hUq35MAzXp4EG8Ba
qmdAbiPSlv/wlEb+cvFmMtMyVwU8cLEFvess4Z+zZJ2He++A9cKIbqcSQtizUWgx
6oBFCBblRi42mi6Ywgqq+8ZCBrmoW+a1EsQryru0ZnO5omfHkicBme2IXH9skyBB
Nl0ue44BzCckcjU2B+jaY/djtkGjGTzj5Z6k/igu5xMsmm/TmZ4uzMkhux6dEs0u
5+/SpSPlo7iHYpItDpzLrilK08REqkc5oH/FKilwcJWK82Rri1sV4a7Hg2jwHxiP
ki7mQEg+4OGBE39uNI8Gxm49xpoXQzwg4ByWdbHaBmQybmMVWojq5vPpa/Awm5rx
YzSH8igpP036eauhWiJ6gsPZkXaehFOZDTUa736k9T83kviOe+BJ+jjGppKSbAAk
oPPPuDOdFFGgO7SNfaSQOukfX2ESj3nozL5URkDI0Ye+6WGhFyPgCfMcZdkAJWV5
hEhcYN394MfLK4eG158419nHCgjbAGbwQiSmL6YX2AseIcollQR6afelnt6dUjU+
4pQCtGsJTwI1vDt8fxlneZYUw34QTP6VSHdnhz4MR/MC36u7wv/VxoGOvh+W6WBQ
Dl7l4jVSJpGswbsXDkKcMTBrD5diI3SmuipkF2NdHwJMsUiI8VZtbFRbGKO1DlIl
YuJIQj7Dp3wG3vnTg8gzIchy0ARQHB/bruKyQ/2er5aUYPdYx6/1hH5bXSkBpiU+
CKbR9K9OOeiPPAPFiw0k5AzKaDWRP+vKnIp/o14u+51CLq4p29CdZJp7iXpiAHNX
Pv8+4K6fSf1U9OwxSN2NsHkQS35BskNDArPwBQJFJixa0s8tbeoJzB2FTUzXV4lR
X+dQeBw1VIyUvnkk77ozEF2cXDoIpbmCT+roawI5NVk81Q/K6SyHeoXILS5/munM
RNPJT+3sL66L/2mnkG9SlRZLIP5G+Wr9SiZNV+iuIcRfCK5z0ZJ96+XnluKfF2Hd
FdhJ/4NHxkAXNQtYsDr6bpLWgLPL1GhzgJ3YbNx+oGQ0jbflwMTl5r9naWuX03Gg
RZz1tKmmB2z/8DMu1xx2eYMfxxL8fhDECJ6wf5o1juK5uIn9H+H0pEXgncj2dIoI
etUYmhCzF1pTUW/sgT/xIALtbg2KRnjHrsERCQJ4iBjc7n5B+qtypbNgo6lS7avK
uvkBcfltiv7ssf1O5XqT21DLDAFxo5AjqoV8qxYG//7QphDTGq9UECqgLNz1RCdA
AyA4Wn2I1zNauYGKIS2GVvvm2KwQvVbcMOe6y/lzJbnC7U95Vm7+NsUQPopEupQ1
V2WPehRL6fz6UmSjULg3b949ikQCmSWb66TI9xj1Ngg2f40KfFp5+rROan9l+Ono
UEkLQ/croLXRRZz+3Avbh6PrQ3qlqg+GtWLwrq7A0Kfg/VWjehSyoqvHcr/O5/hk
c6b55IF1zqiJ4K7S+fnuljIu+i33A6gu3QcII/ujTQmplQPU5s6dHTruO7BhehE/
dulCROffoYkdw6Rl0MQzOXOuZ7Iu+XXmrPKGB4G4K4KFj+Qp3A9V31m2rlT4CJUT
VruqnS9e83nT0ZHYWQe3pgHnzkAv5T1iqWi3q6eJcbhJKdqNwMabphnW2r6UevkH
A2gaMtz/WnheaFdHr8kyMAw/kJ0qnRtdvR3ZPlhM8U2rMVthj8l9UM+qJ9U+SqLi
IKrV+ZP/PesYRqmW5sCSlDYW/vck+KXbGMiTwl27TnK8I8ik3SF7993r4zuNidYF
o03VXn2N1s3Z+0xEUJwv8+tYB0R6I7iM7IJ903AsTtqifDCREHv5N18VcrdmBdnN
01EZGzBu6bZQYZ6m7S9lBbvCJiQm0GBGp/SAEW8KP6j6IW9H6hYJIttfhyLJJprG
AZxR9QEeENFZz+OUodRhsy8ggAhYMHYw89y3n4+Bbva67oTt0xTrS3VtyVb5XzG/
xrxqqaWbE8Ae6wglFWrireMxQqNrlCQIbWWdSN9MauDs54Qj48YqClyjDH9+Qrcm
hk7Me8p11l6nggDcoFDefs5raz+IDDjsLAa1kRVNYxumn0XHZmc4fw0nvk1ipi/R
BLiEgGmY0n5aUOe0Dt2Wgl+s9CBjH+8v2BgjsajpinvXXikOHx+GtMIhnyl5597u
B+RS2JkaJtfBfzfXqddHuUQGf5ni8xuojM9fiKwXXd7fDvSBq1JhHzJT6cpZrEGk
ashrOELu6xaq6ONcL93TQZmfz9c3vFk/SyziCAZTHwqmTRn0dNAtDyikoewhi42+
4mlWIDxj5YbEF6+md+8BfW9/M4Wj6DVMC4OHzv+kXVwRM6YNqQU+LvNhOn/V8Nyg
zvvlZz9PgQuf5Pbvo2sGtZK0E+OWwxZpkcx0q0YZjVtMRIuqBG5v5E1op082RjWy
hGAcjXL591SX6cwg0IgfmZ1yKxP6tUfEgPeWwJUBD+aBYDy5cmx0ignGJhLbdcfZ
y4vwirCbWHO4+y8DE1hIIpV7Et8W2zRvzwLF1m369LwT/QQ8RiE8enG134CvzHH1
v3pAVXLwke8z6XETNsLJ2YqIc8SrY1Vi5TftAZJ+xeI6aKbFoUsWwJiRUvic5ncV
1o5sGvs960zPDKeprUlTm1XYKIhVdmeNqP2Sm2vOP+fjOYX0+c4G2bEZp944OqiN
9kgwD2pTqtIYrkZm7CXCRdjJ4XqpvPBmWyBVhDzMHnfFmsdFndBN0s5wsx20z+px
VKlxw+SYd/r6KrGqwpz921DKV8r+KZyddHRydHllSMZaAz3ZBXifa1LEAGRFFY54
aAwew7WwObCgQ6/PLdeXuN6IUp3qbqutM1bMGk2lVJ0qOJ/krRFq0QnYZ69sh4h1
kQ2fqwEfAy/dC6oZ5rZ0sxcr4Vcip4MUu2A9+QSG2u84NOPC4xe5N3t+QzVMuXK+
cZBM/x0ftcCPqAzm7N2tSS78sJjmLtLhhBdiwZ59Rllwz5Q6UgOrgTZ58hqNTnXM
8qM2P++Dhou8UZXLOQSaotZ+pwmdnwnQh8QScXcuYdh2MQgha1/dNLnSsbQp2VJC
J8nbDulIUvAyVKcZ0wLWy8CutiWsiX50bBgULwKR76es3753g1uH6r/VX9aZRSHq
L2TEkOe5lcLGhIvgAPeFlpbko0H3ZLmhCwE0ZN/GJTbacXC3w6X3hEnQkwxob6Lz
SOD4Icda2G1iE/BWX++GrGGDULfBR5xKa5kK3v1xgHmJ+nHxQyS+TLChvGhCp5sX
4qAkQ4f9YhFZaFN1ab9Y9FBr1PV1JTohqz+MzW1miJEAD7k62+03XT5HIHtw/tZr
eZw0DWJk2Hgb8oSyzS7IpELjCOyY0GI96BZKb4TbJUobX1L77Ehbsp0VRMwKdRcx
elQswpTKkK0+hPRNlIwFGtIc27chn9vHDCaJnyQ2jZqfI6YC93xGUT0pvm8k9zgD
8i94MEfBpGhevSh6GpV3O1AP+lEDy13bolInOyqUF0B/i9ctdEsOJI5pEAUtbqLA
VbjZZXONSqFnEp/dPg/e8xJBsMITVCJ3CfZAunrM4vV6ClKn5bybsrcDCg5FgmwK
14vrdEYkVylqzQPh96U4Ap5pRL/bUFLv6pr6wqCx+/Ia9svdeOIfhUDawUa8YQga
5Rc24XrZZbW+Eb4bBNY3WLrsQcrbNPRQh/ZrQ0VVqwPbDWz9eVXPFOLnbKx/WRJh
29bjmzx0t7JU48c2/RADpngJhgmYCo/b21psnsBVNdFYgocBz/XPy79pTw+L5qpw
dxJ4/5KWdv9QtI7fPSHxNAPGuha8swCYmkVnNePUsSvTp+6PuUZ9DKWlSSQ20Aik
ISxfmCQcXN8vCXJbLIv3trX6bAev05LJZk2Atgr22CGk+uZJl+Jyl4P0IoHF1QK/
duFPBFwbkve96V8ALxdvJQhWcn/d8JbHn1rGaegf9cu3s6DG0GAcT1xYnDZvR1Xr
vXILP2A0SvlDBuTqwFcYbpp/aE2/NHx9eu/vp3rxN58LmXK9je5WINER1FLXfDfP
EtELS86bYSRwfe3xqa24zQ0608Ixh6QYeJbiY/ohHwNWd24oPEA5D1mSghhsgd+s
vba8PG0VGGzd+k6BuNYjWwrVrLiPUub6gRyHauebg0m15i4e8evij6XCBeXAMfs3
d4Bt2+b6AP/K70MJCMyxyMunTmBxZxMmkwk/dMDoR7F/IhuMv8/RfSG+TPz3UG+X
oXpOGTsD4jPUBnd7Y7Kkut+9PM8cJYrWBWuGOp+I7JL3wP1GYpKX2QXqPnKxbGSc
fnAh3A3HoRCsNeBApsEjTE3Nx5sbnxZ65xPg30tqXq16+qyKIiBFBaPlCbHtcDOw
avPtUHaVikShaAP0Rzay5s9HVRPl/VdkXDASQXwi6SW5CngVt1cxld2Z3NEQT6ym
2IVcQagCS4jfRIZXsPvfTCLIZ+WbFaVOi33quMjx3NKwGIiGMnBc4Lth0BSlsCxf
yLK6LhskxQMl1agp+khQivM2D5qJaGIfpvuBVyJ6YFKWi+jyq/4Z1DzQx7DnKuap
c3taBfkmtMEB7QoWWjyZFoxZLTGGLYPPpbA3FRzc9s4NHfWgUUsMPoG1t5Xpjq72
tw0c6MkHVSLrK4QUDKmT5xJUiT4q39DlW7KGyIQ04DjMX4vgl1mUCQrv+LlvHpJf
uZl6xCMh3n2hbZEvLfRthcpgVqGXSq/xeN4UehOCPGVlME0aPj1+DqhG6kGtBwEz
dx5OX9u+9zlXOGUx+Fa4plccA2BXFg8vuvqcn7+Tikn0g1560iTlEPJ1KtS1hWz8
Cdt62t0Ib+gwxiSqkkdzZ+ciU7gEwsIsRR0qpzkI297pgcDKMQt3Q4BH4/vlqP1A
xA2IhGBqPBu+t1fSBUUMqU2c99doC+SVLQ/dsyfI5UookxpdKZ0ZEJGvkp001Bca
zGrczR8YzYnRu39NcGWYsIK+uOZaQEvBlxCMtNLKxk7T7WRZGY/HVH0c2wNbrs4l
zo5hKi0ZRG6V7pj1X2/enoNH9k01ETqcUQKJxz8XwD0bu/4ymB9D7zDPoBtmQgOO
o43V1QfuggFlvRQKA2ZHE/yQIgZEDEF/70uK8MXBzdIjJeMrKZ14FDs4AunmXOvp
D7nJ1x7EKAw67KbDGCYFb3DClgXdC6LHY0Dq3EJ87ycAA6oebh1hverewPImn8p/
YSw8dcGJ7PDJaQxhVC8aG8zr0KWsBG7Ty2ymbKFKSDe84Yl8rZwQwE6GvonvjgVJ
Iz2I7pebgW1juJhrAFepOf8NsISgEAwUmkhPHe2Nb1uE50cBMqy9b5XH/BtEU2Vn
xPbN4VR3WMx/HGN2zPxiH0W86n6R+hQVTRIo6zNFfwIAtKhFolinkKZHv3NLbjsA
kDl1NDDzBt6ndREcHIew0/3mX9kT6LEPH1eCQa5XMd89UnZYxPR8Q7xs53BoeedZ
ZfEGFha39NrTQLtPRX/XDG7f2BH41j1ITQrMBWesKQEGPPNFt+JC7SvdrFvaGs3F
FxDkJp3sI7TXbpT/Uy+bRRHT7IZBxsl2tUIiD+3fi7MQIWvcRxB1yHJ7vnsfyWOH
FktEhCLvlm3m9i07bRVw6Fv/+4jjtBDEHCqRn/DPJZEWdxBncJblS+FEcaQ0eRpV
oLRRlvAWGaIMKKJ02I9JbR8FvkqWaKpZoMsv0LiZgLhkQSNrXbqZJh53EnPfRkQ1
iir5wDDdtLyQESoZLC7d0ZloW98+iUy0GdMNxHlF31ya7kK/u18jRV79/maPhNIy
kY3JiS1TeOPyMvMV8w5gkFggQqaaYgYAYdtyXs9brm1FTkek5xMVAqYfX1n37hAi
PdphDh1oryMszx0HQfZYtyns5VvGPi/lqeBKpf2/kpmB1TrkveUlrmf5DBEoj0ES
atMhDaoy6G8ZTsri96pXtxg4PJhx/xs3xHEw82hCN6TcTCiY+KnlXFRORF/QdYNq
upLsMlkd/7xCOSsFeXostB84v5aePbUMK/OTGc7Xk8XMjqTg+6lljSPV/wMUpl5i
nMOkXwQmzy09JBdvo2H1sU3eExAOQELlS6Vrz2BK5HouUFMWJYAHuk2Puhyqzz1A
KVlyFA/kJ0KZODM8KFtfkEGcOpS1L2Ac5CFQ09ES787ZH6Mvu+lXXpHBfGHjBdYk
taa5UQtAJFAsGcaWwyVKWdBPlukjy5LohVUBANfWMEuzSCHQJRRUK2DaQ2DOSl52
J0WW1jaTYMBgLMXwG0CDwrR3VWByyfb6CTiMMxDr6wCJV7ejmk4hMKf+AIC4wbI2
rAQFLdVB00sefUa7TXmNjKhoVb5iZSDN7zaOZPjzSzAulIz+JQLN0JytOSwk2eiy
61Z8dtZqj3vS8I+N+G8Fdm1k+Qf6MrDp6VzdxtjbasrJFHiVlGQp8sVsPEiWtlwZ
bzyZVgNvZTcxk8/qHjw3UoH8BvAqBWbd/uOIhKBVvq7HXv6jCLZgKu1cjWgKKXJk
G6eBdsfDnpzVcv5ypngGBfpbFmBLaaPo3X5NRA9msf5oufCugtUNFofuKEF1fe9s
GG9Xvs8Rje+1RLHFehTu5IC+bXK8aqfR46JWyOg+DX4fC2XqHFZfWT6ifVWMy2Uw
9wbsnl2QZx57J9UHlIMcn9MrO1EtCceLTJN88VlHqEMZurb9aAfLDGXBkTkhzxWZ
xLizMZyZaVo5XF/TsRvGn/OpU+kClytU3yUXLu1aMPMR96PSRcS4/l8JBIAbjc59
aF01ZagEsQMWzjJRyF+USbspSxMJTdv6jETGQSqaaIOMfBdx81cwvvGhA/lSgbAn
ISBtrjEs+TpQdk+75lfIbbmhOSweKV3/GKavVA6W/HU7mDxeedxDQ5JSfHnwrR6h
k4RzmQE5wLnZ3lYn73FjvDkS9BvbpZdhFe7wobpqWbejGdmH6P6rhEVSBNSaOcCR
snady5JirXWIVSLg5zIboEiyzYWr/Wc9xLjM8pefl97lHNC3QGxlzLl0FcH474z/
Q24IHv5+lUr6RFS89n4x/RtP1gZlVp1FIk+qWvntpMNQcv0w0PsjfxsCGDAEgfvb
mTM3koFZkPyx6TbrgMSuIhpRvJnA1lAd/4agMGHBBuIi8qTIqLOTRy/hBom9+ls7
0y/Dy9Opb3h++x7VM1XsuLGrHBZnk4cloYmDO2TqjGlhm3RxNGM6V3IpJQcGzAeu
ekx/YVV2lm1Xrtt+4xriv0mZRILkWAmehrXG0PxSj000Ggt6Tpf25rbWR/GgENv2
/UjdsmZCBenuDe+wXws8CD2u/yXMCkvEDtXTJ+OZ+g2hcBQxbhDOW12ORYOO0lsL
xo/dkXuDaqzU5sgCxbG9nbqdLHGStxlYawQCSgmUqxYNqKS+zifgsdt2qoZycvI8
vcFfvW0g8Q0u2UCUvI44c/mD2Zm1sNlOOcM1YQGyvWIWRwbFFSgD8irgvfCcggEt
FmQPk0zA2n8l6U37IKcZP2YbfMhrN1mEqVz+FEeGF/De+x5yznuNQm7R1z3+XFn9
XBvMAYcQB7X0K5c12os6rvwTosEjmIESFkSXs91fgTSgcRF0vqNXLJnRZtHT5aSy
6dEQ6lrfuwTugLJBGKikGgnK1p3cYSUSZGI+2mvrIKAf/KtYs/Ka8HE8uy7zFev8
bwSXpXX2B0jTq51kZqe5bi9RrTMHzKG2pgs4uoPI0g0zMes5qIPfz3zh9XeRqKr0
fOR0gBdIk4kY1Ie8I/56dufCbxKajIBEiig+apszKkAszs0evH+Iyru6mnFR0Q4K
gKYvz3QbfBEgk3+mP3uVzESxGFx3R/+T5JOIY5PL0FG6iPG7o4O5QbvOuVQ0MBhl
yuKAEX4LoezFIe23sMh03omXrdSLq1Oq3pxkNfAF2fqgJIprpmN/uYsnwE1VS8To
HYjZPXcAh82LggrhGFAntiBJ2K5udsY7yQu7MX6zabdmLIm72pzhsZQkFRR4fxyC
PdHnt2WlwFlWjMk4R+QA7J7MIBDPocHfm+SGerYw694NVhF8GneaCCZX+pXWy5UH
jql6HwU9ueYjbu4ZxC1IUWnjaBkD5Lvdk3Lto9qOYTGTgIlY9TSMFwF79HO2YDZ/
9FXiyiFT3FS/L1Qk/pJ5u6dN/OIcykETjFwvRy00uF/SLH0zvhaF20jizEa/NtUb
KnhWqgXrb7qvlAsaQ4oRbr5rHRyM5ukXb9h3xa2xdIyEnpaTHeoW1A+3jjHOgby4
DJynOJZEyRu9LF+YxU45U28w+gY+1IqETiwIWjDeWgUYTTp11I2gvOrGSB4IgkG2
x6194aaQQC5YPO/63vKnH6uy8li7rx/5EdWxZjDWYadAQ1gOxaVez5pq3OAvxscj
xJ2r4wie/Hdg1mnWjJcYyXci7UC8edJrHu/T6vuSRzBxkZmJmgE42Yty0rGOw8lH
KgISuXnXZbTPCe2zF1bZjbAoyQct9XzVHowU0WRVB6Yr+m9VRR6fXdumv+lsCXKA
LoSR3FI/0XZ9tsQ6ckuzPYlIDxd7yko9dB1t7lX6Wr7KnvtTxozRMM15G+Qpyufw
OrI9ewHxdzfF/yB4mgx67XUAtWPjxfrDfOOQGQCIjfnaCjv0gPr9yK7S5LXFm1XY
wUJ9JZ+HXDaH9djtgNdgmaeNzllLrF17D9IPHG3tnokov+o+uB7mAj5+532Vz6Yy
YKXIBRhgWi5+M2Jenbuk+MAhg4AMXXoxG3DA7dIRetZ42u/V8I7NXWUgUbmyMa41
OooZAyeTquMb9KoLEV5ljKmJeqZ7cwrN9CnF8SOpFSeG+jmqM1H1agaBFPCI1aud
iFsMBn8KZoAPr0ZGFvXrHNxkERLpXUVw//TRyb4ETUsEe03IA0Q0y2D6ObU57glX
wo0getYLXxbsjcaGa3P0ihmPM/3/2bLgV5n4XvVqJfjctW2I4DrYFH63iIcTDlTM
5a1yXd+K56N4tqzdzk/xeg/zFkXSGXb4+MbFiI4kb0DqZz4kLRpiohockqXhbMO1
c3ofofgkaqHuIhU033SniQuhMwnMaKLek3g6hIhj4+WsBIsL+uP9iyejTlsX8vHz
vvyOir0etOvbxuW1j88vXVCddldo00Z+7V5JZBt9sEDrpXaBMrU6iDq/8C65UDMY
JhUBTIURc5gd7YhRxxZyboY6chTmnfGML10gjrBUbLuk1lkL/xbbwXEFLU1u/QSm
KyDZnaolb62g4b8SJsjVR5w/hVjp+sdobvstzSeKEJzDnA53n46n+bpdB66T5Vjf
ZUqIXvJWkHBZX8xYvjTZflg6GKkPbckJ8CZRj7LSg3SREC5c1AvoRonxMteVOmIw
BrIcghbp/rxLHeZksxuhw32OgwOdY/V9MCddRCijxXNAE8au2A/DNk/4BqwQ1aEr
8N2BEC+coYg7B07wdapxW2ysXUsXeltODasQS8p+qAQEXCAV/+TiipWmgSRaZmNb
LTopYn/hcbGwlTPxP1636sk1J1fZaFT8a6S2Pf8iquHRxORMAkX/P3yVvxSCWI2I
50Zq8W0yH9vfZWN6Uq33oCmqhXcHtNnkBrCkKyX9LlMtaRlcxQjvFvv58ixZ/NKU
SQzRo3JMGbv6tdBkxjBbnvyKRiao3HOF+uiZoKAD2ey4t4Y71ZO6nDW19ugM7YHj
tqI+ShDC1liow1LQCZwwoJlH/wXkvfW5zqpvKdPkFATuWkltifqEZ9sAGagNjmap
aYTyJDqLHMqpuC4sLiSnilpWJK5hxS/gcCiw6OwDwPJOGNQC+A0GPwkDsHBXjm2z
ViKHECttD8My1wyCG9Yt6qTYGLqrZM8QD2HzbTUujK9fZVQGdUD0TVf0e7ZPKMyR
+AlMBaqP4nuhSbg5q7BrSGE7nc7YlHlQppd235jdjqxIblSD1Fh5Wbr/2D9YoIhm
yaH80lfGSlUFAJSbrwoE7/yww8A6a/YbMORWWRTX5MHvCL5P942QFaxCUnYbReTV
9NSQq25xLCyShTKIAga0CK1NC8bwNxqivBov/uzk7VW59lc8cs8k0hHOL8J4hgEG
Ri5bFrY7QrnHeC9ZWH23/IrPIRkfakw18VMBAY8agd2QzcJtq3dMri+QdQ6wpkD/
PPHG0kICmKUsFe2UVslBVNkpOmiSBp4/+eyIWAfHSLH5Wpmq/077KFAuuv/yQ0oV
5SHTAJCgJQo7cdeGPKuAH9xcNQcSp2BzITqYWMGC6dRn8/YJnHBHNnzwFy4ABtO6
euKn4js39WQMUqqDq7fSsfDMN/MAvvwwAp6UI4dxNXdl1rD56pOneFrraeLMmWhn
pOWOmOUJcJ1QI5WBVmF+t4pJXataJVkURNaxD4SN90JTuwMX8bB0QttZG7vdXjZa
iaPfUs7ZIeYNajBn1uu1MmAtWbLFeQQ7qPbIX7fUp+YQ+rNef7E1qVhNOEdnO3SB
9OvnRGIqPn2aJ2Qo53sA1/3Nv7///gwg5J1JQ0PDO85FNZP0rw9gMA6g3LTJJZtI
Cw4Q6nIcAKwnsc7a/7+xfIgVXeu83F/oBnML3qsjtXQoOzD1k0uail8jH3AKDR3u
2sh26VxGYrkuV577D4ofkTJAUpPNnp0irOKRwWFEqMB2OVpQzHU9U9YEgv7UCxGE
IG1lpWKN2ImmWOHdOwVTR6luXFEu4+mK+7seXnYNOMACi2N2+XBSHm52vkuDJvoH
Dy/v8s7Sf+RChaIriJv4n9AcxkqcOxv1zVala/LYC0nQAhHkJcz2vS2pXYHA9+Ft
CW0jlhpIbELmjrEHwIs6n+ju547wPpfHTRw/wsv9Fl3PDK/btsRvAeWijHuVDT/6
PqJfJhJaEqiY5s56kcFf9XYFoXfxjQykvdEe8F80UFfZHltIMM9olhS2F4mCC0in
9FYz3RxgVmV97XOLOriph/tyq5swSeLO5kgDGYXMC435QCyaLtutsxe/BKHKVFnt
IurNCygoe7r5qfre/2K7XW17vyLhZnvPseqamOwyDK5D8sI+AZh7yqCjiq4w1XGj
3EA/gkIbqm6wHYq+hap54Vcbi8Mzdtttr8vNNtYXN1f/UmzK1qnr9p61wgi65dh7
JKZvMssc0YuhAgilVTJh+ic+BWnk2//pcTXHaWCM9vT8bc5j0NvqFkrfGWpNkfE7
0qg/PwoL/+UgHtczridBjF2GM+EWR1lM0i0QlBjeggfEJD9s34hSJg4R7yzrtRzs
x+9wU3/F+OtocLX0NOZqYyqMucN6AXeU0aq68tilCAb3Zf4EdBC5z00yKhKrNacp
4uCb9e2kNJv4dTnDb0N7801BUga6kKWTnuXZ78fDw8O/LxRq3ZVBoZBY5PYHfNal
BYD79QW/M2WifRsDZJGx4C35cIL106vgGk1W4UMCsO1lLMpk2XUh1ppKK3HxRPcZ
5a3u/nYYEw4X6N6OPD+xLhOiV6TTZEH9eSDWEFjwyMzCX1nAGOFcdDQeeJ12sUz7
f7KxZ/plOkPnR7WlkZukWix4yWKoG0MRjKCxkITEr2yX2hjS0C+XkU73oftcmrfY
DVJk5oLP30eoMifvdw1Gi5wo0xYiqnGc2MllhrDZtjkwUkaqcmN1I1YKoEaP3dGW
CEH12fAfntDj0XIPlVrgShRTSUNp080zSjfUWSz7rjQxYJAW1SoPepVQNYyhsZ5z
vTzRpXl2JKNkHOZX08Z5PI1Xz/daH/fKk173NuFCJiFZswd4adlexv4m3ar0sQMW
yW3CSunSWdYHdZNs9DqnLOxxZIBZKnpOWbo17TVc7Kbrvs4kBohNgBWBXYZYO/C6
6X8hKXmEph/MH1tK043N/cOujlLXmUwk9mDbQrNv6A184sZSzSql2N/383yyHmF3
/I4HnMeGpic3HnY9myYVzDZiboljyggsRwlDCL84dsp7sEEDHtI1Oo7KxKuhBR6c
wdbvUuV2S9lglLUuzjMrq9jKyBvsdYIcaH/LmeLBJp2SWce8Exq4wksPXCh/YxkG
dDkGqhTr5x0grzC0iB2Eievoh1EUXli+IQsRs11obmv/SxLMh14edrbsL3AbqfAY
MkRwYC2X9PCN9asR+kTRNB3tlEIzMCT+dhAaZAFWk3NHq+bq8eL41ZhDfi1qP5Ej
8pxw+hOrw9yX2QzFFRjuQo7H57JyPFkCryNb+pjgXIfDnX1Q58uoSJNYueLS8nu4
rZ/0ojqaGXDBx9hJ1D+4BykA2jsFJYs2Aed/JzkrokWNQn6gFB/rScEPPrm5we9m
RkDK3TGm0d1rfpc3xed7Pzue9i/Xoy9bHNbHekh1Dn+gbqzEudOQ0PLXwuRrZyXP
Joxo0KQ5DqY1cnjm4DmolC/76SH+prn0v4so6TkDp56EKAXItR9Q0BraWgI8usjT
GkGxB565bhILdWJ4afvZyDXI5DePmKd3SROgnu63cCxTBnA/JTTM0WMIH8pFKmAH
7dNhE3l5U1IyTPQMnW04Rll8pGw3bb70jq+5dnAqMsdU2Er1D+fwGqNsR+1+r0S3
1sxzYng1GDOnj6bspFEr+r0CUS7/LN/dy86hDsbNgEvFFWY6kSjhOJB+5Hph3uz5
quEI64/oGPc3vZrx8tNV4MW6mCI4M1uwN1bFWa4YnNP8OVtfXM1Va+EWMl6P3/mn
LSg4ACHu7oS8dyvtYsIpGIHGus9hPdH/2xKkDBZLUKvotrSNqLy9vbCV0YD1v7JY
xvLjMkv3WxuahIwwNhYtFUiiCqLwTdW/+NsjYTwjnOLPhCLmFB27RGdbmv2bZAIi
2o5kHNCughkesbktXBGVUSPKTgakFp/JSJ707hpweeQ8m+CT3oWyXBQu+4g/pfLM
byD6ZiyfG9feciaYWMFoZtA9SNF0qhQRGT7uu8QXqOq8PRwKBB4VTxY6YoMUeNwu
hrGUeZwaHr6Fkb3EbtRgFjWmSxh8rZjD59e8iWBq/7tkYx0BdcxzKlD3QPH9vLC0
pBVex1JJVHPE0pUwo+USxx45Gpj7A0Ru9qwX+uXkm6PbrDpZ9rc4+V2P0xNiNbb7
aa7H4CzCGK7obo8gAvS/VUVmxwogMS3gekWX3NfhccwAxG4vdvoSq+KMHSd7XyLl
ta/dj0xLtHIEzpGKqTdxLB7dLdIrqFHX1OJnxq9VOf4/ag52FRK73xMcvfOeXakR
/G/7RXOGlc28K/+lGRZ2epWtlBGrZYrKcyTefh0007FWUSr0RsQtIQokjXE44++K
FPjaGJsY6uXsDW1b9uEvXxa6NGnkFmT/4Iw/0Iy2AzlNxMfPYQQrdLEJ21DtvivV
gPsaGHTEdWyNVpflGx1gC5Q0I9/dDqDg1ofiLnjAfde+BLdp6s2kc3vVHfatarhT
gz+fW8MWZh5/gWEGglga14x84OM1bxe+0ltCAGmUM4dJfVj4mTr1pooJujmYNVDm
p0mitvadS1DMN8r7qvx8HFwMeU47jTMZQCxG64E/l/gkTejaKG4hWeX+uFWMp48u
hNLyZ9uCKIb4+12FsE7uExHs1XIdriAwChtstEJY53HDerBSOZzoecYrjFwlVC8S
Ua9qjMBh/h/a40Pw49n/2pYzSce60U7OuNkDeBxnFvPj3JPRG944yzUpsGPFx6Md
tAodDOJgx7k7bposXFJybeU0JOA9ETxKH32d5WjBZkPmStxpglpLdU3cKPwTOvp8
CZHbqkGWrouBm6coSnU3zgMt6yVoc+wrYQFBHjuGKCqWIeFFcmqfMNJG1hRDtryY
wLUei7uBHdyXBJjG36EbBiehGACVPOJy81z8oW/tRgqNQ2Hb3ymjNOr9ZkTVkxCX
i0zznBVpKBmFlYBuo9VhPePeuC2+msFDaSgKeocjSWMCeszexp14xrwMdIwK/nia
okQFLl/cqszxznAz9DXnHGWcIfHc3ZVWQoK66eXS7bjzUbLbeEEjapCiC6Lt9NWH
W4s3G8bOi8hmRi5poGfsE4DfTFeuCR4yXNl3hm2jwvFXasYZVhcVzlp0yDX791IV
pPBdCG7OvuKTqpA5ZGAIxOQPGdAWCbHmriY9g6n6Y9BcpxoACOUz8jzLQ2uRwOYb
LS3WUyjfVhfcfc/t2+MQ8g5zm1hhlkFopAKpTueWdRib3qga+vNCV0AOe2r2CgiT
yB6pu90JOIWL3RXR6o60iOhjZwh0wpJa/y9wZgBFodm6Af4puImRMB6TLaPxFt2c
DR6w4akP71cvmN7d8JsfUq+07mHSzmPPvficEx5W8kKhovG5wx8paah4M9jgVnkM
LZxSxi0QDwlm1AjjgJmD86SfKUEmXTRBvSXBu9a1aQ8xBOCbXUHmCDM8OnF/Q7Gv
3QTkftYaOyR9W6K6JDIUT8Wky0Fzi6myw1QW9LxweD/scq6M+PppmfwtflUvmxDB
7cYX+KnF8lfCzNKa+kGQoV2eFbOQu++MNS1FXJW1LRc2FS25RL4ASwe6lYeoCO2C
n+uNwLVyuKLznDikEvr56/13kqGviLIs1V2rwuOJpBv5mq9lKF3/ifaAHZoKLor0
/UAZkuuoJjHAQ42rHVw6WCOp5obteanvSX+jhVY03km+5X8glaZx80kfXksfqlFX
XNarLqIICGmQ9ed2qjZ46v8zMoVv+b+GpvLv16+lqgEJ7bd7AEIl7vF5NqZlNaGz
qeieeqs5ZfW9aj2xYGxP2PDZ4s2P7FlCZtRg9/IAR/54u5M9UGczYtH6z7IP3Hf2
7jrxi06V/C8iLEzshdbI5dxymkPHgDYKACoxly8sp88Ojw1RZgizZgFJ3PTD6NxR
75rnoDnkhSTD/mDu3aZ3jwa5stYlER7CyOWzAsDAue6fJ2AzKMTGrE4ypxCPTKCJ
nLlsIo9V9eo8oubJOrSCbPAfcN2vuc8b++vFuhBUBsRJFQC4r5P7jy6wzZSW/srd
H+DtbzfGFgnPU6hCuJpzxguDv5WCSnNGO3uulL4HM/Hzx2G7OJgOjH4kIx4kBGBq
NdMT1N7RtdEgD4kkkRnIka37IRFEig1waxNGCQcN8KjYYN1kHu8ZgwRylVF2EorZ
2hj5ZWjMLIwHzk/TRpSS9kcx70A+kXWuwfKi+9Pg/znMFzjTSZXBlWDXe/qN61Vl
frDRWodOUVzAR5emTmxKtMV7UqKeqGQFP4XtLvPkRvbE2ahYji8iRxlv1RahgmUb
L+lGvMt8EgBalfc1bd99enMc5XkPtot1SXKyzM6th8HlljaX3wACNUNqfps/CNCG
7pB8piQjvwt2/kD6KizQ0l5bT80RtfeRJ4+NlZvWjOJG6rgjOAGsUAYZf76153Qc
Vtsm0lroJ2G2Fzjshp73oeygNFpVpXTy5GBOALWMGOdqiHm0hif7Hn5U/A9rLJda
x+IcuDTlsmZvcs7rvOjwGeD/mLkk2p9DQNu/0VK3iysRpphXgN1iKlWRkcQ0tFRo
6LUEwKrWvMrhV4wYBPk03eEXTSyEOf1vjzTyFySItE4LONDcOzRV51muNXQfMMW1
u6ORYSp9YhYm1qyjUyoavg5hjHNzHLd2ORRnQyVzUuhou4OUMXZQm69uRkKvmsf7
Wm7G9Dc6LxQrMIkjPZhtSXL+TUrjCBogUpBCd8KJPsEpnnojxn4ieZunoWo33e3e
JAuXMk0c/5HuPyfYlZOx/qbHAf0geby1bdIZDXeq75L2AtOjJagOYsdoSOqcua5D
mYsdSDx3d4tBNb9eoO8ny3tGin388JLGvTX5o/ei9Cfw5Ru6ly/BxzIFmCEqhbhm
NUjSVjaU/wK0AA4VU/aqZ67o94wdARERCZLNv74spozx7mDfe8GRpiCTuRkjwEZN
zfAfCqgp8C5JVqp4AR/D3kzJfAm3hSbVieG65Xu8TmTRagkkH/qopHSUihh3BGW5
h6HmUVkZuwWlqv71RZBiyyU7yZ9ZK4R+C0SERZAJpNfPWvB6iydIZv3nSTSY2CMf
RhKmJ3C8JlRBeKmcChxVS1BWhglD1mDS1txskqEGmUwg0OVLjE34PWJBsnE43pER
pgj10DHrBlhuwp+V66G8JVIJnL8CoIkbq1iAxBtz2njmexLXuHKNNwjrAOKcFel8
J2T2NS8tfWMKcu6mV8IqN884nZxWUh8/irlVjO5s31668FaekiFxcsOLUl1c5ltN
rkr/4p0cvM3qXDJvisLo7kc3gXgeiF900nhp9/EqYN3qO4l3ODZq1UAOeeiVPxOm
cLZSMmHbFttMKXmQA60fIyXzv7FkBu+NIFobf6HPGORIok2pvZcD1lRy3aBVUoM+
xeLaQZMC3J3H9R8FT4y4z6ymoOvAUCr3TeV/ul9T9mKv69fZnaS8Sw+vkr4oejMe
MkXiN8Uk6afJrAxFmB7BwQ6WN4lmgoFiP2PsXSyvfrWPmbiYOYErMvUEdBfA0+y8
+F3rGnZ2IVg6XPkZqRODjDz66JZCNy54OYGqau+LrWEYVIz21BRWABrYYn504VK0
ctOKASw/eHLeg6IwMwtZMqpnsQT2v0RhFQJIhT00VLbONO+dUQIo+40jpjInBI3f
Rgb+o9wlxkVfis5OBO9hbZ0y+KU7vpfdVuYhJet5+oX4Kq7K7p3Fe5RtkZDXZJop
TQdSFhAls3o8mYYp2wxEn2wg+/sA43GDx6SzUMAexQt5aVjaPZ9rmzHUix2TVDAF
nBa84PYe+Ydw0cPDovBMx9jPKin0qvZNubbwLOTNRX9M4ZY2EYezpwjOIwBBn93I
Z1VRRxRMTOz2MSo9tPRQm5JOMu33ts6NjQ+J0U6LOWsthPthGsAjAmK7kTgwuFx/
oE3P2SJyAMOepllUaLN9eeaXHrWfWlyei6ssig0cdN+TzuwFXu7mfaWsVRkqh97X
MJ7EjkuHtLRO6dCcxDblYdoZ2Vwuc/1n/mEIw4PNKZI7KtMV4HB1qA07YzRMuLXJ
9GfyPew9EJgZyrHiZAvqCZq5MAETAKk6cdYyvf8pc/XOU7buTov1+M1y9DWcOaQF
9j2kzi017D1vPVJ677s3BUNb3QPDbkP4fD3kvAXc2Tqsf7id9amG+EAw+5VkUAD8
7SM0DYrZkx3NZe9ys7gsOa4DTnOEfv8E5egOyAJch0absa19PbxJbX5o+4lewJHG
KsRi9w0QtF4JPgxcRlpFo2avOkw9867SQAbtR5+0H6s5IU1MySif254E+LQfuCZ5
CEi9iTMwYPn6ACauFCU8JxSQYxzTJDzSeQjN3IjR7PHnwmuzToc6a/ov3uEURFs3
UbRQNmNiEJs1xnbmua+P5x711xGV2qx4YIWSGi/AhGqV4+d9tYQg6yjtaHON8yDx
s2VXqFHr5ZeynTflDw8woGJyHRzYxukTNC5zVfgxljVxjB84Z2aXZZp35O4Y7vri
QR2uEkcUii1wlTevAdt1hw0BwQEkHbFM+fANTim0qV0DAk+lh9NHuIX7nqxq7fia
N5s4I/rAtcGAgw2LEyT5OvfTCsY6EQ7A7SfCNciuOEoCYVyGiw4veHvHf57A3BUw
i8gekf4Xu7uHcZPdQ1hs6ijYCBX/NSh2/6f/Tk7Kwn+XP0QLLPE2ldcXBHTqG31T
5+udZEGctd/JI+EapZ/WaRlwQVFGui1IacBf5eIhzN3jXkpyoRllKCC7lscDaYT4
AD7ishXRHUf5zEY72T2OKdEKB/NsMH0XENsdvn8laNWjgAvg2dczQasIeT6RAF54
10BWhvFDk0aSxhQGJSWiPBjKabgXAshgU5A889DCusU1iS4EDyZkaYuoUseU++a1
uMBrYyVF1n6kds7aqxn0TGvl49Z0Y2cIYn6/cBX7zJgtL8v9mwvub1pjAP35+j5L
eL8WgNf1coqf4+CDt+j83c1ZNy5E0qwT8DYWJ2eyq6rihMolEsPfQBkEsH/qREh0
cRuqMOUOQjKRpKSxEbLxfcJjd42I/k/yf6GllcBkPHtxmFm/FTwj3LFklDkBtecb
fXoBihn8NHGFPmnAq1zyFZOAjwH6uIGpXnc6HNcl/72CA6NQx8X+fihEXIGRcfw7
Pv9sisGoKPRscf720xjfyjmSXYSUixwD5CLnNZCb/xFx5XCNAkl/t1+qphcOVPKp
zBiPar918OUM1HRjL0rgS0knc7xUu90f2fxyn0ou2VtmtZvBOA8tV5WFFo8rVw36
7JtjT9HqeRNKMewJBlAvGdy19qtrGBySACs+QikaiqqcuNqQeeUpUn+UaMjuJJUr
LMB1VKncO5FmI7lrlDEgyrGilGwuJq8jXcXYqqJmH5QDZYEoGsaY2+T1omBF0yc3
VPi5aeQdAVxPlLiNDeklME4vEVZJJU2d0ZpxnCkawDIrxOWec7QPbZ53mN4w3VtN
tg9EbrxfW0n7cfQcVhzRFzpeCtvXkwzG6MwRQYyu76xSibIbOQWhUfBSIDAokheG
cEwbVpI7AdC4vmu4lqCXoqAMdH98Adg9Z/+zs9tJ5W7lnHxGN7A2kyS6nbK7akJO
/b+QQzZmmXsw3D1S4o0YH5KzdTqMyqyctOkYIWKCLJLzPFmVla5T5AinViBhRjFm
a43YRPHmP+EvflalA3oIEsnXtsc9gwpBizShv/QkEspy21ZvftgqQtowkR/hk5Wv
Iab40wgmVsOooj/BspQM88yYngF9vdBB9uJ0vL8JIYW3beuSZQaA3gQ3Uy/jGZON
OJSTEcZEby8zcKQR+r1/TobIbi3/qj77C13bMkQG2sQZIi14x4+5T8QaxAMr4uNg
+AdCY4BznLUTUAGIDR0eL4qK6adI3RNIJNZnekz6sfBzS0DYViywa5X25w/eAW60
/a9JQZvQFc9iS6IIixEkVBwjNVMPifhM+Aots5bzP5UEointKfKuY2mFR+W7b8R0
CIShck1xUAJvohUQicj3vaP/4VTSFHFtCrpXq0GIuOOgY1dyrNzmPXBNHeDiTuB2
LMlg7qNYA7lKAH1IsyxzPWmCM6Wjx/HHqRfO0OIiGosmUhDMIMsRf9bhAct1c+9t
GyDbUF5WtSEDPjtco01Kjph1cxOTJqAosOvirCpfxvHZrOzGq+VwGcVMfaT/UXjx
KQhsNIACdkgQOojKmcAFltV4qrs9EVgMPXSoRquOcqAQxR7b2IIb978QCehEmbkO
YfPQjIpeE9ZSLQTOwZmlPieI6K/WG/42Ibi4btT1E8nFQlNVAtiuRWiljtIKdcb6
FmyNgNuPJRqy4xA8P89M9H76DkRW7OUlrL3m+XpuzpSRB8zXdYSvt5fdWXq9Rh23
mepJDZr0IY0q2J8ZRILhZHBYC5YUw34xx7Ah8WQL2xlbHYxiyGEldG+PW8+Ls37X
OXzKVze19hTn+sq8dawG6AS0YSOPkmL1tHpwbrJvpWZnXmXI/w2Ns/mawYdC/7Ti
KxCaPLIObLLel6R1jnFxKXRrQuHIb7nwVQd+1oRZMkcL8RdFjIEuO477b1lzb3Iw
/m79iFmKjbePor9hiCs5zLmsthblwbQxhTCTt4zArqribioEvlpIXeYBw5+hyt5p
Gd84bbcj8kWZJcBoaGOZp7l1KXcZqcsgTZa+1rt9d+AYMHwc2mM1VIvqOIby5ixS
Uu+IrT9c4iC4cuTri8zd3vxxr+6ACkhe70Gh3Wu7b07I+GdSR2LMfn3UuhdYL1Qx
YcvsWCZx2YnWZh90nsouBCsQeeW+VGnuHSXyYBsEJOVUVPTTrluLgpeQE2Lpj25Y
kXZ3vv0AF24D80XYfCtHgzqYmSIblUgSiWmZNkl8FQ7kJ/DLyap/Oepfj7B4da9H
/dIwfoiPbPeiuZ3SPoUoT6qNRYvLlgxA4fjZ5IiVKrAcRwrXjCepSOQFsi44yLsx
pR1Fo0nVOw3H0V/mb8WiZzOgSM+BDiOrMLmZlnArTW3F+qbQW4Eb6NZnn/nyriOv
cbn3G/2cs4zzmffC9RWbI2oHajwEuCiR9ql77Y2jq7rDXSFX3tefDlnpKz4UZg36
mahHva2aTppQ+5g/M3Lxpln8UEyDXhQYymnNmTuXcblA7Cd+DVXixCkyomK3YYnz
zzJ0Em0lWNuk+iDU/d0WVnqfhMS0gT/HM2fX6uBbnS3YMiBOc8haxp5zgf7hS5fc
dJtsplaPUrEkc9dHPgRKE+w0D+VfHhnz6kT5dhu1FecUGMIlrWfAHt2KTda7Jmq8
USW/8o/05NJeJ2pSlXDP0uizofwu/fYIePIUWYI9N+LNBceRzDhjdjQp6639aO9s
M4Rhgc1ssZRiJDEAk3lv95AwgM9DUGQ0Gp4iptHq7Ub+G+FOnQiYv+KMZK3nbiRX
j+VIhGy4cM9du+Nt9yQdHNNO/8cn3TdtkxD0TAT6a08YvhQNFVq/7S2t9L1y3LLx
jT96joEYHwBY9z8bxuuV3v25w7cjm8PFKFh2GUwccEo8Kcu/lQeV8HJDRa4Yoxcy
kMZM8haDD/5f3CAkJ9Cnd6DlZXoXxR2CAspMXwxwD8I3ZqNw7VYr7kJYuXx5Gaf0
REbaUE7f7TmfxkHk/JLFnm+ud7hd8IqLLXxM9qEs/Z/KdHlEa7cBtByznbl2/XLn
BjXiq/48j1d7WCIgyHUTG4pblqRVco3BckUQmQzDKG/8IRgQlVkvpjSxu393nPTy
KXAvAwsiYBy+ktegPybgGK1wrlMAaRUeLh7ol0aE7Oyd7XjXFh3iLhDUNSQO3VlB
VNqs1UgTSOgFc9b+0U9NfyuSJbLm128Q4Z/mvCQCrdWsyc/y9jVbY+48gaKX6bXH
I23V3kCgZFi1q9luO3jeuuHa7Mg9x8dWCh48N0jkIDkTc1cfJSkS6laqlYPvKKfe
eRlYnNEfR7FGdqhExO96SeQY9xeEwJ+PplRExuGBu5x+/XK8IRn4G5rkgUfpIUCO
rEvZc9f+zP6m7VKmwaNNjD11jpqpJgaK+riFcWM6aadvKQg5oDOXXWfpvtf71Zvi
2ZqIJ8klQdcMaYWT27dAIl4b2oeVMlYZNo1E5GMtl1KgfeAQG+zKLQbLTVN0CLgt
hOo2dmcaGOLt1eDSCFYLqSRNCSyqI1CzNA44jp+2e8Khp/Dc7MxgLcuRDpWVXfF4
69CV1QunMSAFNzZPm23R333xxirDXWtuDWxvlKRD+51m2rRtiWYCVyNmN19JLsXt
7to3zzjU3BhqWqj7k2MvcH3dFqBiVQRlnQjZfuOCU/bk9PV2rvqJlNP1WT9krEDn
uwkEnL/EzqeUpg265cNRMH8jlW/9+iDyBMJ9jbuXEGmqoV2dmo2xZ/ZluspcKx3S
0F/BNReT5lcJjUGhie2YWrg9yY8i8HJbOdm8XKWQAMOOPfUhpTT02X4yFv0H6OdL
yyDmhFl9thlHlzuWho6YMd94gI+Xm7Y75+cXBj+42i4HSnmgopzCEOGYYWoj67ms
Tz49A5aQ3FiMzVsM2G8mp2EqF4psfQ9cE53sjMy1MtE4YIocT8cAwpIbu39iIRkp
HZYb2zjUOx6RezzSLge1xEblabYwtAiKsdXr1iVGOU5WWlG+9stCcyRNLnuNp1sa
O/hthk51tC/L4Z9aAmmEKzpGCxLYYUguBlolQlAa7vInnT0xzB7p1eVPErVS6rMS
7PHTHGf/nkLS/S1KsWuxs7QrjdYp1LP8Q1bflRhIMqYTDOBsJSdQjsyRdDSOK1VS
TmphwdShJbZVgx1Ws9eyklzgUEUVUP7QuTg7U5RHesb6GVjgjGZbR/zDUAiGo5iD
zoHrdY4jDVQl/CGLheJoor+Thrgx4RlmIwFON1Ck5+6/VpEg9szkuNQ95zI1ZERU
hrS08OAODs+pD8+UvXCPVscS063B5AoDEPRgPIZXrNDGlLab9Wa6qi641hk8LtBv
0BgrKon76MWoJ3Ew4yHHp78Ssgga2wNmRX+BX5LzVuMoN/iwARrpBNftsu0jazv4
H8qi/mA96Z79tp7DPrZbezj95fJ5zgnXjehERJRRJ+f5pGsVC47Mh7dAYbUu1OX9
Ch0gtQYTbh3F/qGg9SdVnwQLtWlyZB078Sn72Skfte72hYBULBfCnIW/fu8x+BCz
Af+RhIJxZ0ZhruGsng8U36trJlRBO/cl6uBgyEgg3nB+Vvy5urBtC8AdSwvsjxFV
fppk/HLAePjLjKgSgqzbcIvBGinDKvtH0TLf6DEMOd9V0fkE4pXTDCeRSztlk3Gp
ekIifcFyhltHSwyH8qDPeYGmGB0J0+gV1fhVYbg95pPt8CEYga0KfSqxFpC7ZFcs
EpZBHy9E9IdzNfi4bjt+CdFKEt6w9p5m98mqyQvCeEcLl/sKmSG2ynkWYl6/0qUR
QgaCt7vgukz4DGkVPDZL8EPs3ibxvM+Koh/szTOmdLRQEZpi0NOMkeLXTqRfltgI
Rp6SNXgjUsIoL995yonhOn4GRKFy5tMMk8xGtb990wwzUfM+hj6G8/nl1ksYVO6c
i0z6q+Cd2PMl6gLFmV9V3UuRQZg6klOdIFdcY+bQ/dbxQg8O86DWZC7L8Omx80wf
ik18Wb2ATB19GALJJzXIflfo8bIUE5VPOYv52vjxGejBMWCAkSJgzGQ26n9nmsFO
bJXxnvLVWwMT7RWNQsTX4OYoEiExgKeoC1Pn9PeDm23VkBBeTyOFX/MoGYCCr17v
aEoqwjqn0ILkR54yk/gtLR1QvV6AEQD8Doj72G7BH4JvYkWoDaQu+fcPDP6nh2us
OCh/PKh570Nb5FOAQfqi5K/8t5GfWiEUOvRLdgJKay1NAM2QQr5osuBnlOd5Zie3
GKH/8hxTRp3HJaEw860a+2LluXNwqflsT86QdYBFUazVW01+WK5tq9ZFFNfcqn7Z
cUU+48Oo9ToI5m4AgYPv0+QYB5AlpcD7cLbl7J2QGzEz93OcXqJJs9l9MdUc9E89
P29fKr5Znx5TBnU0dvIFe/Jjh+Q6TvxpnQE7T6+2ZuaCKZjH7bD6sO3k5KoLM4yB
fZygU09pGqg22bajUVMvsfRK59Nv38iMSemhyHU/jLCC6IJi3jhhVgmGvFeBDFEx
h9bVhPciBPBQumYpuFy0qNCLIwstGMAsdsfTvgge6BCVGBQESdRCxlJ8+FnNbUk2
2VUmskk5atxywFCgvL8i9nfrrSyBOtdmNswqIZYtvt9vDLjJpTJl7En2KYvFfvHz
uBnCiwP5DrRQHr5RGaTi2gfNyUW/PmlzQkhCtnmwDbgavfhMoSwxuyCl+L1ODoIa
9/90H3rAck5zRdz/0RQGdOSmPuOXtDL1EGir63WJLNJhZxyyiT7eqS4vl+MQLI47
y0DIKIh5Sg0lTwDg41CLiHnKg9EPCV24MssJdijCPJlBeZW7Fbo7xMBtfX6fkLeu
KxAX+tmo8cbbrmkkbpZO5jxoH0T2p76ZFl4oJrjO3eTpt+FXHGT6EUJFWLP8BLtN
83j2a00YMfEO2I7f2F8O+iRz61NTYhSMhzU6VrdtyIRJ3G0d4Ya4JiEzRxyc3kkf
ppcEhvoe84HxnPak2rfHdkX1a1VgZLjGHKhwOenQFdm6JI/zsx/0WaZvXjgtHcJp
DVTwad9ssAsSR5D3xlTIquoYSTFLSEcCf6Vu+stT3987P+yRnlcNJaZJ34+SCS0I
sFPreI9zGRNNAKZxbcHci2DHQvdWsLmsrSM4Og8J6XB2NC0i2Y+7HdraB3WaIbE7
27E50Nej36o1DzmYvTUvgjIFSwLkSa7rM8mXobtRCiZmDFsnz2YK/3iZjANKFcVC
o0as1HN23X/aQc1hBo6wB9RG/KgpuWCWrgvwmNIECz+B42IYaEeCpZa+itLzp7gf
LEyxAR4E9QLpn6pq6NlHeSnkNptE+/RZqVCTQYH/y9EvF3TA0BQwnMjFeHBpkrXA
wSqu9fkQqRebCq2f0Z4tk+Ni9LX5dEQTbY79T9y42rjN78Bt/feuaN4m6Ddv6unv
LCX+L1zHbQ+CuSATTm9FG03lQw5rKN4mhNydDvHsnB4IcHXqmJ3o9iZNdvf8f7Fj
VxSchAO6tVC21/jXhCp8aHroH3GOvguViGnvWZJ5P12zP1eVABcPcjMz+ytW88qg
KLKE0WgQaRynK0lg8ZR+YGu8wIdqdFgcAREt/kGF+uiuHG5vmLOp42YTcap0jcR+
/cVWIAP6h62ZUsXcSW9tOswERbE66QG2aPZCyc7BB70ZvrTR+AJFyEnU1KHGHzv3
dhtj9KZRTjpS/74xcQ6PB4s7OhyuRwWmUZqMMcaFSAFbc66N7y6idmn3MyqIKbqf
Tv1L937M0duvtE8vtjaJ5Td3oZy8zRMYaaiDoAssCcUeQvGGYvb1kA2OmBtTwaNv
YzxongoqlL24SbbkVXXVtP+lJtPhzrBtUE6I1m2MQgrvQJ1zgc97hcm+rXfiGLGl
8KkcOFuRrRBs+AQ3zQeSMnmWzbdmFQwioi2pWMBCQwTFMkB8D1CNP3CNUgnDLVhO
Micp/gQFQ3I8iUKsNEi1lATmtMG0MCdaYLuM0O4IG8vwbBQidi3DLT6GxJ5QKaMA
F8+Q5+gbyM8wF4+FyfGiEj4kD1rtY1D6dYPVe55Mq/9tdibW73WEFB2Rw92SL8Fh
z8wWA6nq8zV79RqE5GuMmrpD/ASkCAX8YFJDA59JHPn1FmpLzrrMFBhV8UxeeSs1
SYAULdx88cHGGnbcl3VLckFkH92lDVmpvvaSeJ7hqzqovhcmh3oOn+Nb7pG3ETQP
6m+/q+fbNYrg7ogibHRLsV2QpTcInW/9gfg37FoIPtA9PMUiOAw92GamovT2i5Ob
eXc6kIkcWGa98UDtwtWX8qpnSU8lIrG2kTc6dhNtRdIBLib58T4OVmsXMC11/FpU
bf1vqGb2zriudACB7YGJMfcAe2/EUl/KtwsWPeqQDQ9m8LDebN08y/xAomDQb8iW
MQO4RcU0p0Xbx/s5bnTtVc7oA8/KGMDBpRx0r4A4LxDKt513Ze2QWtzc/wqUyvNt
iORCglRRr4CnxnpgzqAljxy+1Hh1ch1z0OxU9GZK++4qMjpRW2jOMv83N+2AjIsQ
IQ29bHIZkLwh3wy+pKFs/v3xDznR5lAnZKN8rkLL5uIuIkSYDk31B1ArQ2JMDV65
ou2g49boYT8omUDt4Kx2ThkV9247m/Yq5j38JlqA/Ug0LdydBp+fQSiDncttGiPH
/Azerk65FJ4dcy0SH8MvffJhEMG4WTchjS6j899MfZiRn0N/v+tvN7aGv+WXHHZu
4H+uSnpzRmtvJVEeCSxuU3HXg9IUkzBdulzKftbLSvGD6x1madIYXdHUi847Yqm0
qZfMPaYM+RywMV768ACi/EKAacyn9rCDwB96lpD5Re7NK7oBrk0nElN7w3eJuOYj
xCEC8R92B37IpNbs/96tnvkWrODPu9S4HotopMMyiyhKHngFIydLo6tn5YalbtfC
yq7lQTaWlThTzo97HxeV3jxAEoZbWjqUqSXtJccPyDY9fN+LD3K0hsoRdJkGTi7I
JKF1597js9I9A1AZVc8T7sq4YGCD4ZMVdzrZPWSqvkB4jF6eNokc3+kNmCHSQBwD
InJeMYnkoYOjFksmTQfWmdu2xp9EPXIId7Suhly4lYGQpQXL6z1/7B6bLzHVumlW
yTi3PbidtC2GoJ+NyhsYcnmC7lTwSwwZXl+1hr9ninY=
`pragma protect end_protected
