// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:04 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oTmbVMWKEbrH52Ejb8+LVvutZj4n1//EPoFwnYdNrFweyGiBkDpOhSDqbiPV5Afw
q2Xs4u1hmVbIF0+VEW4le1nWh+D8tqlr6ZDLnYc3yMcxJJ4oewNHLxST1twPpfNo
sryAGCCL95K5gV2j+QIusV+aSz/A4K8xgq5wQ6WvtvE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9984)
WjyxnizqfiboAz8RH5EenuWKZPOAphHGqH8TqHqGK12Y+eqrLqLTR4zGlCp43/jP
ZMNRX3ayIHggpmBCoOXYKhNQ7fCzbb2GjQ8K0cJ00aturmS57rBdeqS4Ml6pKJZF
WLGfD0SgZ/AWq3U8JTTBRXmvVGBTeTDNrbAk58nL6+mwd//7vU4iMn+fnxcg+ir+
84CkkiLSS6a/qDc7ZlAHRNz8w82NqPv2b4/soFm/3ITwBuPAwBGXzNVAaGa17uH0
+MZapTdtSGOIFbYnu3SmRo3PQigjB5O+mIKskVC9/zEhkQdz4TA85B/kVg/ZMTk5
U9q3jW2pZ0fS1rodMK+PNUV+o3Jv2+E9wFc+AF07e7lAKjCZpwo1QGSvLhESjq48
J6oM7KmHs2IQqElRNmTQMXxtgkdoA7/MAxvH4gNtTcYlH9t+4WQ1rIEJsJ2CtgRC
s7tgriCcnfrSWMyyZeEmwBP25NMW+DuhJciBZdF7OQ8CKYOEKBMmTDJDwXXjUKC5
Mm+3x/NDQdXqo+/Oa2pyOG2VjA0raDbewIaT7d+GUSzVO8o8lfiknxwYeBbDrlA4
R8OuPtJJyToQ8i7Tz3s3WD7Kq4QwndSakJlnIauJTPZ3BxuzdeKCMGpB/iWmlp/V
RhrtMYs8dH0wGfiB3SVf3AqQLMwkfUjkuzQypqRHeaaKq+V6zh0VGRgTVLHHSnze
3VHjE/Y8C9P1T3v08llms51vKm2fDy+H9oydNPEreFyX5mXB4rjRQSPb6KjZbqf0
+taziwraVYaVJN1rsa4ITQHLPdZuAl/Eg9g7S1j6GSfKjC/blPtQ7XOYaNz+E+eq
1Vay/rBptRsJmw12ydg95zo6zUjDGeu/focXhQuHQS7YrLN37vgWw+lKmeK2k9RD
svAkUcHkbYVzsTLXYV95HX8rHCbKZ3xOZlrZOPJQXNtQE5mzM3sdnKjzF0XOOACo
7pY0hhs4BagS/f/LBRpU7cSHmeIHm4XPY+17mvyXzgQSxCO5nXySmy86PMdCtQGY
2XASR3kq0hfFWcL4g5m0wguKLmedlQxu3uPhq6S3sZflzdgpjeQX8RUnWnfi75se
2HHMhRjvRrHf9EmWWVwx8Ew/DghMs9GUAYqdh0oFzlOStzhrGgDrW0gIPPtRaAvf
1F0+rLB/+q9xmqz5whqxSJpG/ANKOmghwyF6A9DVG0Pq6uzRWEL/e5inLadC6FcI
DmX3msTn8YS3BtTKYDDoumFPwZNhgZkxzlSpIlH59hgX2pADo1fuQ740b3c60FXr
J3UZeub35qx5ntOq2+jK0wnyzS/X7YeNrOYdpa3RB0lKZGpsKlSZ+XW4H0AjYdEG
m3wcZrjyATV2aBgOkIoukZopqy5q6hhPYSpXbEFNqhQUJNuPB1azt07RbtdWOave
GBCnrqu+kJYiC8caQWaP+vTJVzYWqBJM6u5bXlfWywqou0U7DtEaszNLmTMz4CUr
ABbQbsCDwUAbNmUCJnl/CgrcC5Y32T/9BQmjDV3oSL4r6MM9i8LQMuVzbZH2EXz7
IB2d8WQo0TQBX25KoSw7HVWkO+/AfINPIWe1qcViBaB9D+kg2Bfqeq+/8PdS5oSp
SaLHVynfjMRQ0PtC4PAnyLvlQo7783BEkYux0sWoyyP7mhVYD1qwo+PpfZwvJYKW
pKeElLIWKeKyilZUMJKTQHK3PQ0CizBud/nMRW124/p6CHdNDytv7TbYGdRsfAqq
wJEWLHP9yn2elK0AMdmX+jGNUtvGqxkrsg0B4DtqCuTirC6vk6JRDVhbjhjEdzgD
arh2HkFtw5osiqySTfZXNWXQiKRId9KCJZwtpTrYBJRMjEK9hH0IAVxmpVdWqP2H
HgDR4QpwjP+A1smeXr4CZGYQJR4VURlmV/r6XtkRJhJFHNVbB4ER2zmL7KsNbhVV
a+W9UBYNEI96ZS1fPZcnGlRTwJf8usMaMgdtR7dll4XQJBfjeYYBfWWE5p9n2C8v
B7r1kQ2nGKiNEMIokjfkoKez93HnGC/1/dwVTr44TGtVGnUyAIUHwEl3AFFCj+h0
OF/7LZ9Tf3Dx6zxAb9o+Qmc/U8SIVb9jM4t8W6M8bCgsvpte/kOwW4UQHPFI39K1
lAi00pnHEo79X1cGTdzqBdFgBx1tOnVD0HM2O0fL/nF8BDYTh0Alr+nJpFaOi5L8
If0KVgFMprFubViBU8A+hGuCFDUCbWFA4SNRRXp8fpFQQ0hgqV8BzNEImCMjpQD0
+K99Sx2RwvZ6/eZY/gQJ9trf8U4r4Lddi1qRK7GOhc5CiP8K7fcn09RDzW2eXTQY
IMpwjMwk9emPtew+v8imhabvWDvR3RWT7QzHI7xfE5ONFHnGvnbJYgznVmvA61lv
+XJRj2zpcROXammkr3FEWxDZ0VyXuhYkBTjBY2wNWwShFE6LBCfuGSQqTVym3gWn
F82wyx6nycYk1dLEQuCxR9zQro8N1L0aN5th0qWe7k6lHI0t22LD17d4+ZDOrnY+
21W+EAB23MzRhfxYu7cqKshy48coLxY9ojMQ/ctYK+R/hHYJhAl9TFf0ppdzS4cw
7oQsib9WS4PW8mt+hFD4pyUi+r6n4g4mu6fPHXgbjDzhkKjwchLQU6RqAQpNd3MG
IsjysUWaKJ8OTmj4EEzJJqxuruZ137UsJsk7icmTZv+g35ujTNbAh1V9ak3Kco9a
V01ZVWJfUULAI2CQN5MauPyHMWKFC5NwQ49a6Xyaou5oTh8ibyeojUZENESFejz3
3xQKFvZBC4lryKiZT799De2uOxywqE2GkP1mva5kclYwvTBXwffC0JN/HPyhL0Ac
FLd8BWiL3h1FavRMFsvwJxy/ECuZ7HsW6O8ZgoZNusiMTQR1hIej6HWSRdeBSBfZ
TLWaDw6VuGoQr+rhCwQas2dr/VNay98ea5UN3ggqFF2PigB/2tcrff90JGzbZPaN
P6b87Y8F/l8noWikxCzXxX6kRPwR9+8YzxLZWUo8MAk950VVspyw27x3Ql0qSOnS
VpbDEuPAEvEgjlc+8u35U3r2RiyVe1Rahz+mwnzyQjL5TGC4MBnx3UWBtdOy0vML
dJu5ZLlyelOhH9dLMCmab7W2LFHgkD6n+4es8fX5k04OVT5N1FPfbjWZSiCu52+2
foCKYw55rTfqJer9YeO+ccalJtQ2ColTCMyFgJ4ysGy8wxHdQ3N2kpac98KoEUdg
E9Ih0abcxB6uHedFnNkSH/WnfhLce50VxOca4Kv+5NTXskL3FEYAszAnnNQXFaSO
f9Za9Z/mj0k+2VW5woU0tXCFqbK2O53GPAbAOTDT/0XGWZp70q5dhwqb1ntq3bAa
Lya96HgGZ4Df3i97xRsl9FypG4JYUIouP00S/YCh2++JjcPHFGobvSO7x/dpW2xh
UREDLIh/Q0F4cFYiU8JVPatjQimTfitVWDF+p+FXPsldlSesI6DPJze7MP2U1tDA
MXEHgTY/bkk7ZI/ALpg2Ki1szmufz+GPU7YVXnemsz1asUiDKLFun955kqOkXi7P
VSf8bA7we38wYSAH1eznlrdtCgpcJPbWG/e4BIfPdE/85v/6ejIW9H+3yryq2T1x
aiIzovVLJC2PhDOTovciR/jLHGCAMum8+8IPJ3bR3GD2oNhApsd1qtIMsVvcIPyZ
muVxZpoC7Ca/GPys+Reon5HeLk9e7wOo2HX3nr1I4hfI0IcNzPToBaki/qdXhdRa
G/ufiCSRDEvmeNCNhGyinRvlNQDxbUNlO1+jrIWdb8GKKs5dwwPR9jh+owrY2g06
6+GHcqbDFyDurCwFZfnbcl3vq27kfHnB+KvTfcCZu4sPFB9cTnawb1gYtko6I/K/
mPqMwSj1TpjNxa89wyoYh3c2SdIEcEl+yA7+8VFy8DMPUz1dd/eHzq+YewLcx1gT
q6GOHC+Gz+JVThsWtJIun4AwSAxspCdZkGAn/HJCL8BpRTtGoN3DT8dnvU7U7ugX
q6ASanyicaRbrURNWSyPGQbMC2uUhtz/4zxX4aKSUZF8vSkia4/9MQOdOcMWcyxJ
02ZC35ESinbSDWxCa99bSUU4CQxMIrb8kyO6gDvqadUToWnQ313H4hKmjl8vaiLJ
SURfbTXOoqSMza/44hKc2TZX5bLRdzJVEy7l0FOrMBZquLENdcu8FLz0keq758wI
FBliz/iKGdpZZO60c0yvoNDPZDR12T2tVVsBnfdeiwz8/FAd3xuSroHvOgCDeGI1
d/7DCsIN7jUjixejMFC5kVsjfA69cG76tXZ3itDxhQkAxfAYtGj5dT72FlmW6pOW
ycfxHOjE4YRLQKII9p3hhVyMoQeaW2479H1gKBmPU1gxXMtywu4eI58YypOXRsJd
A99itL9ZtUFowan32SYhf2i2l6PdUBEsbWoN1063SsmpKihQI/7lH4OFBncWBOXE
nDitsgMbavhymdsUJIntH8uGvY23zE9dbdwa92fEvEl6be6sGYLAwgpxaR1M5yTM
oEj70AHRrGhbrF1TlZrs47Z9icAhhgy0ecTJwQNnLC2WCrhv8YefxTKOnFA+Zb86
fzNDfNwjtyEEJxFlHozoFtC0Be3NCMY0SuuHrpOom+hiYsrX3r6uv+Sl1a5IYd0Y
J86yvtJJP/BflwDx53TMfI37pGC3vGo0usRmPISj1fKbWSVA/JfZ2xGlwrCTNMIp
j9a0yhhDJoPvDRkz3MWfg76orKoA/yE4kII07SbM2p6xPB8I9aN0JuM239wunvds
hKL2ACRsRYZR3+EnBJT9UsmcbruiCjVsLzzJfTVJM5aCmaTQJytbEQOyNvXj9grp
l8GgAxSa6/9wq6shKVBhk+yY25DPQ2z0q5l/wlq9IwV8vNk73Pxxk3ZGJU/cOZT5
WOmhEB4lkfTeT5oWZgAs6h4cEP9Nyo4WkqZlk2Wojwjo+2E/+10JN/yOZTM5YRyA
WqO2pd5otkHS3AcLBBd71mlhnTSl1mcTQeyfVcyIqSMW0rZ5eFIxV+Y9KMS0a3W3
73ZT2t+2ZV8CQi3SAPp3Cgv1k4xj8BcGkJ4bQwdZdl8z7MBVqSfiBDYup0FbHDgB
aBc+PPiV2ZfaYUsDSdqNw5oFxaS037rsmgt6+Ivr+6CJ8GiSgasDCXkKOzD2ePO/
SClS4FZoqHrdHinZ1Hv+XUUG5V15VHD4cVEi2Z42BknURVT0UJLfsVmXg0CPUatJ
x6WS9T70lbc/0Zm+Alv+lTyKKtffeSVopRoZ/V7ek2ybRUrxh/4DowTqBowpWn5Q
lXJvr2AzMWpWCGdP4Fhu6SZCJgaFfpUZp2Zax8fipnh+92GAXC3jEWJAp8zI/2n0
a6JBDkn5+aQGbMufuC9bKzFcPabPbEGa23Z3TCnaGqxvFv744vrL17ZTgtkp9NJO
pjwPgopQx18mNavp7ovDIp+VyYed67Ut0gcAm2yzPG9ZvNgZTimsiIKVoHaizDuW
AMVD9kz8gL4XU4fyS37mesoOkw7zMcHx+M50XJE622ltSTTyoJVNSWUP7sEp+Wv7
FPpCXO7GI8SxtTOXh3yTYyprHQlz+hCdFr/bcTDouxhAV5uVaKAdMNmzF1ibof48
qBhXIvtuzt+1BD9+B6dnLTWCVCDXM0Lx8851KhaONZLMwk+U7mgOyMh5Sc8E9Tne
yFol1exHYRjn6KZY+er/yz4f07T6U69W+N3dTl/W3s8PX4cCZzTctB07oHEBDZOQ
D43Qc9dtH4xaCtBKz7wsJAPMpzA+5Sle6TXIKPiij8ZMOE0EgaDynOHy98wo++hp
ntducAO3GL83fUhtuKG1Z6mOm4AD+4FsuvHpc4JYDpNesSnDEDoo19ozXJbfFfAQ
+SoFXPuchLG04XeVET0RF90kG0T8vBBWVvbS4krnjb0IMDboswPpu99raziYboS/
PlfWEumJ73fJGxWbqNC7vm5iksPE3AJiSyLRcW5vyJ7JeM6xiTaCDVATOVEB7o4H
tFNgmGvXZZLxdENCEubp7bXtk6TGjjU1ZEsbBALmHt8VckmOPAYCY6BLhk3u3N6c
N3eHe1b/6HC5m0x7nsEIi22ynLxwUYMH905CXGpxHweyyZf222pTEry1r1w7gqN/
u3/N9wqy7MiATBMpLxhGlJV0H8i6MoNOBPXzggyf12WPUX+z9lnIkpZ4KcNrBYmK
ssQLJwNAZCEwDBJSYHjQk7rmcFwWGmtoGhwdW6DZkHkJCc8lGe+TNe3CnQaJZsnH
5PxaFZmQjYEdSdT9bt1vSTiQdOFuxLsVB95vBkXHvlmfKnKIEU9OiNQ4l++jkuuF
1ZO75I68Vknye9hd8jiKtKTG5N09WLffyjnsNlgWIOEL4xd1sN9sCftgEmoDXkZJ
sv5vM9PHzPFTZEGsAtcbgItRjNQdsQTvD/unHqTzbY1QOjc+Xyj6TkaiMvFp8MmP
/JXrFOXPfSRENFqVaaQ8YWXMiqMupeuf/L7cpNcWLpTumPpEE9nPcpCdjLXE1875
eAPJbyySi6ytn5ksoTgx0iVoW9uJ1dJu6xtiumxJrw/9o4jVyJgFBt47r+G8V+kl
jLpCRluoeTNFRXdM8oV9LDLD/DrYFQ9V46/EWdVR3Sv1cdHGuj9WGtmlLgBZ5375
AQaZCI2o6xVV0SU4XUaPr3ePwLYwEXeX3EOlddTiOpsJ1HOsXMZCCpFMqA6qehyi
tuxYZaVw2hfMhNHII1iAy/Pnprfgt4z/6rwqCSFU0LsGMRHwmUy6W5qISCrRgXFV
5k/f84TKX8Trxt/juGqXHXPKJx/7N9yEni59XAy+Ajaf36/Ok3nrS07DGwnl0qgC
5zorhsx737Me7JZ9nUaNYpu5iamrxClDSDKc6jGggRcc4I9Lk1x/7qIZ6NEIFZnU
UPNUeHVVNoRfiq+V1lN7XLUTBH7cHOvBz7dxqluK7diIB19QS3r2hIn4X3ZzA2+B
6BhFCd55v4CH5cQUe53Kwbrer31WNGyVlGQXz+YAy49d/T4tRG1DXfiuC/xutRuq
JbrTnMQ17TkDgmNZOn7hvNbruF3L4RYuESdZZHbjxn/g1Zd0Fc4NKX6xmMIqaeCn
HTTwEOnGzN2TdGwZTiRrU7S+LQ/sQSBTzeH2Nih3FGVwPtK64fiDl/2Qes9WkUmn
ajMM18JF6LTrHpSr6H7q5A0xNkSOTvSquzdODWb1WsIp7/jbstWLAG7tt00a6Nsq
/U6WGQLbSLW1xVOp7s0L9p1HgXzY4WJCWx+AmdjiuS+/oqUSmfjZQrfvdIcUQJ92
gC9j7DQkSxjmgaR6GOF3O/2aicCgCGR0k0ORT3i34/sm5BT8Pdg+zJkK2xdLMWk7
kdRvf9AkjTEAYSv64ocpS71QzS3TneC1ACrDo32+hq+v3cysEvW/JGO4M/EBO+J1
YZZ1oLd6vDeWO5D31p/PVUX/YoNyEYEVKdPsFFYQZPDDjyVIBuMeC6UsNEB2QjnC
0WirdfUMZGlH+nQ4MwcOpJ+KXIWSGSd4om7RxhtvT6oGDws4Vyqxe76TaAgtB2H7
eARXGH+LxH3NkASGDv80WL7I69aaN5cb4SMFM/VnjHTX5Ji+Dv/zqSXaRzibTzOL
7FDH9DAzGFSLz1b4YedV//pWSWgnJtDowCYayR4b/NsIaJMM1L9Ny0DisMv6wKGD
5wHsXLuJo5Vr4J1Yz8Ahd/gYfCsf21Zgw97to/5eqC+8j5DqgH+0HV6FBlGrqFvb
D5/m2kda/YiWeZlpNVPqP66w4uSOT0IB0NWTmjoga4W7wzhP8qkVD+S0XJVtu65x
YvVhkiUDIjhSfkm8NDf23Go0gIwUhDHbgmFBrghzLv9uwqawJyWZooUw7OL7AWth
GzF3om07sgivMaaMUaW3dVg0V3O4dHnrzgMx9UOzFEhjAcuC/L6Fk0/nrS1ZmNS1
EzKLd9ReNI18ST2s9HwWEy1hBP7GEmznkrcjSxSAG4U60SHfxX7GgHWk41bjoYah
i6SQ/cxyiHssmDy+EtLAVo/sckAt/pbFanTtAWUrpc0bMvxLVT8zdQhyKhfmR67R
xNaV5OzPE2tmVBU6VhkDECQbKenpbLJNmxX8OMzY4a1KcGMouNr9rxiP3Nr2uvKn
HJRrOA+K3P8gwK7GPkOACxsLepiWXFc8KYntYLonl6E4qkB0zZUJ4MWuIpGnKE/U
WKwfmr0zzP0dYyw00vcwaauO0vAIgXxKiKIjCywvOZWdV6lRFuH63Jzfhf7z1bYS
teOEioK9d4lbwJcU4bx1fpKiSZtO5WtoWvgxCsJ8hQg2BArTErrtoGG2wuuVvpBI
Y2saakXku4lrDsh+x/0QADH7Q7FdWuzcwG/+9vZgySyMHvPdk3WL9Du282/cLQ2R
xvn9cA2lKpxiqWw0YmonhLyznpupsZCyEExuxJBsF8gCYkqD8k0sLK2co8++/IgW
FX0bGO3TibZyKjUFMsjgCHLqYNQSxSDSw0vqd8q40Fxn8wQMdUaExagVw04bY/cz
cm0DU0P6XhkTEKkSlnfJKN8VDLejebZ6PTdHS9OaxnKNfk38Byp3BQdENf0GYXLm
S4Mi3NVX+lYmHCmunNNEZh0ra4lS/hRjGXtfFI4E0q39N1rkQSuwSVTj1Rl0aRP0
NTNpIOm/1lVKUKyZ2psHGO8V0245Qamy/ZnAx3/UdSyXAMVVzZgK+9pCQR3W6Ma9
p+uogLH2ETuvjh0Z0tbbesakWNvoHPwV9Jg2VDSyjC0WJ1gaNDRzvBrVSaH02u23
BpOy+ubUr9Diy2B4MKCEd7/iVLxWV1+9LkU3HU5K5jep3uHn6okMUMUO4oQuUD/a
BHkA+yzCp0DPvYP11W+zEPDaO9w0N/2ukghp5rbXCQe+4VD/mV1thYRPebtE7Abz
mbbnkbtF9ov9hID5IoBzdtSewY8yTZbwMzrbVOmj0ORxHWv+Sc4DpxmJE39wkGRe
j5153Pc2IpDiILLQvcwL/6kaLrrYIt9MURy5MD3xXGokzOGFn/9fHrpYwvdlKPB7
FuRczPj28aC66iG3c/Ue/AnOKfUSsm1j1Xee03+JlxiFYFnwDs6JzI16PF68bcoA
Ovw2IVWtP2NJeO9R4fQcfy1M56/2F7pidgNvdtCB7OnW4UXg+Gev3YwOck9lxzmP
VCAdlDXALIal1w1GryMSJkLgkwPqBrnspkVsGHA7eDN7FMZZWWKGtaRRdCxX8zmj
Tpd6g3iNjum4hD/9I+QtKzyvc89T/nGWyM7cn7P1bFO7R3VmYy9EpnKs16JgPSfg
Eu1TvKv/h5PBQZS9SsW3Oq/juwZ72s1EbM6hKMAZcUJ0VE3NwhiMIA05rQB6exrV
5GyFAnHwodS0Ya8MOsT3iQnzjijk1xU3A9xOJZEveWVtIS6Dnnfgd7qnkESliYHq
MXErH/rnYhPJjJaA1aAo6PsffE8SUaxKyj4KGd+PquSInO37krMffnsRf3oVeCx3
x1Gtp9L2G+kvVxvAHoolUDO8R7h4FrVfIK9i1og18Rm42kMy7N9e2uvqKjTljcpF
FfNMIfoPYvAedblZYkYBiba43r1K73VL7QytB5SScxUVPq5bLMl0XxCAZWbBMDHm
j73tRQoruRn0o/6B8d22pcvrdoVLoCS3FJbH+JEHW02oHCBc4yVnVU50vdYlJY1O
XK0hlgfXJC0/ENIBYCPpeJcRf4kzvCWvFA1aBLcdRNiJ8qCuWe3C7xx3WK5QXl0p
Y91k2IpreGWxsBXroT9DwdDALgi0DaI/T+TfGos2xHfBSUgT4K0E/8ggLIb45rHx
78LLYdtFzYXqT2QkPPMDKgQ3FPiPcNQdOmlUqXr/FnJehhS3gKCpcbmwoYVcvD9J
dsocuaBMHgu5viIkCO2TXfMI9q8pF6jlwqi3wUFaJXDIrA/Q7x6bCE4CFPdMCihk
Z/3l2fupOvOQCrfQ6hn6y2VvH4poAav9JL1R4GpI83nFmN6dj/1PLXCLEHwO6ewM
2F7Od4ITwRZcs4PDbNpE0IsbRbpxtgLVMEdCJOI0Ce0b+8CR/WXVm4qKoCw0pI4E
61ASezBL5zRvFcba/kLROfmsxDi5EgwafXK527WEWawvgHfSeu4Qr2ue0J/gB5vR
p/i0uyNLOleGxR5X1m94wmKXGXVTFQSIzncwYedEOgIDF9T5ypYEsJUT4QmE9Cwk
gpQrtfdJDfMLmNuYXAuBWpY2sYkCgCC2IPL9jIl1A2+cbuponIJ8R6VwZakQ6s80
qLgwtEIAFK/QXYxqLIpFRQxunJMxL4hKckx9sfLALKyYRB1HDGIsduwfyK/Hi3Ue
xWbEkb2JX7oX/KtRa+87EfdMuE3lBPKRugvdb6/Cwg7iB6O/RhE9H8teNS8KO/Tb
E94AFOK6obL3bbmyk8BjSHZDO0dl1l3T3bDEX+URecrveA5gcBvyD2rpAESSphgv
sMzDXqNknZ7Z1ze+DeEAGr1UVQ+Kx8s91SdqhK1AErxsYiC0nz5atJrTrYTjVAsH
IGbEcp4xEU6zXsHtGB/WvMwxLrAJsUHulhXSzQBJNyxhO7VLGT0cNv8B3vhkivr7
Qr7+ltvQT/K3Xkkj6/iFN/MjutqMKGqhRTJY5N5Ei3odwuptAJqgWchzGB351IeD
huix3dFi2iyAZjHOy5fvlXOX7KZX+3x3lAtZFs0MBS6LWeH8i1JtQxOvOXy3HhZ0
8ka/QlA27Y2oH/QF1UzrYp+KKkZGBfMMuisP4ZDzOwoCNUnJVPDwXTLsziofluLy
XKjs8/4beiMhMMYotwlsIztcfbp2eigZHMVbMutwQ8UO4C6GiJyXjg6b6N6g9QSS
F1pKzREx0J9A2wEeDwSKYC2fsm4jga3pFBHdBZwnp/8WejcgLFKwNVfa5waHCsLN
gfSu9zWc0+AYSM/sr4cuakupMPbnBCzvBpjDAUmnzi1oLa9b/7w3v5fndKdmQ1Rn
vtVgDUdkhZigyYs7yS7MikQUtAP+VAVer/PFRzilG4KkY3Zex/VTaZfLzcurSKQJ
ZZki6kWbBCLgtgJ7HjRQaYZi1l3uzq89DzUYCEwY3kS7EVII5w7LvIAYJKaWoreT
xF0/ZbQ13pl79Cu63WQAS/ghBZUWammcKyMA/fnO7fcN8dWysFzhBsGi54eA1EkM
0Rl5+pCIyFfMd3Iq0wDY1JSVVFUP4aztGakG1Cj5qsHXfrdJIs46Mk3hJ9AAw8VE
Jq2CtK+2gcmjZyMS83uXb1GJPSuxTZ/uASbQdoN6YnVMvL5u5IoVkefSUuNOoJNW
c0oy2IePJJkp/Zm6h1mLdWMnhkUOMfCviUQwmEo7umZOgmtoV/ih+FxiBmBU5rfe
HyTtlOZZQkupQZFm6P3PHH7gLIXLcT0p+uBjg/N0CAvDfJw9gbMO9woQq6X8SF3J
ipAgopw6hvA9ft2nvCgmlbJ0sBhTv0CibCUJVnTsAxY1MQuAD3E70nrgabrS5OSR
YKvYyqzrNwz13R4puBt5GAoBc/6RgwM8eMzdcuzQJeZW6/XCthBt4hv/NmZPT8mo
Uv/48I8yTK74tqSIJIi0i0WGoIsx6DjAByepLtg+Xt8bPiJRCsAUDsQverev6kl2
cX1+X9J2NUx5Rjb2uIxriqec8BmjgfvYTenqQ2ulrQAzSZ5fXCKChyBbbCDi13rN
2RyK3Y1SkTjhJ0jUOsEV2fRe548NC+WKyTY4pW7In2ZzhiiaMzcyo00YvtLPhjzC
HW6UIfmotVpT7g2A5DVyW6lHoWWGzguseJXktuiFJlA3boGkKWmavARnMWeJ1XKB
cJJE/P3Nc8sddlIVBqH6QqVdX4+oBXbbrwXWn+lV/JBo6NnSj0bsRWNvkrFbDYoX
5t1HUKj7JXBr83zkDkXwFquonMzT0VFfn2cDolYbOHm4ZyE/Kjnnor/G/1/4THHZ
UAjKAdcB8voE4D39fe9rADmEH1CN1iHInfbyrJO91Z3VAjlJS1sZLjuPSi2n6KTk
qxRwJ6SsBRJOU0l/LRg54k+0uqOHpX8srcbNEzyE88P7Vj1WHpJ5nA3IjJhMSfFK
au6H0oNn2Qof6AKmfAGaiVUzt9ev80gRtd3OVdq9aVWZgmiRtnP2lukKAnm0wpx9
JUH0XTrSHbb/BM8iuRdBWc/1Gx3GilzOmwhIpUZM/8uj/4CPMGv9EodZTTdj53Tf
ksl8hDs4g9QjUjclRF02JnRGVJ2QlP/jLtrvaIBwdVNFXQG6quX5OeKdxHY8BloW
CKSmopCUM6fExgc62noGc3D62Wl/zm39unw/ZFVPotcgWNK8dHsjYS3XSTrvtQGZ
X/qe5lWz4qtHMU+zLgGeUSvIVxWSW7j8TFKB88QOIZiskIQn32N28dhhGk3nKA88
ZwJakeeSwGMCS05GRJ5rv2s2aRvx0uZ/Ezl3a78HwIwVEmz7og6SteFmF5IBkikT
j0GGiHtx4JueEtSA+i6dR3JQaPmbAM83ZcFFycHIYo7esRgU58NQpwuKipTroNYL
Gt1R03yHLooCe1KtePX5ou9AdQhENT6KhNmdZxsi5ieplkS1326IVCMr3FYf+WZK
WZfSkjpY7dKx6Cew7rrZBMtGzgSScSx2YZaTL8Smqt4QEr16mDIoetgwHTKmnuFF
XruI9Po6CjavTB3BFHwYsazss/2HhEdXOWoQ0fRZop0bLV/tC5/zzRO1yLbHsTJh
a4/MiPsutEbbnt9rLnhXSOHYcAg0X3FnBoT3nxuHtIFjc4UaDqfHmc2gZ+jp2zvr
CFFaLFwbIHB8XLgeLvdPRYfy53ORi8/pmmRYvT/Sv37naz6wVo4dp6jlQbkgdsaq
qCy80FUS2dd/FroIrwv+muqgz2Nehb3okp7N8R838qF5fXwMkVt2nwuqoVANOIkQ
ttcrR7TZSUPujYXZGOalh+BA9xQb4lQkLHYTQ+qYlxC6lfLghmieZqmbXrAaH8fd
11ccfHTe889kYFAqNffNdl1SU0wZOMlz82cp6IbUr3mfYVSJ8zH3FUvSKBQmkOpw
+/lbb5tp40Mx2SPgyD5xswfLSEEe+xuI4Ky5ovStNHmCLiGLvd4YAX/vNWBY6RVX
6HuibLju2SbOJyAhVU7wEnVVyt5XiPhhuxFMEA9EIlafkS77JBlZLQATuTxDfFtu
oC3K+APTT6Xsk2nIMboRMC696vy1QxjveuQKoIKLksAQEpdwaGQ1vPhLMZ+JHUBL
7M/gTY3X8gvXqN/SlYCXf29vsRxp5aVpmrX24/CLbAkubIsZPCaAoXUXWZ0kcFP6
m9TZZ0k/joONfPEMSPXVNRYlMTS1mPuRgAQko4k/W05JOpjrRiLwcWDUnPSjiEFP
LthnSf4ogIt9Jh55B0u4fQ+q6g/o/Lh+2dXbKJy6RWsbzOOiRj6g16R3bJuOv1tx
`pragma protect end_protected
