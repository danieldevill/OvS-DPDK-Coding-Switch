// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pU4uFu+wyWJEHHD9550PopNxz/KY0Vq1C+82iYdREZn265V0JdwVCFuxNjLYxE7V
X1i7CjzuWMixFFGTVAB+hK3Vz+AqWHPQFdKT7mRtrL5QuVgsXbHZA/L284O91vvr
JG1v8rWf3Y34DsJXPftdWjpZ81BskBrsifXwlGodmFw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 103456)
w66DKrHwqH0j3K5zy+iwVDwTdoWuyy6OlD8wh0i0a8SYB7Wbvqjm7C5bfTnjKoEO
RMA54yNLxh9IGFcckCVo/cBP5CC4eYPwuvxU1n0PF89BHJJYPmmwUlrjg+1pxj5E
IxjiBJjmlP0e5mMrNEme+rkV8L7C1uqDv8d5TJSzqriaalyLhusoMDVO9Q31uTp6
cKlomoM+FdK4aMxYhwY2UngPgdwS/s6Q0RPg20IYsPd4Tj2OshIu8nM8XFEphC8v
Xx9tqMXpae453OfigN7Bc6nBrST2EpbIDi+GGlDp7nUI+8WDy6voRLGovnTYIWXV
qSq3G6IzjKkUiRBMS7ssKJqp6OzL0dI2nim9aU/NXUQnZd2aw0gWak8KIWbrKFyU
ly3W9FVO4OIYkFOHeOUZPLaY3oj4a6vwLm9W6ta57RS2AYippabRuGZa7F/PhzHN
6qjxfhG/ksZsl6kKaD2jDaBKvUBdJbXwl2jvWZYVY8G6aP7NgOMWAdiXwx4q47by
eXKJ4B3ZAZ6DRFXnVk3GeAq/rmpbdXWUnM4Cys1N+YUmlqvD7QnU6uUkyx+RGNp7
HDrsg219jrOxxPQWbtCbqgEAm9a62/ntcmHS5ovpKrFa8FWF2F15DwU5sqN2QFRq
mV3fvqrxH8YAhVVVCCsANOEIrUlnJl2U/+846tQtIzVkpW0yxirhujBj4IykaHel
LKyKqJordw8LgYXL3ibqgglbEsH3+6zpzwwe632QMlKljJCa5iM2JcJSO9Y/PWgS
yP8EgDBsdgNzF9sEHJNc8YUuihDErnQM1WdT0uAas1YAv/ZoIVho4Hc+cRazpgyK
XdNGv3/4ruadKuWM1kuQGc8WovKDzmiwCIV1vT4Fd0Q7IM6GYvLInXdZ9pua0jgB
qvm/JWkgekgZszSIYCbYlYTDFMzZf5l4pYw+XycOqSU09jdgu9vHtlLH3Uv3u1nm
sHEE3WYw5TjCRK+9eJQMDGFt6VCnhUAzKqVFGyXll1HSJ7wEtAsRiy5cDzbBwSc3
vgwXtWHZe5ZhhaQBnfpxegvRYVb6u/3Tq9eiqMkPINK2P+DZcWEay3z2uJ/Npxxk
RtScFDsp/hs9DVKLLukyMWyDwXIwtiHL001LXsLMHQhfMkHlVsWIj+FOV8YEXAV6
JQ7t2uLmJJGP3426xOgka/J9fDimT8sNPY9jTm49UzpRMUAIp5sMhBgv2jCAQ6EA
UxDjsAoqes+Hd89eO/Mr51NhSjSRFB7eB8w4PsdFqBnS7CS5oj4rdzHRv7TJlJXP
jTax0x/0XXYyNTUDaAfC3XNzWkG+ggsMNmv7EVv6u61HN5XYxr1WmtizQ8aGCLai
fbMK41vp0vwoSp+dJjtKL9hoFD6HerTxCOv1adXE+RhztcwDM2mMygznHuVmxZEA
HRx9aHEcYilmyZrSApw8+tH1RDUsvZEv/FtXpONPhsYa2U4DCWTsqcHOdZug+xsa
pJ8NyPGmryTjuLXXlAkvnMNLaNi/o8RP99VWeYf14GshviqXfqLKCg/Lo0h755T6
85zSu0dmEg5IInizo7Nspy9IoXGG2S1l8FNlgxVYma2ku/oa/BDKTcxk5ag1Ij3x
/0QE+ttoPa+tqUH/axo0dW39bfKwiPHy5pcAXGxwuu3+oi70OiT0w5mt9Awwx/v4
3W6kCXEYGD5fdmhM8UnVD7DIf7m/NDekdI3C3bT7vx6vXwaHjph22ABEIWSn7Wh3
f6gPBsRJq20hDg2Ixb1h6MzqFOFOrtUWCPwtyjUuVNcFuhigX0zjdDVNYNmZccJL
biGgugOmkPY95N7DuGEf6SF/hj/skRuecw1X+d4z7G4kAFhS4Enj8eBvx34n5B6/
/08FAaTIOUyjlxZaGO/qV1DYa6FvLY/aZehHeBlScA4IwfUqJUmKwwN7ZwHXhpp5
bCBaIGy0U+/BKokmiAO8U4Pvvkq/YCeTMOmWlsQNX1Yj9rkSrBMziMIQdFS2CqZg
PcV/Ps+KeR4Fb01WQ92LcaEGh6qhIVPdf2yKBj52NPKt20yJIImUbRusC/J6xf+Q
nNxbeCg2SZlJUv2y2cMTCPcI5VlzukZVWjrio5GIiaNfB1LGXkvbb2yl4DC1FsOL
J+z0bOUKT0spcqkjQe+mMFCzwpQzsqX5hBt8HP5sKtqPXQSrjGYc4eqmtghs+nK8
hriQaL3CDHa5o2dxzJKiObywmB8egtTzuKZeR4/7Rl/Os7ykyXtUTCWWteqzN/wf
AA1B7yUdMWKp7hiXNqMGIyDGjcO1aANShIuSG3oUrCWqveDuH81cmvilMa1XNSjA
hiARpi+S+GJo/KHOXG4Rq9wO/Tgax+pf03eQ6XMWPvTQ5LlSEpo+RJBSjGwcp3pv
S6rdYO0VVKgkXCid2BibnWo59fMkgH1G4E9u8Hj9VCxe4Oumst3a5uE0VdhTWov2
jhduuQ2wfl4MMcbf3/zb30iqACEZmaJu+OQbT75wKVsrMjoPWf+SoUD4XgsPes/8
Ioyvp9PL/5RFeCrAy7tgRB8qwOUhGdh8N12qG+pLWE8oPLBdLN/fwRnheAYtlOAT
XWfG0lwgV7uEQTAbCDGN++PcNMrpoOVCXj/N6RRDH4Q/s9IA6SoCQ5NnJjwhNB/q
emuNlD2MLoxGgWKJMCEofTo0ZKUK53oSL9hYOqLecd7r7qYKJur7c7AllcBCN76D
tBgFqVc2vHOgD8j4t6rCISeprM23R2NUsEvdOBmkYV/f14qSHL3EUmFl3c4dxNaX
g9lK/dN5vKcZ5QCgwIBJkdz6qOwAG1xGEa15qfFg8EdC9gF0BeLD7UctiAnbH96R
46uoCeKBdBTFRiaL/sDSouEIUkZqFJn0L0YWmuwNbCks1ighK/mNBb/DhdIsqUKZ
2d1q63ShMQdooOs8616VNJ8/5yT30J40jSIMt8cIQJZANbYZ8FzWJP015DBXD5IA
EC50Pgf5FWWQp+MCZyud8y/umBAf02t21gS4o0AeCi/bnbf6jrsVoYVh20I2P0ZZ
NwNoKCWwfXliMwc0UnSNV2c7cn06LDw0jol5RIZ1Q+rJvxF0zVj/WGq9LVcXu8uH
gQtn8zXi4+Zscddeb97P9fkZ0kj1WwEj5stuUpzbx8b1Ju+HdF8ThM2jsyaPvRCz
/bOxulHcieQ8NT+F8La87IbPGK1hld04fjRDHdGU76IHLoF9BfEi+WwyaClZT0zE
6qqKp3EV4m4OllzDq5S+vM9LtC66V5NpCkfLwHd2JUpH4JjjvJC3w5i0zLjgNj9t
dkjV4Uwmovd7POLLTR4VQwpWDj7S5zY+Dchz0gLp6h7mD0J2A6jDo/o31rnn+nQD
o3fFzGMcyTYWdUYIAea5DmtE2fkQsntQndWgMqK3scVngUS1oqQpTwvEkK6Y1RST
W41zLbybn7r9W5VH8YpufislBzuvbH/kq761M617pQqKFfyaoyzHzrwxyvAFLcOD
BHHwGbumdSpyZfWBsxytvUw5QjWv5n3iqBB3fYVFlpGobxPvgV5A+Z1Ksq0Synx/
cHrIIL/bDe90cLoAQZ72/W3o3SJJ6+dWAmWl8114EExzDL5PvRG+YlcqJLU7se22
MUOuG7aTbZYIPZ0N8ib25Nri7ixjFCZWol3AFg8J6pF9o6oCqJOXbZGpVUpwqdRI
ku7Gpn8TsNgYczGoZXd0kvXd4XJ7ukeTj90VGEaCJ7l5t4+c0vv9vE+057hWAbZv
D2c8t+3CaXHNVQOPvKAagc3L6qnZyYMWy9LROH17ETEOhkyiSV06/1DM1BtTmZvK
VmQQ3rJAt5+hvwlGUGhKHtzJNtll56OlinUQStkwT96RnVsuEKH33lh+Q4morxWn
8vX3iI++QLCn1oCgwGyCqg0UD2YK98VaZwH3MFeVOxFXNzbu91M42F1LureE68un
wFxfZRENYzEz97Hvfn6KIRd6VDPoRU+xqNsMIiYI2LW5FIsz5kYfusn6TTnCTKh4
XaPBU5PGKo4E7UzLwWnfm78YYoxtvrookrn8M+ZmMcauMqW0ku2pBSJ1zSucbFDw
2U1g6jjgszzbPkN6tqXgi0THU0wYfjB/JMd773SCpv6e/xjjztQCRfQUJlnAzvYj
KH67CAv6DJwd6IevTa8Z4z5G5J+sy8kiDqBjx99qmhCeM1FaHD0ZhwpjcwL5T03m
dYmyof08R3dYM4thuD0/B0jjoO3lHt4j7RZADRlNxhgco2QUhwtdMWEXa2ElP4nK
z3iOvU8MiiXsKPnJWkduE0OSkobIC+qGPBs2d86ZzKJ2occN1BF/6TU6g+6l262P
PrC3Is7gqxIpr+AUskbYD+fuyKewZPxeLXTppEzNoFWtnMAyAMaNSknmta0DFKW8
4/ATZnroWgV78mnh3fMnTsi7QRg4+OVVjWGqtuQLSOUv7LCin9f3NOb0HY7cbpsB
wAJOWXD+dWnbKDVfxjgIGZHUt8DuxFpLlyqsz6USlK+g4wQ2Mqm9UeFYO8iq959d
HIWUD2a4XhVQbmZhGhZwBW3jEljuFBmwxdkRT+XWTIl/cZtzlBBaDnBBA1e4n2cR
DfoxrcTWz3vXhq+14WwZzAsIWF1U405cODZcc6gToSIgBiV8qqbTTwUneh1yDMY7
zdn2tZki60O1sautEc0jpEtYmQMB/+cndk5fjmQ4rmGCm2NELK5cFe4POOJ5x7mn
YpqvovWUFaQ6tqoWi27wtrs8fmotPXtE1Xtdy2Gqm1o5XFu6LsXj7/Tb/1jpKUvD
l8wLs8upONEXYd1jkl2RCdxQYVh5xxD7DRjbH95i6AZ/9V8IvJe/0fXvl4ZKfNn8
gwIszBp9R0tkNZ06kiqBJqHD+MfLSXadS3PnilqaoUcfeq93vMvvUTavQoticQA6
qdmG0jbbSI2xispG+8CuME1E4//R5hS3ziWzErFXuNudJqpIUsx6+e5xaWm1GrMV
6GeSmRQx/a7sYYaisT//9IxiFAfdWJTiCz4/zKIdP6201STrEtoZLHxmbxPtXquC
UiLMN3yo4TS2GUa3bP/OXjYkCb9DmqDAR12KeztYdn7ppSOEJ4MKHPCbJAiyfmPz
Ts/5BtaMVn3+jX07Men+5/M4pyMwHP888Lbgg23i/Z6YeKNktx9/YCTTZHNZcvWr
juFTDTr5SuXcV7vLiYNrL5Y+xoV4c1ibencB0GmnygEOTClcnRqQ4/xQcl2R0+XE
nMTyIH4inhBqCXU9niaJ/njA16vgMn7bMOYEDRYSbjXuXYc/GEBkFIZIfoylssz1
4g2l3fBJYvjM0hlhNiG0wac16EeiJXKyA1f/meoqaORKF5hyPOt+3zVQ2a/azsfQ
bKhRvxyBRICjh1Rry/+ctzEZohmHXIw/Tl0bBiCS28Wz506StyCT6jZkaS0liinT
4ncHwrjIhJgjxFflyBab0FvRkEwrugM+dzdcWYMfW9TYy03eJ4pjhyIZ7WqqBo5f
YIZFW1ASkovI928UYIfZBFQpcr0Gv2Gkp/OULkirtW3aW8zWpwG4kalJPNe6ZaoT
SqIu5OACrT+P0/Q8pY4YAX2H+8BokuGJ/oC5bTJXd2xZTCaEXUn80sOwBxcJeA3y
STd9bXBhLHqRgWXc4mc5Ybshqor4od9PoYKq6v63VdR/SpAZE2+WmeKxcxJtjJtg
NdqyAGl4yvkMJtHK5ISB8QDGhQuJENVuIE3ojrbM60MNstLEDUEBCI8/76EJJLth
sIbhfVk0gLrjZKXr1fRZZg0boCfTNqeRQlInYh+N+/QvbA9I5oRQB3WdpCAk7fBo
nh4YsDqYqwhfTtAuGhUZvzByta3djFMLIZo6R4Cz3K4RJt0Wtk9lrP2ScFmV21gV
CEqXlMsAe98+yydrkYb6TI4wTAE/XM2v1AbMY695/D/6oPQ7Zl5IIKPzCypiKFqQ
ZSe1Q/16/jSsSI0RApUUW/kAUWQi0vvUgu2jmUJyBz0c5yNAQSNJ91IopvTj/zZ7
3VMD7wnAraxkn+OkvQp0znEbhT2iihKI2XjYxUxslFpb9kMo3kHoEdvDN1cZ63lq
2fc7/N1IB7p6PInL7fda7LAU4jAl6SumMV+FhtCTW3x7ey3tbaefUnHk0nNLtVQh
QlnelzmKSSCoEms+FQlvMeBb/2HxmFRSlGLNxnWCRBXpI1oDdu7F6pjVKfwxVkGE
dFvMF+e7piS4WEn7WnYQu6Vq4Da/QFyxUMoGp1+USnENFoTknuv+RQeeUXl8FnO5
XfFmWNBjBqPx9rfj21c9YujngU35IvHr8pXHqd5Jc5RQrNiSsIqdjJfyTnztzyTS
c7geUzrvFERVUquPhxrnuGMalghsPFmt24FdwfxZ6SeRq87301MWgDAHg5OkEUy4
inzr7DPzFmR5C/kxDShSygj++529T/fkl4WT3ebMxnZdr+o03zvD4YSVdi7t5VHt
mmD/i5NXkzQ+RvKjGKyn3K8xvpj8ZTQs6j6cfuX/ysz/mFafgLzRB5Pfh3xKslcf
QXVXALP54fnIjK1q6LaHD4KYRhkrziafW2kRpKuwfZns4CM8JRymLFsZcTPHipag
p9TzcyiDrW9UiGmcdhrmwyg/EJPU+i/wcvKeUXxquUH9Sv9hpLycEZDt8ZpRnm14
cf43wwGRzi/rclnq6pfF0f4i4lxEgsX0JcRltdxLwT5pVOeMnQh2FAfeJ47Q3kXb
0Gp1Xo4RalVI7k0tvusxBNv7O3S+fCeTZcmnj92RaXl/XDlA7BSPaB4bcjgLEFYe
9Dq4nmqs5mGwMLM71R7VYyQeQgErv21YvWoGI9JNqXGhm9/r53iMApVnzL9LfVDe
1HCXi+d32TCduixDwZBoTjWOyGV7JQJEwDwXJz33QoNIaR9T44HUl/3s8acr32bh
pY1i4S6qknDyeKj+v1EkpUFpPEU39m2S5DldV8z8h7OEimbmEUhyqYhwn3CkjOTK
NRD9F9ruNbaVwHrOqQ56Nt1cdro+wTcLbPZaMbUTELR0idDbHMbzG9WIFTc86MYS
TSjL1x6zVL1rWqKGHTDirAdcIl21asILiU57wTcjkiJnh+rk7P9SvHeKNNK4H1wr
GxVJhyJww81mLvTrczPsduq9P6klci13TgLOw+OjecEnVc0dPBZPGggv+wKZqON+
8gSeaXJTxDY0HLzax3pW0pC2XOw573CIfXkRbElPT3gkauxgmNImrYMO7HFRiaih
/N22LeBRDiNNYJxGrIK9qc7eybJu213kLVdRLaz/eHI+tE8Ko6Az6Fz3fUp23zgy
EGB9/QKKOAoV7NMVo4WvCSsL6KIWMAlAMNw3pKSGu6DfelKHhmPVL5BA4hn4g07w
gwz7A835y6HpPgOfElkHfVn7g+YT2uGN6oHSo8WLf43//dLYtT3vOUTHFgmx8iOr
6uLaK+3OaWhg77f6oWDNrkCVdt3E0UPr8KuqdrE3a8eDAXPztO0ciI2sGipRH25t
GC6N8vsdO0WrNu182yslOSlRyc/ReFkS4Mj2q9YdgqwS01+gC08JOcEoBqwUEN3T
Nm9ht22Pa2HRQQEYR0sMhsfd9CrZV+5hbOq90Je2DmYuERWb/V1ca4M2IvvELgUg
jUChWyTLaNIn/m96a/hvKTGP2kE2wFUbX/QQJBajUQ2xL04ysA08Ah3sWafOklIV
mwy4geuIsd9edGV7k3yPd3rYPvm1AcmDu4UabvC5DGen7iDc+l3kx2i4VqaBnoRh
mu1PKeI2GYvNYqTLkLooJMLeFSjn0aaVS9KN/gwMtvmOODFFBc/y9oPN8OSL/OC+
SlWIYkkIIaGAdMPKOpwMl6MUXWbmqAqy6iAt5fuT+PDghUtZz9847cUWWpllklVu
L/EENF36zY2rPOx0cDsDEtESLQiP11eUT0dE2TMPhL2GIsfy5gH0mh4EcBN3LOlt
nfOC/ciQtiGobYsZHM1BoT53G+I1wjQnpmCoGm0AT2hekapsPjg3WCSglMzrdGqZ
83PH1dsfUf3uVC3iLvvJsP95LdkC03MnKfM4AET90ukYjD/dZv7x4/mAwgJ/XzJs
4uEvP9s7MlClOG9yCHG2Jcl/yK7nUh+XLdIk8tVYSmh2UTluUsL4TEP76dAnqCdT
oDa9exG/Dd7e3tfFu7Q6GApUc9y+6ybkYp1PAooEWWowgRZCWjyV49dubYiHlaDu
iaFl5F0Nid3z42/0sDZ3nMi/fkz/cJFT4rmZmrKHF8/K0ky+sRzME87CkKKzd50Y
LdZ9q+O9YNc5WNkYPnsc2wIZnZXsdIijyrDObt6TSOFTV5wl/xKHMrfDYRREfQMY
2QMW1UHoj6dkK5EbUIP/FvDnKivSdj0akPTeRSYx/nA8bs6v8OTgl0Q7mL/h2UZz
ubxpj8umR5t5rK8Ye4IpOizhiDQR5/phDf1dnIMZ3ceUHspTUfmC5PPrFQCUrvQP
SvkeJwZFIliu1jUlDhUSnxRnMk3kDdl2uDQ68xh2OiaxiSVlo5H3V2ahqfaijY8U
LwWbesSN9tSlsZOjOYGQDu5w3B8Fj8zGa7XOhPssXUIr74t3yDCOPUX2KbyzMTNw
H613NsWv9I3hi1EAAM8fqRhr2LHlL3JlBzldta5kDGNw9BNywdqWgIZ6RkK3DptM
atmEGmgPcHySbzrKte22/8JLX7B5sAc71P1WdhsP5/BL4Be0CzhBGuGO5FUR6iev
wpe8cXTtIBxZ+XQeFJ8UfwHhVUAwgog/9gvZPMVvzk9yepRUPWtvP98xiCFAs3gy
GKhlikdbN2bC1HA5svOngcu4vizERTIJc/DuT8GSHiaQD100nTqmx1ZU+y8veyqV
z5apRJGDPT8F5SFE3kmr+hPZgM19JCN0EeaHrDxQ0+rYeNfnh3APew78obBHBUTc
UTceQkZVS6CuEoQa/uVEzQ84gqNQ49hXtdtuoPkSsOzJ+feblC3VqyPDUE1uzl9Z
KcHyH8/OFskynE8gd29JaBK+/yDOFsI+eWFtVL0Q69LFUkJOQb9a0tOvY31GgAKg
Makl4mknwq3lk/rKi5naTA2yT8NJwvKtDZIUpL427QaMQ08VWxUCL+qS3nI+aUHO
ooTC+3Wqkd5Xh2flzKCmy3LUH3q2VlCoy8ESqy46Je24XHWQUCjk7VWwBlhoh6sf
BKekB3WMjpje/xPhre3+6bj3a0R6g9w7jbtzuBWI61T+WwXu/7SyNIX2oavRQNQg
h2VHCnbY+VWLDZUGb6MwO58ShG0vT3Nno3gqZdmZCCu5RSbybATwMeUyrufgi3aQ
S4nZqNW0cBEuDCZS0hz6W3LDEoyrX/jOXGhpAGGfKJRcsPyb7nPoRKtHso5sczJi
SoL87HqwRImQwfJ+EubXAUXIzLhYArYd0r14CvIzCBQuNZlqV5+dJpKlVwD26cxi
e2wpJ0nuglXijU0kMsFGRMjC46GeO8KICyP6SJulST1avhUSJYzhl9g/IED9u3qj
17fR53pGhG6aPiROFmGF8Cq2nyNyEdUUNuPoP/sDkxkV8Ex6NlzebOXAHxXYx0oc
V5uT+iuDouZsWvxTBD3h//VXBmghDhvW/QQAGi89BjvciV9K8tPP1cqgelJ1UCbA
2zY244CIbcU9/HtB1AOTzd4/ERa6riYSQdZ8oO24RvBXP38Y24gDHnsEb3SXgWja
kwgmzC0JkAISJjwuJJ3X4UntSfZ+NQIqtGreMiQeNYbzMHqb2+mhuhmMdKcLk+Zq
9u4hHlSYCkkfHdUW3GfzXQvIeb8wfnSc98HKaKUdReIz84z70GR5ekS8pguw9ipd
3QiysG7AgcSwl/oPYPEFyeac13TSpQQHDRLJwlIMmFLCIn76XiXgU+TXqzWPpKKD
d6FJYOsb52JrNbQnAQtmjFa+12g0ERrxOgZu/Vux/RVl//N36ifnKuIQjemsDUkq
GHafaVEJIqvXKPmJHxp+PdhmhtaVsn0xgevuJ6RJJgIla1Z8Qyj74V8F8zn4v17b
/FiLSc7GhRvZxpfk2jWqcyh3damY4i3xJC+wvoN8gvZw+72d//V6yNXcjWL58rEs
hEtzLTvDy0OY0GXg+Rdd+oziZSDeAZbWid4E6HP2xuXjSmVO0AKKhLKD7JWO1jLB
LJI4iKeRrHl1IF7+Gw5mihhv8gKJ0hWQCJCaS+7pmZZiWExj3horphUCrYwxR3gM
LbmQ8LIVZKfLZm+UnTl+RHoNIDJ/uN7KxZfapdqP71opw7oJEHx2qCw/Pkkz1yHS
cRd/FXLaJeNK8HGqWbH+Jr84qpgZe9h0K9RZNsZD5tU0gzOWRfBFu/DcylPS7tEV
l8C6DY69XDRo1+AEuj3GannJzxfIs/ykkFpszZpyxJXLavGtKQfpuaf6OwASikDU
s5v4dMqVGSEUxkSTTQkDclk75avp9lyv8kJx0JPSOCcSDUwvsCRnLzSK8gwZ7NlL
VXywOqX3og4jQi3CwjfibPTwBHzqIfXro7Irxh/Pwm8+jEBUfKXe+Yq0Wk+SFrb0
E3Bjj2kOEMglMebr9M6H9PzjrvmcqU5UoW7Vuptd/MdGS+RQqi0n0aWU0JT8RVr4
zzqZflAV3SYLZDpHVSgHQlHEQEpdd5lAGlQoFMaASrXtzYhUDLODkR2UGRUmOekp
7Zy4QUJtmS2oV479iKmzBfxF7F52AtTyV9cN6/GUnvbZ3XEE1t8/t7yeWdDNcMbY
D/DOKt6H7jA7dfOKhlmf2A05kYFsFezlEG7+fnAZBEA4hROndTELn2i9Mrp/aRsR
Y+m/9+FllIol3fvjbrj6ssfNhMS5xHk41UvR1FTRhnEIXevH3myayP2qob/wBVDR
BIcmlEErNVqdtj8Kzw7xjw/Wli4w9LRO3IeU5FMePbf/mfE2f5rMo4KNbkmPLM7t
41/o2Y8EX+kF9PFFD4CJ9i6hzz6jJFoEfTeSfGbvgp0SrwuCn31FraGvOzVyrGMh
owyqMcjMRTek1ADtksG6wLF3XUXzeUaPMc1xBF1a9htNhsMl7waiGhZh8PYLhpFY
vggARWYLEGGUWFfqkU/Ftpdc1+xSxhUgYq/bIoFpFwLyjccs3Sjlm3moCmuHQggp
fJXAU+F1v6oHOMa+SnN8khMKHbhgfp3zO9pFNoGLhO/S8uqZy7Mcoq2HXo2pwPN0
eEOng4WoEMnS/GT8lYVtY6ZaOOB0ZMTquwHYCc5PGcK9qwjY7LYVdXEoZ00jJz4o
WdaWJcV3E3Vbnt/xsVwrSNZL2gwBw4/gxIbNGdcj6xbqjQ6S37vnz5S3BJO8z6xO
jEYEZNH126XXZGbH/dhoRd6uqfKsrDYnhdQdH324UxVf2WClokdMNpF5QcUtq/SN
OMEFlzh6bQokpFm1EiXO4k59LIA0iEXfXyUDu/+jcWNYmAzhVf2vPa2P0N/vAXNB
UQdMSU6jjimlSc62w/gWtbNrT9hQeQKEYddhWI/NanHJnMcgT/CrOZ7RSJ6gO1kZ
/Bllck5K0AIe2QfgJPj1T3fYm+d/Cli3A/pRfZ2ZKDw2fJr6UsN1YzMi54tp/poW
shaA6711i83SWmzT/iOKSd+m553F4gpE4iw0I9l0Lr1CtQse8/Pr8+WLcS+vQ5dD
HIq5fOyN4Ltv3ulRfOBz4AoMpHbEHoBUTlLbL0dbiV824tcBlYuzXI1ted2hRQHH
puV+FwLZ31hnzJFIlZdiSWSkuiuRguBC8UnlgG1ZDaK4ZCsBKh3DGLcAULahN9t+
MvPNFZCGQCtdOVhyNKiZFxDgFalx/vEJeTrbbSfdIHDJ5Lk5v6ZYkkWeHBTxoTe4
0eJmxqvQwO/MmQ5uZ+feG8prBQepRv7Qm70KMHUNmAjadqygKDQS5kCD7tEaV+7v
EoxWOGVvF5e+DiiVK/NCnkb5CSBNrwjauzFJLVwBfXoXziItCfOVwP1Q2IjctmSo
wvQetT23Bpa6JwiUB6RRYRIBqY2Y7pBYTt5Ldx7OHv+4rUxQe6rEQU316CuKOQ99
iKzneIXU+M93MYj8svaTJb29dwazDoZ4Xpc4DQUk0o+jVsrhq1UhpoMc2LJZaUwy
3DuK8IJHSRkbidDgX+HR0oG/nK4xBVkDN3fy4WPLRSPap5CncAqNN0BLJBESyuVU
R/KuhK3emk0KkJLoyIH8tSRcslCHs92fSSRYLqYmwnnhaf+OMiwxc4WJ8SNetVMF
FVcnMJ2gCaBzC/l1/bXkHiOKfn913QcOoGqoXDyfEXnBUj3AJD3uOB2nRNTVA0yp
FId2AoszXuFq6YvEdcSMoiGgNRavRN4oU4D6HALbOmB7qgoAgXW0MFiCgZF5sXuJ
WeFDBiriZJi1szWmMCZjirKxvgxCJ7XmsL4+h4J0NNOiHNoQS4LQsjmS/k6CsLs3
EGluX451DTbTuJKaHPSVJbFHjQc2Ri+s/Y6Ai2BaGqxqcZVC+78sAc5n46jV9Vc5
NXb+ggdj3l8LV+58jwbZQ0t58cr9wGCdIQgapqvHUwi2z4hbt2FVXPzEIl2Pi0xH
gtMbcCJwMrqkz5hgeTxW5uOsO1Pet7j2QXqzJ9+bR9ZtjaRHTkm3JOfINZyWcqV6
b1TM8bpm1X6KDZ+BfZsqZ1S3QQ4/3uyTvP6Eg/GnOcvLD8fOG/wzpe2iguw7seuz
uqKT/cMqEgJXYygSE+gE9qDp88Oek9DJ8bTIZ+XJQUELRhuMlsAkPnDyFddtKfI2
Y9FJMWl1SuT3wkxW72QZpmJnsG9d6V42B20+/ODWGpag+LpQpWsB5b1Qr4z0jRtX
XuIotQIEo9Sn/FcGfbT3+oIVFRuHfBVAr1+qiF/tsWKrCQ1cdCw0E0fZ8TVYMq0e
OyiNkYtcG5ALllRzsvs8wrSe52NoVAQekYB2CSRlaJeRwqRqydTTbgD2u3APaTzz
Y7Tz9CcCOrds7oFJEYXaWiww+LcGecz7mPB1gsMK+TnqWrwaKBSqQ1YUN5JsuItB
cRVk0vLbGOtKXUk0Hgk1kEz1x9tSul6+mT2rggxFoZENr7FwgX6qQfSbycSaV8Co
U0zs3gjYGaA57kCID0Ihy9UZvoWvprEQoLd4GeKEOIg92j8FqAaoQflu04E72rSm
+/6cEG1CBJ+3iHFwcuvZWanCCLEEKbOGFgWep3vOsjhVMDJWHhXSjlTonZHoOdkh
6Xcv0AzUPrbYCZ9Pw+yi2S5WIavaLKAoWwynOpfYL+MBUJ/3ufJKUNEXmUgSNPRn
snxTi66ADLDG894bIwFMB07EdqdqtN349pm+KM5vhaHjem60wn3O3nTE1RikNfHc
WJEKBiG+l8/6dbQIK8s653AEZQxnSaswtsxYq1Kimw1V+6ZkTVKgqRPZ/orIM8Pt
hvkguTOVBE85r7bqMlyGzCqLWSMFBXrl/KYYuBH3m/dQrtzfscau0aDL6QNqYe4I
TSiufTajbvQ0+bBUVMhrN561udpZco5ucxV5sRufLcm2ercJDxFTZb6HWRhFHMUm
4HIa2mPYxdkxgde1IYh7oBL8pJ//7P6IRbj8gQy4gY35bnCkWzoDD/tgKehcChKm
FaolRyZpyL6ruHIO2eV4kKeLmSpStVoHHAcDIlTpz3/UhUX6r+Eq/wS/d5Wlt3mw
9oCcHFEdvQCU6s92pSSVevKUuzE0YEwj1xJxW5o4pHMyuviqzxic1GShaRTE/zLO
Yelg8Oq59m+XkS3+1f7ed38LuTACtAP5rVDlgTancRrSChnwylATETnMVSfDF01+
0u9EO/Sm4mmdILTAXDdM8h0ORj6h2IEfNdAisiAmVoUXcJYVeFcp9vgIAw+aNX76
LlWNQMFPFrhOubPZNGQWi4+TbCQFku8NBaayGDHoDXFKX+JwCmJbOa4sa5NfqWC/
Su/Fm+xcuuiIsX40tnAo2wNkMPCzSdIJy4pbmpor6+PKIxICde25lIlnJbxKvKQf
cBKO1xrmn2FIKxS8upoc5eFAk/GWXHMsJSrKazztikG6YTgZ5llGooplw8NCrAUL
cgBe73pXbw6uOSy3Kf2ERnVKoIhJsIeiwyLj7gFRaAcN2PI8BzTP1RkoQ1w/AItn
g/nSnOhGDmSq9KZIl0edzfC7hUriZnjbw79n/VyBAWmqKL6nrTzu4iKv8tINjVsw
VAGD7gw2PNj6YSC/Ux6MuiZct43rrG8lUourLqXH4n4AUEqYpPrA4Kk+GmGBEaZ7
V/Dc8BMU4BoWJ8p1ZS6SSTDMbcbXxzCcoEIIMvCgA21nMe3VWrivxijX1wknh61+
uee462PJ4MsM6B/gbYYWjnsMa1n/3mnqYaUrXAKIaxYhnojwz3CVRP9t8RtsJCUb
TF9CeTNYUPVddOAuIEdPgV1sTNwIQbanxROcQSulYskjzOvYtiWMXPrvuQOZ3BkU
bgXqzqrwAfN1aZqVqsxHBjqoeXnoAF2mRU8BSqmwuKeF6dXPIybG8JEz7ofzXy3A
xlUEj8zbeQQ8PQ8EZONe8hBRg2c83ijutUUgp4Rh2B3DAshY8C4c7hHUlzz/gcXU
cc1T+lOLkBFwU+m9kfq8LSp8TDtKZv3+i1d/w+/MQuqGkenUVFpETB5oLaIk0XMS
zZwLCDIbvVwOKySz7s2FhbuDKV9MS4Ytum5UVETMrRk6o3/4fOScrTSv/ZFkYMBe
7CdaNC57DSKvz1xVxahsIXw8LU04f054rmjKw+IRHeHLFTgf2pGTx4Futo76rS6P
ZVSieh0PsVWLdGPTHsg6yAwhGgCaKEmRdS+Dx4muoKJcCrvw13NGpMSAh91aMLj0
ayazsy+FiBiGEQlm88dTLDTnDOkg9wadZyKsgJffpFnhSTpRNwdoOfbJ1+Q6IJvB
Mu2MiRRfawebNeidcBK4I8g7WkLBpcEjny01ISwmpHN3+E1N60iZSTCXRyoKXkEf
tohU52AeYTOduGA7mgN4xKC++q0N2TJY1MOf8zwnRX9BnekKjlFd8vLg4VdwJ24K
4QOqbji2eTxgHxkIrRIrlNFbV3zkdfg2lKtfVMqcSETm9H5PO/f9+WVEnK0cnu5W
38JmRqD7KOgdUukCEm28r6GOp1hvKKKyIz1IyGSnJIG+SeiB73PiH0PaxosnWtY3
E9FHZ+d64En9Cx1rBnumcMhiilao1bdWcE6ofGsTA4oRirjFukkt+laR6hASunnz
hOt4YDUGKxlbzMauIs2PzDjUEy6lDMCZSdEMkI4Iak0sMHOADSQAEw8bWTEJ6275
jd3H6Ybbh6kLzOmXjY7EgeriWPBX9yFkO3Rx7/unMs9o8Mr6t9mS4k5/AoaIA0Rd
ut/ovcsthkAFk1TARcbOnRxTy3CrJsEcMrdto2FbPzKSHXy6VGtj/V/BJCYl9f/B
pba7tS2G9oKNeok1Uls8/mlLt/XX9XUD/eHBE0OO75mBqcgZgiANeLBXbfBQFnip
nQSC0Xf9Sw28VTl2aqlrQFRtkRdHQxcS6IhYO3jhtM/FhuEt/5zy3/mZkYg/nvAn
/e9F6g++nL+7pOgcVkAyOGd/IAhY/ptVTmgIHY4O+L6Z7R3DHj6QVB8NDpm/nw/v
C107jgg16LAdTEpTvf+kkjmyiWR58NXlZUJxIo6wvsQ2iTWzalT+QWKDzbw1wQN7
TDRcjn4fwH7xHQIy4yeVwjXtcuMhmvvWM2QZPlDDz1tye9Li/C0VeGgkBfJdkNIb
7G06qSLkI5mYfNNNO/zo7gk8W1PW6QJJ7lygmYh6qhxVd58x3qrXaQGUIgevKHen
GoGcMX49IXfHEYfChViFgSqG3vz3HKU/lpESO+Wq1ZFekppg+2pL9dKPKBK3TCqz
yij1TP2I46XE7luvci2UD6R1Eh4ybeKprmpLZs3jlffWvgXSub1jAN7eFiTUs5f4
YLQwIKscaObUsNx0zPj/D1b2vEWo3spW26fpIIgTBHPzgm+JP88r/4+I7nSQuL42
ewOrfzAlhQ1oKfwwTIf5AgVLymeYSHXD/4F2h0rzb4uFdJk8F8WcQqFqeldqPWNQ
IQ6LWPHN7XtZQrxIloMaHw2rhxiR2YbtPfKV52VO2xd2xfGI61b5jrI6smyhuKyf
qg+QtRcrdBniYpOmcArKUxrOctyKO/CcI18rXJcCKYJY58fGSB8qrWkvMsHt0HrL
6GgVqItGr4IQeFjAczCvoJ8iEbOS0XfpuygFVNCVOO+MGeq3g3KBCqK6ZFO8KHsp
aDXB1X+zJp2ShKA9t3gYfxNUFhsoLKUxZ2HDF9aaBswYirzGljpjt9sXl+KysOka
1uFyU3RFUhs2Mk6phtwasvnSaz+T+FNPX+yeb+EE5dw3YK6eErJKaWaMtahNXtpl
OGPjxv/XR8n+ldwGxnMylKznCbFlTFPF3nRGsP/h/6RMqtJEhnV/MjQ9/fDSi4ST
Sg9/IwO/y2jnDqxKcP+aa9YlSAWxTdl7SO/UQ3l9fKBK8a83MdNGdYr57tBCXC4J
DZ72cQ2JU+z4G7JkqvbBumuXQwr4yHoWcKMh3xKBJf1kLnznKISjbyjTKCwpeIge
+D29YmLWhnnBAYDDSHgQGupHmRshRCUgSFFJWYo8aqL0mc1/Z4mKT5CHQgbc9j8Q
WKglRMLAidCk0SEKXwNvSz9Wz88ua8mjlEi8XyUYIhXPbZryJNaEEypGtcK8rsjY
s6jUJXlc/CYUeuEPcBY6ruEpFALn1zJosvyFGKN0FqwBQmuKkifis9dcYFtZZ6EC
55PwZimbATEr4PIyZpz2rXoNpafSRS1/IEw9o7gmYARcGckJB3Jn0yZQJgkzflRo
q1dwV+PwYX28dfbSn9Ww9dAH6f4IvFUCgp/DAPHvOF1a7PAm+wf7bBKJfDnvcG/z
l6wjMkfWyt/+kcAs8MzUarpsPCWsxl94YkLi6vnOiE8kN6cPCCZAkc1uqFrWivGH
NsnzshoymWXJLcn9m28+5YC5KUT1GvLtmuhvrf/6yzDNUsnW7DcYu4XQLZ2U02oU
9K1qftlsgrmvnTebUpArcOyOHlVWOgEfnnQCkmt3PgmONSDepLtSFWtdhyFyAl9t
ffEjgSM9uU/DX7KmaUVW22hN2IupdqApStPw7yWhqDJADyfx0hQkERexssdGe3lY
lU0VeS/xuPXRFhh/fee4GBQzigblbSLDGZwKOKFLOL2JjXvlQ/eKq3tpZkzMPeO3
qXX4tqeA8VPPvAU5oiZZTB3N3XcElhPW2cvUPueoqOlwQQOVvopUK/aacJuEnFCG
h5Y0DCIp8gWsxzTRnEs+g3026BT+3n5SmX5tsW1ECZscZl2u4rQD9w1nhgSaiGuz
aOIjcIhPZMY/KXzx5ZzSWOVzgvrI7XHjmWMBWEVh+rsyqEjDRrTBruzsC5hg6S7v
EqTy7CzJ1NUvFlJsKM6UwxOECxY2wmSviXL2Ej0UTQY889gZHNunhf7t1bC77NrH
pnlD0t0OjaQDxUZNKJKjblN9tCpvPBOk54lY1zzpuIxOxa+1qUxGFHA5mwpjG+gF
o5NZF3zNbXpdpx53RYCNQrf3Y6FHCsW+B0kVOyVFj1UTZBXt+BaSltGJCyPPAvvB
gzjtWYZKy87vhUpHl2HLmYXU9rO9hulWV7q0bVIPFgbVH1ShEs14ddHuWufeGdcR
rTzHcuoySK2d7KpIXBZ2KAO5h+xrgS6j4xPCkjwTb6yJloOmKTfrwWp3x9Y7M96t
5fsN4A4Y9TLHBLdN0DWIpmSNDY17CFr9o4zVbeo3voAcsa9xkFEDe0c3jwowbd+2
Yjs22GLWom4Z7FtjI9UdkwfnvNS9Pgc+DakazarfEDAQ9IwOA4GFhmg0vj2Fz5G7
bfCLbAzl1lu0GH9MAzh/p6wPDwIuf+iqYSlNb1uvi97ciZTnUrjB6rWkv78BiIdL
aQnjqrLzSByqyYLJ79IKvH/1x9cWulXlGfK357At+o7BJJRmSTen1Nnrwj0tSonu
ScCINrs0YMYo1f/vJ8fkpDQm95obvqXs+QDbdFzkuR4QN4TJ/vgFsJQ/E4v9juYJ
RSmZAc70x7CF3raIR/hc+qzy7T84gYNnjnieUmoebS7YUV/vG39M034Zddrdh0aN
y9VepIq8eCo2sExJcLhaUiZeLoVTiI6ljCiGQcb98QGG7aL2P9vVvWRSo2/GZJIm
8L8ef+iWm8ejE6gZnPdmKPPPj7Kqe/bQcUzYqxQgj7A43pheF1PzC9gJ+U9mWwgI
BoATLUmGnUNBZGOijgHhAHu9NYGgFbLPsCvuxtJbGO2TME7xwCx5zZdfH7Mksg5T
TV0+WJ6Fc5lnjSLADYiHo0Cd+r3MApPLQChbPlG2PeyGe9BYZbwAMPcnhBi9qoTc
dBeAGXdBbNvh3jlm9xA1VyY9rbHkUL3euCtLsfcAGLP9D9opOuvxOcCq5p8KjktZ
5+HjfSHSKzptoGodEm2GXIGgbLRLnd297Fjw+MtyIm9e5ID3B2RdfXnAAzF0PRnl
UHoxU/F5z5VEYtZbJxumwrChTvwSiNAcdfIoHFTNEV23XU4WJS0WrHbqWIIb9VRG
JDZ4kcRmlp3Tngbj43Y30m8IdHgIlriboDxHRcdprAOVnxtoumugeJI+bI5qpIdn
7PUv3RVTA40c87bVdxBBzUUO3Hxq3THuOQtdOlFiLOwXlswE0tZGs1uoRMnlcu8H
7Xs//1vI+adOB5oTSsz3YIotdWn+LQfVfwyed64JmmYvfjGEzoTrio0x59nHrVX7
R3l/g3sGoeOeELh5ncHUwrpeIsDJy07Zm7Va40f6qVG2U5L1pi97benhLCTlhLCD
c6dr1DhAjPPwbTjCdy5NiG0oARCWW/24uK295zamb2Odye9BSy2g0tRzMg6hrycL
K0GJQ0BwYaRA2X5qGVPrTrJYPgP1XnloPrHIESBUU3A3/UJiw5d/dLnFV2+pMGF3
LpTC839n1UiFWf4/AFnCgA1SVnNK9/kXE/aMzq/SPr8jxpFlISXRoTbAZd7rzzFn
l6rLcw+cjcC1Me6oQJAFCWGn9j7LTEbCkoPREcN30FBrSC2HqYk4nxDVEiPojSAA
voGo9FlAc5eCqzK3VTlk8pForGtYWi84u1Hmfa+/zmXt3RkskL7jCHS6VpbeqLsk
nY0lnERaUGV8vb/RQ3svFdPxIu7opzQ+1OXXX7RZliGcGGc9n/OHwHlhpIgSj/y8
UAiuAqpDeUfxwYEoNprw9xwUfceiDzacWxfewr5fz/VlllWCaZqVYUktMunVtSrI
AMSRkNTUrisFfDoOsd6Wdq1G6wNB9yhkj0GPjWrZKi1RnsdYu3oCc1xY6H0/Vixe
tM0nouYzwRYldwPRtlKzNteofTomjOjdlnjGWwaKFb30hjHzq8MduGBbBeX/W84y
u6z5U58Fvad9zGXFVRRMwG5RzXPsgQ8ka4LM/jZwUW2pJavPTqYu9EJzJI7SabAt
8a38xZKGa7niTV2OJfPOkNQXSBuJO2w6nlZgRZipZoFHGzmonoADY4HBAK0Ci5Xw
7/HqvLlQhENgjtycSEQCZLdu4Jyz6ZSRHgVO3ySzBRy4B5XjqG8/bFmr/gfVvrcH
pXAzYQrJux397XHYvbmAO/tIf0yzotRbtDMUe7yJ54h8/suztJ3hgrnmYEH0Xtk7
cccARbyUmjz4/usZyK3s2KQKzIAanMKqmiBHRmdPGJAQNKHz2BlBvIM8Neci46r8
aUeohFtlYUJfyrqToeKDWE/RhV63cu6vdnj2UQPKXNspogZbD2o0CRNk1/UJhYM9
zxxHckm1xHIMJfM1s6ztdFc40hs04rbZwWbSChxnmfNimU/YT1WQtlblDaIMBGV/
oYCn2femSFpX9lhPnKI+/HkGZXEQTiU4WXtKK4/kvzfaIqW3pTgc966v+Hw4cJH7
PCKpGsbhsCZbujXEjk5D5qdLVaxHnsK6ByGm5fCedCvQXFMFf71HaIhGemjvX8Vy
QQ4QMYJYbrpzMSdDdElk/Tky2Q8217AGzg0Jiq0QMACurflE+DjjPvPKxe2EurN+
Iz4WVhDeumFRGmQc4n38G+Aps0MOSzc6qsxBH2nLxFbwQtwRxPXgATqcO/+Wxi2x
fYYWTHgzBIDq8IZBpapKF62BcDiILEjDNu743t8AR3VepPx2XAuX+O5LJccrOgvu
RI4nCiNb7q5GW/x2Hm7r+GqozvrYjxiekTIYIq+cKWTxZRQVlosy8Ben6V3Tkna4
QJ8B7msM0GkSPaezJZmWSKVMw/ZINGFKfaJOeInNhB6XXHMSz8Vvq+1z+Acs00Pd
YsQ6wzkiL093xiOnf6p2eU8XMYcH7MoF7rnPS6UaYet69n4NUnwbRK+3CXVJQWVH
SbU3uFEDFFIxVd1vw4rIdVWC+pDU6KPSdqP4HeLJDzDOIy084RhEIE5GQBkcCqK0
IC/p+8lG45Jep+tKFy3xxZEU4fuVoG59Ur7OeHGIIts/WWcDZDC4F7H7kd1R6pfW
YXCGTZ/KED/JoIhojZLkt9IadYE/MxNvC/QxunKg1ZgQIKw/6qtdypWVIaiwkWEu
Oszc/yyJudGxNClcxtWclt9H3zJjCWCy5utKH97I4TiE0QotBGSFb2hecTpALtqF
nsfZatWLMgmQ75mZudGeYmEsS32DVVSOa1/gapQsRbLKPpkuQeJ6dfX4ooVcDthB
izny2kAPHciJv0krLclCK5g/bIbe8d0ouyO34M3KvthWOqJbgWVEDk4n8p9rtF2X
61LsQDaJHfujSWLXCtAbPKywQjeudaDMb9OdpBe7unv5L1M5zn2TQftpRJ03PBw1
GwMN4BKLV7ZB4RyfwInmXusHofslrh5FJwMfKd3Tpko2VHHsSgrGFQ5lZrA+9iEN
x99fN4pNINcDGsTtQUOQarSW63WSKw8JwPR9dLZHhvNc1+FJ3qD6Pb9G97GXSSxm
SXy6XGmrHlUdlWEMuQalAHu4+8oljDS0tlOPh6BpAr5MiDN2b92oLS4aUeYYHxIT
lMdL7G2uvswoBtPyG0AcAW7ZWlc/4DUGR4G2QK0DUo6NIxSkya5QfW7Jd4dDe0Sk
mgZuGKNxLhlppYpzkKKwryASXZbCJTMk4nr/NIVRmY5pYHNRxghcLLFzu+5Tr4ze
4RQcvXwtc4gM2wPB5M6upHlzcgxBJ7VtNwus1qmHEHSmIaFM33TwQzZ0yj4Mopmc
XpL2GxORvIC7LBvD2Bmi1QqIx4CnmsHYTNfMOQs55PtbI9CeBzC/nAq7DWL2PG5H
DVaV0CqUDXg/st+MzDl1btj8r3iHiY7GvrMFzt4l2IRubJfumhI1En4vt3P8FP0s
Hgicd3/V82fUV0048eb2aDOi32p5yHAdA6OkWcSCbHIPvxzZ14unZg+b3hw+IvDG
ojns2FRnb5yqREA/3olqaQBVU5FjEOhb5YKWiJqkl6xOXamzOix6beZ0QW/hsxhp
igNdC42Ek10zt8m7D1IldzjRcRqDJdEl0pcD7qJ6j1h1D4Yw6U/prfGP9SL9NW1e
AsxlnIm8njCRtyb6hsOKIIuSTrjX3VSpQKiFd6/6Wiiejh4UrmgWX1AwXaK1N+62
fxqbwSAdQCXmzbO2pkOKVKY9HBg8TCcql2YMTOXUQEVMDaeEo6tCiwn4MK0A+Cpu
25Yke04YKzdVQh+7Y5Nua1dml/l5l2aMcIr1rWqWsMyYzOsFyCyvH8L1uAWjxvRG
6ZhD/cQrtBeJlYlxe7CKepvBZeOumRMLi1ru8gsFg2jBZ7zTl/ALh0lycRMZID2I
wuckMAHSoe5xe2s7C/IV6gWB2/nWm+EebTdiJ3K7z4S3BEPMly94hIAGZSuK1etu
15KKdDqcGPgrhX2zY2JvM7F6CbubI4+oneoY6WoR9iXKmz206KS7Rsa6HEEDsACP
w8+p5xbnzghsKLYm684bGl7ZzMIWZvYE1bYGsxu9YVIBl1E5wMhclRRt0Rye1koj
ufFh3ca3NxCpi8aIi4MO0Kiu3slbAfCM6S11GtCccAMX6DC0IDBYQkcu0/raldjy
aPDvvduA+iWFg4SWTqaVg6TlSC5VMyK0fGwOK4PIZDQfbV4YaQH5tp7uA5+5v4bH
cluCnuPz1kRBucAHz9/ATm+Up8xdU5lqYPiRhujvhhRv8iIAeSjPhkoMyzGuLyp+
zAkq1ijTqgGIoII3Ze0//w/3t4lqJ06GQQtOgOCg5ZlXdDE2WjadMfzZ0rDDJ84J
BfTn9m6oKL6Vv1pJJPZ7eo6N3gGMcZ4PVSSNd7Nix/+iszOnVA0gPHUomU1a+/Fg
2klVWVNfkR5dyN0ALf2blCUC+GUGf2MIdqnpcIvcP4WFq5WDgUrk4TV8Q4XA4Tfd
x5v7d37D7RDxtRRcvsLkbsGcpuri9LvT/jRqYeK84lDl+t7v0qrp55g4LDwmef5I
KcX9GacRgocqkWDBJCGH82MCGHUE5x9WwpcmX5Mj4ASWuQgDGshl/ayhz1kUdvnZ
BXT7yut5oeARDG+J24JzPvBCUHHtRmJoLdIU0FQvRdtWIerQG2NK0pUS6dwCY6mt
nBAhRRMnv8ujsP3uLPusDwL2g6NSaiN+88MbJupTSltsJQvqm+b8mSyYvgDLYeB0
uYBOqhYFIjRrashejEtObufg2Uax7i1Dj+VSqMYmCsxjgS2oS1MYtjV8FfvAzZen
aEiL0z8hzUT9wwD2GEfi3WHioveAKFjlWig+UHIudFfE+47/AyujlzgiNNBIgBRM
lLE+hyHLKhjN1ZCJL2PlEuQAzpFCMnxeXGSLxiXrHOOD8hkOXXBpfep2S+cUvszn
dW3BtpbqSKChvwUycbbzdvIF+3glAHmnizaByAjzBMzNy92lBWX/p9ZCQUzIHjFT
iSQLeF6uLpBdG/nslWLHGJgXLEZL9BzrwUx+WFYi5FeiFreFSvXjLg4SneFvMClO
febdiYfN8wMwZUVnmNBUF0cUiaGY0/YDLiLE5A/QmNau4NLsNBeu1xv1lBSCdd9v
EvpL7psOsDmTZdwZwvZTqaMlbGN9nLECXJc6qza6NxNIdOU1i33wn+Gt9l4n1usm
uzcOteQ6O0+6f8MTL4ws8BDioUVIMTVLJWN6kM/pvImS7KfZofyorWI9GElSfLxY
CooNs/TZKiCModmg+An+j9WCeIe0OgV3XWK5jrdoqYcsViOHwCJ054ISEMauk+Rc
m2wmomtjFALuGZlhdYyRyG5/hjzcRG/HQfZkPj1vfaWaVu2yyVtukXv6Ifhfc+yI
+ZAI+QqrCpC2oT16o9Ur6mXJeEwwsqoL/AchGzvzc2z2LuxiDr4OPDSlsekchQ2j
8vERwpyx0hKXzTqUFRoFKEgbsHeyBAXjXs8+OT2T/IJ4vmf0os/i2Wq8WUkuysXc
ZdW2VwGBFa2OHn3ptJpTSxhVPjgGr5SMMGYTz3okvb/tVdwHivGhMgb3k4igZuLo
eVvd2z6HhkPPZAnVUTlF3L2rtrJw5muf+ofcXZr9me/9CfLclKuDReeiGKkWZWzb
ZtiTCYjxanrvYdDPAhexa+o3QiekJepmV0SSTLKCL91hK28o6RRVHgegTysX2/lv
Pru6O4Mtzhp2DCU5SB24SC94wuFZ2BieLurqZlISiPl+u5sLPEkrBhPkvH7gPQHK
hUnMHzKm37OiERR2wG7rp/E9z1DMGGtAOYhYoru5VWZB9EUH7kCe/E3mh+UXf46S
VnWvnd8I/b7X//jgNi8ayY4MJpK8FbDtQcuX0EZrevpG4MTbWYnVVmFn8AZ40imB
g2Mui+xUeQtNDB+qeFd2NC1T7t3PBfm1f5McbZompLR8CkI6e+FpweUy73qxuKxy
4OfVN9+2CFmsHMIgfFRIk/gk6FawCJ0Xix7X4Dfo2327+tyrFnWisFpJhbWLzDtT
/oMiPiAF5yjOYiBZPZlGPv2w4/3y/GIHD924Oc2Mm+QgrJyRjIRoWE5rboMoL3LV
2ITgj9b/HLNQjvuc6gBM+E4uWUBZFiat403A9VITDuVaNalIyvoNdUCt2ntXvkE3
BkKlSc/ee1R3FLwwDvjZaWmpcziCk6RW9F08eFafY7HrpyftpQblA7Gp1j6SYreP
NwR7TaU9p8cG4L1iU4l6coy8NaoTSZny46rqalH2SXfioBZ9saoAwVksj2EbfbK7
Nqa5Ctw7MQN7IE1oCR0Wg1Twd6qJNXxWIw6wiLFOwvqUmiL21zgkEyqkAsEUP1v+
Akl1boJgVr1I1vHROEuM06kWxlGiekbcak6R1rAofT05BqEzJNBoSjunrn+eXHam
NkgKC12MGk6YbQ04GsD1fjxYSyuvZG/Rtm2HBkDBrb3MzpVZ/jJVKSdkzlqVBJfH
gO3zoiCEugauUJHw3cLXirI+pKtgp0J5it8V1qlSm+UnB6x2kF229CJze8ITu6XN
o1w9mpu8PDIQFyMktwPC64UJDsu31vrdWGsz9yvctya8ZZv474PK3fJ4T5BJ+4JU
qd6KZQ0sS9eAAau/mvha77TnmyTDxH9MlGnVsM9cXYjZDDmv32FoUMuYxzhacxKN
0h8Dbmzsb9RGbTcppGvg8Zo83aogjec+Ng+Yu50rsqgO/S9lxKbiBAPWRaL7yYlQ
19mdL43a7/NbWDi0L+i3qQ4QaLatlHDw4gnVqLJLDLweHrDiYTST5Ijc7OgKFPqs
Qk8jqs8FgPaaCi5ikaI0JgviKukQpwtB3uIbHmvX7Lpv87jep3b+IE5PDmATgdC5
27AJ2h53rMkm8uTGOKtFR/BTdSm7GCfaqqUjSETO4mMXPFC+N0yjrrfl2Y1w9CvD
I0XkKxClBFTvHZjIsW7sL1Zp3vdXiv0rBsVHffK2/3rBfj+d7AiAdU4r3fR3mtHX
6jow5XISo60zcstKGevCCe6A5bGOPoEA14yKRvsF6GaxePEasPtxbziMWogiikeB
a0xNW4wgrhYZpbIgytS+mR1FZeRO1mhW389yt4VfjkJe+5EFnb3iBFgDMo6qxP4r
j2ozhWuVl1qQB1F9DET73aX4AyS6y5gk4gaOACVyme/tTjp0gt+wtCpEqVhJ1PF+
ViDGRzVqaJPy5WoNS/MY55mCA1U66ZyEIDrD1QyeBvkL4Z3t/lFxfqqj3jlsYMAn
iEXV1VhlHuKPB8nDgjPRjpvfkqSw/Upp4JH8Z6B2OkrCgHWwxLMRGg6uk+MZWhoV
0TvzSTi4AF8oIITzQecsBXnd/O1xXGYzPAKH0yh6gJNLuMhnP9mtBJ8/CuSZli7U
ZHSUogwBbRHprfkQJcD8ZMxEuI69K49D68T8BL+m5sVoG0JNH62E26jtJdB3BJH7
1d9c0v4X+tiG7IFOxfkyy65XDhd4P0uVvu26ypIfVrvuNcqv3SicWy45mTaNvfEh
r7je/rTBjOh2N434Qyu4CsyfK7aC/huQdUKjCY0eettIGfx9218H8sskBWL2Ec67
Jed5KdIhT3OPcmNwf/9hqLzqaEFjPMgobrFacsiEhUQf2l9l8tCuEjyH7AXn9TD7
IyLYzDj5wGLNmiYtBZpvhFRAxaO1se9Rn7B7Lobpyabjfkk/mw04Qw8NEywPksJG
0fVetxJ07MT540Tt3M6Wi9AsU8lobTHzgtksFHWA9fRWwPUK0EVwiEe11HzsZmS1
7v89Wrrol6HbBeTqxZAMEp6YW+WzA8YwiaNGcA9UFfOIfo9aCXURsco5k5vV9wNX
52tAyCuCOxLCPnjSKuvr4D3pPqf2yjRVjaz+4sQTIpfM6aZmHHPw5c0BiZjBFD7T
6RwgCFoelL0MP8kiUP8rHNJB1ZCPNH2AhQYC/JbdAOWOFpEmj+gRuvCVJJVWnTRu
0AI3/twt2QDg3UQcb6A4RfTR+hHAuPsMsmBDWep0p/kBu8Up8MluAD5dGkgJ12DP
6uvH4fNp+ImgqwUNAINjBYDIrua5r77oWJq45Vmc+G/hlVyvqgS3QyanxWrvcwqE
mrEv/wzupfDxwUv6kzKQo75qTG7QloYpUgKwk7+oN1ZlaITWV+zLXlv0Xf1UV/Vm
CAded3gt0KCn8c4d6sCEtu+8uQ0hT9dEMyrrPruUY1yj8MtmFIoq21SFCS6SSfmT
RSACCWKcYzaKUvcrP8vDZwaQlEIriApVxemsqZkPke6nalvCh8iKZlXM9hc24Nj7
U4cgzmCaft8q/crCJnm8FRpoACmhCBIM5sdpT3/U2IDWykF94qaOyWn+WHruTS9O
zQfSLg9VqkW69b+O33zl598iAVPVtDiw/Wh+brIwfYUbgjsaNs7tZB11MUUo1RX+
QreZl7df6o7MCzePK1TKOFw9t4mbUWM0uwFN1gccNnoJbc8AVstHm/gTF46fIZAH
Oq01BgVQlg+5RZOSL07H+I5shJUYcnnCrbzUbJsnYHZUVnQyNmI5vCbZ/zXjOiTl
fGgoLjukEJf9K9PPvbov6xjMrhr+kBLsWO5RHG83sNn5ryrHtugfMXdeYFbwi8oJ
wVYBmNTPyAGrKU+Fufmu15eFoTQeNUCep8aBRwk2/xDWFTux3i/qUAJ8UYXc/gS9
U8nITh5S75Zwzg1nujZGpVKi436ynYK0figJCbfgyijchRxGTbTtd8U6MlvaBOHC
aL2JDdB8u1+2z9rE3XrHRwZj0YX/EGjLTRRljHimuvgCq925RBhZ0+bqQClhGA0s
pdj94NexcZC5TX6tnHjcjlL0Q5vZigXafMvQNmtHCsPLhRtnmLm6MmERCm8pqxtZ
pBBXISWwCpBb1wTQ0tej0NF/eRDQN8a/Xiy2DPEDsVGRWgAdjmj1vrb48EOcRwn9
CefCBMl23hUkOTAACVdW5FUF+dDDN1oiWKKsYZXIl38dFZIS3GhM6OYk8oJdmmCE
RteooQlibX/uXoK8FMN4Q/GQX3pSPL3zMpmhCskvEuDroH7reyHL+DYmSON6BFYE
vuKnu9FpqqbojQ9UMeO4aLVZYi5rLkz7fRyTKLIxC/arervq6RcMHgKurLMxKJoG
w8nqe29mZNerFr9JgsRt6Zah3xV9Q/KiiBC0+h+yoOHDXzKvXJEFlJiPZDrHLxkV
KQQQld9dHQ+Q3QeQWK/rR4G5PZuL518KSupwRZJREnfrwG8rIocZhPiCpg1vQMKa
1dHRPb7Ud6REakhQHLUqQ1SS/elwz9HQl82dTeC7ZQEhceVA7QZv10rjDPDQWJpJ
l5gckDoKMzXpMJ6ILTevAQY6jZMqt3t2q+WIry4HwhA+nsF0pIRoQSQOH+voo86h
8I2YADNiSGWMLcNYobQT7/7BnJbIzmYjwmTCbkRHdROvYdLLaCMBY7g/212kW5OI
4byDReWIpzgqph9lExXlZlIqVlUnNPANAFM/1U6ghq+djVrK7277uHsnx4Q9oFZF
UfdI1eOzs4BZ4sRmwEmaRaf7cpRx6KuBDrET5mj1UHz3trb1SXx2KsHi5I3PQoxn
no1BGvbnXHlJ5qHMpzUo7XGZ4B9lqJLd1Zapq3palsg911qKhuvyr+jBdMkZjlMp
u2IDf9fkQwTKZZz/SVvlcaLPukYilaYB4D7s8MooHqvvOzv4EvHku1c6CdoouIih
f9nh8kkn7HklGYuhg/BrvBCF5oLIyeSKL0ZG6WeyJ1sKuQQkhTImPgcgZNN50F5h
WDHI16cJFl2GAsJXwIwbVAivYXGlx0I+A0bTsFMG31XAEY0ym2a75b5sWHAXDY/z
liaT/c8OUddMDeF6Ml/8+ZM0vMs4VVIqbTdrS8m5X0VtEnVPeROn9hxK6gtgJueg
sPt0s522ALpCUU3X5QK8MtIAeX21L53CJQbKViDjR/N68EyeeTl3koj5b7TaFqvN
N8sp7OttuHVeR0XldaE4j5vt/NEnzy/RoA7HZQjUmD3/B98nkVA4OIvuOS/ULaD1
mEvdGs5dwxbwm0i6w1Me1zqri4FFsjtl5axzZ0PyQQvBIF/4Yas5ulx6ZObJ5JPC
h4p8tiJIhSGa7pqzljc814n16FEA3Q3n5cCcC/3JmHeU6OUdJQoDh0Ue404W8Ja1
CUgMrFwV1rroSFEYEhlcuJfkfFsECexsy2zEkU5EXYgTZ9cQ/PJZ+7yqPyeVC52/
5z8ojbVqHFjegj5RMon9eGCVOQGx7tSGn5ml9B/X4Uy3eNNGYjxM4l6+oX2Un0O8
F9e5Npindzt/zY3ux6nrkqP8Ra51sUKjo5zl8yeJcZFaEjofHrwjdLQzwPMYDQeP
ZlfM6DqCW3Hzatp8Mh9O3DqSIiaVYO7jcgUJeMucae3CBupHb+9sbWIeAAgQawLM
m61a1OxfiP07GHtnDDzNF5K8SnWKK1rpFH4UAgPaqm8R5EHJDdidaNR0Yg6Ms8jL
6r14MamNud3AgesIunjcseACh/bWjXQuPgr9nrUU0HI5VhUGPYlmAECNhG+nhFWM
exN/1mC8WcQhxhxfD3lnDFXJsX9W093UOUBFhSt7ZsyUAW8K1YbgDIozufAbbUSe
MQpvID4kP6zF4PsZToEoVsVpDVCkr08LWvqHcxwn2NXco8OmfPnZZKlBwo+Qhs0i
JEY0WgdHyYNfsm5GIaoRfqphSyBCC7jMb7Pa9+63xl/XmoWjJS4nL/32zDRfUQJy
ke99Ny6x5LRQamADcslGKR8pTIRsc1S9s1nfxioDUJdFmGRYfeG+vn26xAC3wi8X
yeVYHgWAu7PYb2Kueg6rXvGeSC4Z4OcR6bhg/uSIehfqho8gfRmgSAq4JIUcFdqH
3+r69gflbnCLezuNQM8AuOWCWvld+IVf4aPjzl0ylbrRPclMH5WRlq1rSrsZg+7+
r+P+AVNN1G2a33Wv6Bq1GbJ6h23SJm/1QmxNu53fRMtVQZ0G4D6inNldVyhpG64A
i6tZRc78DGATAYcqFu0NkzHSuDGtuWv89Sp1w5R6lfxMsZM5X2rPY5FDJCXFFM4K
iEXkaZiv64wfPBxfd8wmPJtp/mI6zNHR+8PTIauKBZuK6HnTtxCuYz6uvunF11E0
jbrPLV1svVtySKsiI8+GAqf20qXrRn5Fm93P3TPmtnMpYB6QzBpY6TVzOfcF3I5Q
ChXZDJd9IuU6n2Xzrk/k+6IFYQYiUVBFwg7RUTxAe3Nayz4U+cKttS+XyPGkJwVe
K3ZnACyaVUQhqz/U1Ad7wRHFCcbMtjryJXmrl/1L/5sgXI9y8bqJ9frH6y3I8EvS
E81Y0ySQ5TWxtyLkbf36lkI44bpdOUdEyOcT7TQE5DhGzAS9Ab+zfiWGYugsOVjL
DVSf0R27llhFrYZaL/FIK4WK3BeVP05Ia4TmA7x/BxMOON15ZzrkSSlGaPVQMOPL
yT3pej8+vG4vb9tJUMJqa5wVwVi+HJ2AwIWQZ7urDroUX4yvnvrK/3rs/l77SA20
N1cta/wRgTvyIHX6cTF6Vr+ytiFPXW07vythnEeq5fK1e2iYlHQa8MRR/yScJVqg
TNYZsD7UvuaaM3xYKj2l07ynlBj4FmfuaQGG57AaEVEFhJW6eBJVMae8jqEtF7Un
vHk/fBoOpfQbTH1OsklSmZs9TljjU8QWKozvGQ7iXFF2w0qspt6FX9mnhJBmKqOI
vT9I1MVFyGBUuxmo/sl2qA0ZgaqP8wHHBl2IgJX9Fq1GgGIFa0wkMO7U8i2TM3q+
rMnRv+pwF1HzFDHGpe7KN1rqgZKHX8lxCnQuVNCZRmAVw+KoIU9rDmfgdo8MiPzU
eWxZ33O4Vuwovz2bf7kCRiyiU5W8/EhFTM6HqjUhvW2EeWij3/Ne38/a4ieZYElx
rBXnC+vK1srCvJFYSeFh1ptHOGYNAgT+GfZ5VVVa6lTNbtw5WL46zuQXdkUa7Xyf
jgejLFzN8hkqDEjlIiJ+DfIAECqJ87squeUK3ZA3urLPI0SukmWW3uU8bDEKst6t
amog7AKI7esbbJKzVUfaHPU7ZSGrJtEyzTwobCXDSvoVrk/fqCNcrpksgU599AdP
yiK6HV3S+Jl0ua0Nd7odtCXvLuBfKt1ebqYU9GX4L3sYuUSekGUdknP/MwWai4qR
PWgmu/6M2hwjBosV5dN9HOHrQPXiDJiB+w+W2/i0nLLDSZZa0qD4+0U5u32HMaR2
HAJjSnVJget5jYlQbuAr8BGhuK/QYB2twb+oYyt9H5/1CVjIU+Ern/AvufkFVMQe
HvC1YbhmTR9aGPoOZ+g0iN2EgbtXJ5gYjSz/fvnXYH9SDy7z/ULun5ijBgNnZWGg
/2zuljIIrNABER79BxZ9o8lgb7FPrHSsbgmSVMouRHSXapBMqOiyEMR11G+nELOv
CP+8TaBJtUDpr5lRWLHryq68bybSEUXheaD7jHM/M52+Hf1cgY34QL8VDr8kYRbt
8d859ZT6bNreG8q8GP1W3wx2lF7IdzeDf9ypfqrguz63Ck5xIIM295sJHlGENKMW
hT7YKfnYV7gRPtyy4GSaR3eLlPyN5MxKO4fY+Zfgkis7ciRWF29P8ScyLCObIafh
W83le+k7Rx8k+rdwumt6h96AU2gFFroCQJxNxm2kB1v/7yqa5q03vyvA5bLXhceV
g8jHW7sBTnSrS6K58mEjayMiRAOfD0hYpcv854iKzAdapBJRPhcGr8R7fnGbLEEC
6OnoWP1iyTXSyx+t9IBEGHdUgFukA3bARnuZH6TuGFeuGHxNW248s4V+dPMvMXAN
yZqlkEow+cjQ4/UuLxsPvurE+/N1aFhb2vYLe1K20x/2ZiC4eXwfAJhrp/PcnJ82
MlCDfgVulKkGjsxA+nyc2pBsHn1uHdtAtiADpE+hnsTSVRGlg3euj5LzcC0JRRTz
5/HAF3c7otNhwxfhA7AwKCJ/bg6ots9vfhEijr2bCZDTLj4ub0Wl5BoWK+RPwZrh
kr49U6o1WFKoiONhag2/RL7TOK3N2CzB2eMYVQj445zLxN8NQ8so2zw4rQWDjA+q
/QLK8kDiVYn6bxeM+ToXtS/kFutvBUiNBLcbKF43oPSpGUH7eaJOEJ1FttnJZedj
A+I32vAm8QBPpwXZpzh81RgQZlpbnEg8s+plvUd9e0VPdUzNXnpMO5UGwd3R1Qpz
MGDu10zMVjlLzX1do5o/d1RqrF2a94E/y4bq4sbwkGIKJ58qTZvYFa1D6fp7bAur
uPXCERV5P8klyr4VV9SsS/0EEHBE7Ct64UN8m6mqvgzHdg8ND3lVtr7Np/ky/w/W
LExcWboDfjnd/W29fhcN42Vcm2L2k2fhnki2whxeq26CCG1IGn88D/4EZAND5STr
rHHCXUqiknksVrCzi9OImjIMvxOWAQ0tqm1J4jrwYBJzxyHb/i1DxkgGOLNUfAQF
KEax+efj2NSkPhNtyChiMVB0/CqUoRKYcpps7/V9LpJgmTaQFgEiIPy4AA5Ng44o
MwaMpfvllDTlh8x8uWOnOyFYiIem2WpHpKSXUB/MdJLkFaEAxN99j0Uy+py9AYQt
vBRy5XSnGsTxSivyEGozA1MHjSF1L7Kw78VCYSXLPWXRSIPgVqTzKUwgr/xB8zPB
BydsTLlf0nccXRSnZHWjQFqA07sRDl5jRjkMB/mOlkZgh+epqeIvQMxrgVbY6pr4
5ApY+tPRTYbFIIe7jfEdt0nZKVlSrWXesXuCbE8dQYUthKa1Foul5lRR0CMKEDs7
KQLxni1+oNEeOtGc/dr9ktI5g9QzZLcPEsq5d9DpstwXgNx/yu4C6tsJVZjXs2lZ
tJpMLv6YPLXeM092wG7Nola+rX4IMlVg1UjB/abv4O6ioWLBCBnAMFYvJSmTjhm0
OQWZ4jXihJUHKg+/L0EBHLBAA1IJwQsZBv2tHpsyUG8OfGTD3TNc8CoDEJ/LMy04
1KP0VnTBHrArujEPhDSdcCSexP9/sOnDE09jdoAGPgxInNJQGAxtq9pom9A4Rz4b
dDkSR3cz85rjj9fI6QHIB2vFibiO5RNAxkz6C/IaAliPCGYfTLx+CfC+GvaXV+h+
oj+yEdDMHAqWbEzCbFRbL/tY9aYlvTgVtrP63i1zC7YtNe4PDjV/nuMWiUzciVXq
0/trxT6QzNcGh5m7Evoa7GXWUy7HtnQECLUWmTW9+nErgbF5NPsukjhTBJpahieN
wI9cKzBP9kPb4Xh9xISf3ghATfXfpPDymWRYDkUr5sQ1LZx58FlipJSufxwwP8jJ
/hi9olc7dW7zT6aPSyYdzDfgnUEcD887DbOQ4KXNbSzAIHt7a116vAOasQAeHePW
8ogW8TMTxgp+jlTDsAqgH1k5/aTfY7/46JibyzKMM+fL0ahxE1QHAdCtthkvnaPJ
ynjG9d2eR9vhA/pZhEi3aBulZzo4FttUQeJQumJbGlOPg+S9lR+OkmWmDEFF77Hf
Td8fC2nvrFxKZJDhOR9yZFnNsZ20154JpGUDcrRwprqtuU7a86PWuE7YXqVEqJd6
fGSg6uBcyvLWKAkhuhTb+DmBSNFlTIWadgxCR8xUbukmgJt0pQEyEp9p1cGbVjd6
NiG4s3Dno0+GzIdzYEqygGZzL6fu9nfkBfJjbEKMyue3MuQxx7AGxGf1JxCIuoEx
HSedpY7rNXySAypdvuOQCILg6OGmbf7Vy8ohC2XtaMPXXp8E2ec3pk6y3yUlW7WT
pbVrq7OHzfz9VwK4IWZZsBFTiyiC09u0deNZlz21CRAwuSQzamSBIJtCoYxyLJGA
Nz3HEiUM3ew+KxLmBGqNNsS8HkAopXyO//3LGufNnQ4STAyd05eYV9k4B9vLMEj4
6/Beh9DBLcXE+Uxt9yxZFuGLP+BZogGfW3sbig/lK0Z+Imv7E8vymBjZNssKJzq3
9bC/eQhQhrO/7VOHc8E4ZvDdBSXjHMbnEdU65SJAO44V38/1NRa6GjJGkGTOZjMz
eMBCDTPQJjgKl12OxP8NEPc9RjluIr23G9C7Akv8JXx2Fb5d+Ph+IwCOkTTHRBfs
3z5/vDug902kqwu4zZ4zIJokrCSEOfdexGZ0BDs3BXq0NAQA15KB2oe0vMvCr7s0
fhdstPiecFthZTZ+osNhd13NmnKRftCTsYonb7PCFb1T1rPx9B9S48H3t8GcTHEu
wdUlahjBxPLACPGcsKeqLlarSIQ2t6uAY/hulNGtMqZo4SZEwEgeLHgxZAM1rA/n
Kqv+YLAG4yd73O+YP0brJvzVROklKzJBAfl4wSSmsAOc3DUaGF4YIQu3jM6hc30u
QqfZOss+chY1fYJPaPGu+5R7c42tBf2PpJUn5b1P9FfKSM9aakZKBuYAQan86+mz
0LobtZPJrq2klutiVRCBkCCFAKpkWAAwFa2JrR0HOUIAN909e7YfxatdJPRb8i9S
IBpJXf32XzYpq3MvdQevwrd9czMgpJ9ztQ1Yt6+XKfKT/92ATnDLP1qh+2gHdmsI
WIhz0oS3q/AF8vuO8ruDAPq20VkABx2NjrxZUtdcXGTf/NlLKXeJsarTJEFTT2Yq
XjT5qp88ylyJuwG+k2g1fnQuPI+C/ZQ+sO2teg9MnrESwYEIdtjqqqdj981iwkDS
ODRRzN7YBdf5EY9cLr9Kx2fFWn0Ycdv2jPtNjl5NaXdLIwrUnexSAxZ/48RF/cNG
l31JUooYMStWjMdY4Gr5bk3huieT3KwnLkbr2cKC5M562TzGv3BjSSlmFNM0VkJQ
Jbu0WPEfn2Qs1QLRxrlqsNLa4mHzxA56LoB34zzuo+wiKqmoP/bkpFFEOyrU0gBn
PTDQR+5tZfeAQ7N4DV+jhzOlAPdZlp7iUWQt2YNuNJy0hcSgF1ayMphsaUznf1L9
H2dsAwFZFDxpL/3t2/mHDIXJGYunFIfRBBAq8WLhUrQg/aVAv5BNekN4JTV9xL03
P/D4F9XpBbSG1Hzl/t2HpkR4RRxNPzekAlpfqEo6Tumo5je1QWvFVCPeTknql7Xg
V418HIbyFm8u6dxPpCwoVg4jUd6yfsfULvei+6e0GKeC2UDumA5wDPJQFXM8bF8B
7zpSadoOrIjyGSyX9n3JKthuhZyhP/wqPydRPotju9z4I4UOJqA93SMTai2D7ebn
qlDfXPMIuJdp8ZdofhLo62KiRvs8KmWEN40bMGbSI4RGc4uC4WKy6pHcxig5H1hn
Nql13PwFqfSTttvWEl+etmS4rmFuYQrJbie47uvBiAv9Gepd4XQSlpNK2U8cAEga
AZ9zDknwszqeHMWYsFvEtsAFsaMBKdMns9MqiDSlVrWhjGKkU7emg725Ic98Kxlq
hahZ0VX5j8KPJ1VlPwgR0ytSr5Gmwy3mMOwf9HWerKTeeFeEHg9HKlPMFLKvB0ga
YhH3NDbNKWqV52Bi24kuE+xzx6U2Ol1USB2uPqo3nr9lKh1eUDgG4dRrUikQtcKl
XF6KC+vqjEe80EKlyu17qNIFOak6qsfmiXW/4vMYBlZlhU8WQUL8LcJzrG0oQJu5
58FvlZoqgjEyE4NH6svpvz1UgiYxa8lMcVzeCT4XbsGn/rlbwh5Wbe9OiEgifAuD
S5Hlc+KIMdeBHf9R5b7VBn1b+tEGMB80Za/JrJvvmAbNTECGIzmAH+IdSLci0iJd
dnrlW5Xm2sB1B8S35e3P02iqG3sk+OOAMDGtnFI3M3LRrGDRCQdaLSItsabrlOna
XAPHm3Slt1dqumZYapS2DlYz7cUChEFZAx/x4Ir/qahtEcQHgCx2E/uugM9q5+GZ
eo6O2nyvTcI/PmwDLqhY75wTNqUT2HeuTvXnzVrgPjXHY3PSKxhaXgDD8OgQpYWb
shVz3afxpEU8PVu8hhd6kgVnuICxxnSMZbPCfs81iQoDHMWH9Q4HoM//LtTQDrej
Kpau840PPXje5ns48fTd7Vj14TP+5EhJFO7lDgd5BV/abKoSV2OWPxMSxDxSqLjU
Clo7HIgRDaoEn9wnLZ00RV5rzOSD1J+0S8czgSGduK+TgDz7Xd+ubTkGzS9AJxan
g04A5AmKx8xbc26NTr5iDjIR3xyECfWsJ6B6zZ/PYpud+H3Cldwwogdb3TltW0Xc
uGrcGeQo8hOx6WDleJomVr4F9lKwbf+wW8lhwDg7F4b1Lb/S3GdS+DTHtgWNCo+6
wS8cGbdfvi8XGPlPoMQRaXvKv3zZTcf3tsP7Vf1GGJ16t/rdYNlCsCrH8la7yPTL
n+tMD9poiXohvOLG6vnJh8BhdxW+muX8B36Rrgxis+oJgqUvmG77MQLLZ4n+QRqb
GimgVJe6wPeWqfg4cDldwi5Q/FXCHGou4bpwymyN569quStaKLYAYMPNALiCLtEb
dOVIkUYHg/QQlT5rZkUD3IFvL8AnTz9Ff118AjOdj8JyH0r8d3Vq7Da1Mrbjp31Z
Z7/+jNSEYA6w//RgvwxJeDAhfaAlWYEtXrvRYhbiqY6LJpMrp5ILTBwYMF4cbiy3
2uEEZ4lkthdmdgK1EwhpDUA8YKr12T12nGG1iAsMee61lhqR+dgqbifXzXkljG+A
N/pos3Sy1mm9SCHtQgprLHfyjTR04XtEKAh7oZrwbU114smu01De0m0cJF4kdKYV
UUOGezcYuC82+0xD7iZw58BZdqTrjoePc9yFTXhB5SrDBHZaezjHrBHDKgRC+egr
PzULAdxe1b0YtJ24m9oawPx1CX6CojAbzUwb/ciPkZj5jPx8Y+HDmyoa+ddkFFnq
Rkmm9ZtXy5i6nPgyH5dxXjDzlHula2klW0vpowpsxqgg9kFCvdOVWj7Ao7QSxrhw
YmxiYNe2eybDyjjUfzCRdZ0Yih8dhzqFpBwHBamgNW4XUMU31eqolpSRfT4uSzYV
U0MxAa/nER0Dq/GziICrueMMAGme9Ax/x8HkhSW48mn6TFJEk2zVkjUhnZzdrGEA
gTuS5yLkmSKWVBIjih2ZfCNb3VWLrtzzRSPXO5ZUcQml9888wxx/2d+jIqvqzkqN
kgozcv7Ysulz+DssH7aHxKa5GY+GuKbL/bgwqHNCNq9pjZIsC5JC0NtzHIbYRL+f
+7s6jErth7zIiO4nZxAXGbsoISU7Fv2tyH61XcXshFcftqJpfNJKF0/qw6hsm2Jr
OlCAEKNJUGXXDhgTT7AbUp7AmW/EbU2h8zSak39JIU5QdT4YL9VszuLC7AdvTMHV
yxvccSDfGrkRgbZeQk6FKlYOQfY/j/Sl353Pegxo8qAg26WBj8gIGLX5CT7JZQ40
9sWviUxb4Nzuma2a+XxiBgfmF318I+4JAgWwg8obT8Pf++Ll67LwqrxAEZPZs5e+
yqJPa77bSWzDYMVq5iF9k9kPNMOKn1jjMl5jrRpCLCICbwUbFF1gkvJAuQNtxMp5
JNsn+uq8eB750Px3laghM/VY72JfHyE3DRgU/uS2aiX5VOYhJK0yz/3c4y/h3cZq
ZrxsEiDhr1V1FivWQz2NQ1BnYPsdXZPh2xHAQXg7niDB/vlJ3fqpMb1IMgpKnfo2
80GGByPCgn7ljHVeKwbWyD1rJr+UwPTMgdeOxvvGcuPQUtOlvC2gnM8BAf6nrpj5
AExwmfd7xDG/8V5QT0nJkuRufvDIM/KquhKEaaC2Pgva5BLNnZn7HIMWlC5EO5+/
hdSbSL6+KqcZseQCi2OYJjOj7qtW/KdCZPpxY5kqGXN2siswNgBwoWcqvL+FxwhW
j80N8t906cEtCj/r2jdKZUIW7E9FpF7c58cUGbSB58xGJzObKXCHpx0NYP0JBYGj
nZ3TpsAMUGXIm5/Zc3vhQdrvz6yyhNz5iEYq7eWEp7J5Wa8b5TxZ1wxnN6W11jpS
2SICkfDenxlwbcbuK5y5gRgBfDsnHcMRVP4nUC4t+/RVoRjv/NbmWYTcQxPH+9KJ
wu8I7rRJKf+6V8nBokiK3TTLSg+s3HG9PaSZ+B1ISyDACtlPfuZqHVKZqN8ZU5eo
iAmZhg1V3m83c8EylOjAnL4AuqkbfYG093f4udvSyMgOevVM7sbgwBUEK7eSk6tg
HNBU8dGucTUSzoiFYBZ7RAfUG1UTiBHsJ6ycHAQE9Iami+120Knq1ykr9wMbKIZz
IdWnt7FkQaiCBrj50NWf73S0XvZfWUCu+Fmo3W3BI0y2iC2p/IFmPGbbl4W/h9Wv
naHWC5TGwAZjotZ5W8D6+wabapb0T2Dean217J1txS6gB+Iwx9O4ze21Y0cKYqAY
i0+GQjUsIzdRLcGwANfP0753tmr1GhVuOgXcBg6jhhzUcxaxYxzXiB9deKuiyTzk
BU+KYtMdV4oC/wc6OplssefFNQJfwI2o6oznLWuUFPNRxUgCKzBRnmPj/V/kcrly
re1krxA4TijF3+CyZv4/y/8vCLJPIf0xCR+cfWZ3xQY0e6RrG0oX/axh9datcKvy
aUBPJd6oXgPZPmxp5yJbZva0/4h10uav3rYabEP7j34QUp4lxm6h5CZZdEJ8CEGU
Y+YZG11x26vRfMphlS6lgcdCgySwkecKPIcXfcHAeE8g0U3G4lB5j68vXZLrSgah
NjoVLjkI9k4Us38MHzR9UpA04ihdQxlIGhykE2auNJ7jqiI/nIqZntAL/KJe4V9W
voHO2YtNEFneP3nh3sg+k4A8Z9Kmumn2n/X42+zD6a2a4eT4lituUGKdUqi0xjNt
61IkyrvhPsKpXDfmFHPExP90YRZ7hglZpupioqjmbNBm8V7gZUgIaQ+BKxVKDtg6
qJX8cSqsge5fKCuQm2DQIeB+EtHy8nIuRsn4ecwVWUg2Ts4bOIy0IFgkb2lqY3o9
UNNCsjG1wBtFpeWcJeeyFyy90v9PS5yyaU5jgUggr2tBJDF0Uo8yQ/mVYcXwDkOl
z8N7OEuAByg7LvEdtU4IraReMk/k3xNBLte7h00knzBywqZ5/WsU0UTdznTfuVK6
S49OHdUZ/DfVwgaR8ebx1n0MnZRmxwUeSDBE3d9M+PAkljJ71/AUV0ZQnSWrFdkJ
8GOyOE4J4wKO+widCvk85arq4mdcDXkbcmpBjm53aEBIVFoMRjtieBWF7zHSaB98
wq40NOHVZAUkXFbEjl6UYFFKR1k4sLfIRT25O5pbfp6LZMhjCyI/SCHWyjqj4BCx
fBOS3jbjfmqPvIQVk8YRrTu2oxDNhM5/Orj32jIsCOpBQXbDG6c9tdqyek7atucJ
NgGKs6F8NH5iOE8O0r0vaDEtORDIXtgwl80LEbOK0gGmy7xKfWlqOohobodEvYGg
Oc5UOdMA+l/lhbOEZ+NFeVyrWof+x4yH1kBl5/K36oeHbU0jfLHbTvv9z3ea6mxm
ikIUXuTa7MN3ApaTvmxiolJDeUc1HawQgtdzEyMn4Qc2yu+/2ib3TUkF8HFet1PC
F/yE791yi2TqhGJ/139XdB2ccaXiSuzZFH98Nh+Q/LTn3QNtElJKm4whcAfOnSqx
yXVBAZufKRvCbV9hb5d/w8o8XHr+8cIHtR0IsV+Y8VebiKL8JyXRDZ/mhV95FBdn
OUoSy+TcrsGJuwnmm3oskghIV6Afln0GQ9Dyrfj04wT97cgScSALCEd/1w0k0lYj
OxTqPFBYIfmUtupC9e1tDDhR1DeUAvLM0ESaqdPPbYNqeyhtersCAoGWwCAfWmDD
JveUzJRPgwYG3RINWD+TlUdokQgSUlBoxMVYPfDLAThpENr35ae5HOH05Wq1/cDI
0M3ZZqQRQcTDuCqykZEl6S7VHdXcZ6ydCXFAWMGB0dPdBvUdyWcnlEFMCDJjyyME
DM7MJt5sQPU4ZoGN1R6fcersqR7IAlEFQNrBVENfQ22XhMzF6lh/45hkqgkGDH8G
JBEUjR91hp/veM3aDTN4B3QfAW5lFeEN332DQlwvYjPIkrRUX4upCapQSFTdS/jA
PAFHAea+Nl9XemGx19Kug/YMzq7k92Kw4/wkK99fyHxe9uEkWDKEyu1bq4bQYse1
2JRr5vudf9w3Cn+EDvLFXgwtzQzRdmi0yNm4BunD+v7njDZd0YuDDWG5p8YWWcWF
bPGGgELexTwiQ6pE5AuXu+ADIFX08pYFeOj9A7diBFgWbhorJjhCkknQSf4xGhxq
PiIifNxUzCEOYhzbPalezPQmYB5nD6AGGdinugoC2VlPYLolbPgVzQd/eySsYTje
aMbA3ukvzP6oZ3ZC/dbVxGiy0AYLSpLb2okZ/InQdwzcBiH1U2JIUIElo1t/OfDg
IKX8xr7JPuxqlgngPKIRM873W3KAOlqEDomR43j5/2BkuwgjqV5i32wXQIwIzWU7
UUUKWiPw03RnNCCteUcrUXLd2/6hP7/xFj1eCEN9Cy2rs9BrGVTyKHHNlmYILZdV
quTAeJ08tmaa7Dy30ryx+yKRrz7WjhtE4+rpWxQMgBDvrQvWm5HLPLclwl8XMaTQ
tk+K1Pfp61+ZzxZtGeHllK10/vWFoCQ3vzSHv3R2wnSTUejZm1rSS2FcYXLpg8iu
OvsDTX+rhGuzQjLN/nBk8r4G06Lc/UnaW+0tndNyc7EmjxtXv4cijpBhY7jQacYh
2mVl0R3IlnsRFInh0X438WvP5eGici1+upIzdLkDpymthV2HU00rUwe+ElKC7dCe
2Dg+9RK9ki9VUF1Q4lr2oNWKd0+1c4JfTrAxbPIOPwUNYvTv8zkJXelmr5yAo4y7
ClFGqzuYqbHkBa3yTDA0DEHWl2BUlJ2LgdQFjuHGKHrdZ6q3r/TfqhkwAajE3oTA
TGcLo8we/zgihklPzuxoTvKMOTM98nzrO3/ngAQYR8q+XDLkWrHk1L+njNT0gOhh
iHAFvjseXd0fSIS8aE+p0oyZOEBx2k0TwyEGwNb8LkSphfz6qwSZxIaNJSxPN57c
LpaYEH0JhOAUoYhLF+g+QCPRXmTmYjqAniGV0PK2OE0qVbdK8rRgmkIGlSqXB5hl
XaaO2m1gHAV+dJYEunTZHl0J9JX88iwIe5in9hQxsGAKCL7jWH++ASNzDuuglTKu
N9BtyIOf9zVWYrNiP2YpWWMZ/RhROj4tPpSJaDZmT0ygYgc0joXnj4ZUwujx/W1s
FqYRYDwfNEK6lvAuaOi19DUKwpK2DtCg2X4OD5tpgqiGvNxwC6ETaSpWYzrgvOgn
ibqEg2OSy6mcSRE0Axiy8bXgrATiLSl9QdCEusqjTTGec1AJMV8vm2FNASqazzFp
lv5BtnC02hIe/mdOkGyakBrCqrl4yGLAvxRo5T21ARHcgwdGjI2XhDdlsXM2viMR
JdoDz9dzsK3+DFonPpR9aUN7e8qk0gKn/K7dM33+3jg53lPzESq3ZS6Ydixyg2qD
TvVgErZEWj3WBdlYM8UFvbd7GpVwZi9ye9N5mUQkcP4IxePWk5eycb82PEsM5Gad
ATnGoks7LEYvBT70pNqwg1ejQ1sMy6ViDZPee4P4aDegF41cgESfCnaXC3pJ+aRn
I+msbBgzR2driYWKfyi/yh+HTGJZRSY3pPsQ+YzPSNnhHiZPmusH2ToZjmAdfgEx
Jp2JqW0Od4hfFSJlF9c7/Dz8ulYp5sBke0NLXz9ZCGfW+sEDlSpDpeENYWHJbkDL
Chz42jug4TkZpJRE39aOa3XCFQi+MlXZg6Z6xmVLzjqVY98jjyJ6CA8mXebgVFSl
/7CZ7enXuJ1+vMix+G8e25fTuUt0LUCIJC/txMK+yB4B0kinHSuUa64Gci2tGhsY
TWRIekUSK/zXgKgXo3JvAWL/Wjpj2j+J5ZH7rTWZmQxUqA/b9DUMv79Dap7dgk7A
RpzizILMdf1W14JtGkA0WnwXeuiH3F0LVX2HewzPjFEh6CO6210KxZZBouFJXaoY
3M8inT3eL+6UFenk+Qc5C7zwC3ijLbsoAtcNz5erkcqwCckPWawPHKM6vWNVdoAG
7I6EM9+mj8qwFfttZjzD5Ny0VmpwOv6rPybI4tPQGX9uKoz3Le2n58iBJ+1mDoXN
PtEH6vmvQInOsCq/ESruH++BllxNe7qde/0WGcvad+F4f3hpw2pr8CicYUFrivB9
sAPDNs9TWfome93vZJCCZX/VXbEc8ub3F2qaAX3XFZi6Gcy/1kjLviOjC/EmsPhs
vUVC/oSbY4pFIQ8Hdusgsy94AXqZKBu6fShemTVdr9wX931Qa31X0C8yuAufbuxv
19lZk9+wQicGgh8dvO5fjno2Cmo/vk5AQ/24aI9xL/IXHnF3/N0X8Hc1kWP7k93C
4wXD6hXQBVhemfAwVbQ9JPPpTtOvrUzZw0pgWN5xmIkEjKs1zKlyhUWdxuLcc9Zq
3lTiXOXk0BgBBV71vMyaly7Gl5QBqBtdNuW/qUglDCvHMGPyiyCNo6/iLPd1OkKz
33VtGl57rUFgtXssqpF9RqcgO3D8zYWXaZTaxPz+21osATCheYZv1UDpkdmIlONu
tjM7aTFtzXZi4a18bujgTPDcVU+iyqJGLjfWjSCYXPxp5YNzizGAkwFR95hsvZo2
CX+ySGIEJscC//SLxEnxw/YAr/XNKIwsHWEuK+WNvUOLi3J848zX8yDzE5EAV1fx
JIFqu++TOlMhFdJZdenvZv59XEpQXXiJPagjV+HiCdlpPUyEKX6N7Xgrel/ROp+U
3xONZWWn/9K8M+6cJRijx0MrjekYJn4YUAKqd6ypPzO+HcN7gYPg7zMkauwVaRfa
kFQmZ3lpxCr3pHBlXThW7ZTLPUosnUnYGmbM0oN533VtV/pJUwUkT/Ys3abBPe5l
QXto4M5pV6uk5h74j5/4/5lmQA5HlaUCCjwI29yaiRa80rs+bCtQKO3OK47Nd58Z
nPHFxmLxSdpx+8w2x4aK0sViKHX3OxVNzdP0dkazLX9yGr4g/RR90B/9DWniomCd
I/K29vQMUqVaVuWHLI5G1ZQudThfRrifSmbxgpYq7Bd+TtGwD+RZeJmskl7akW7o
aUboP4hI1KyXK10bVpGMNZ9FOU9UGngNgM9z7usFCJFIwYBQ9B/XgbTSTJ79baUY
3+0Mzws+qYL18kti2EbZx+zXjVtBS7x6YrBuOQujZyDYg6TMxyg8QFhLzvRkW7Rg
Mg9AsB6Jocv3AYr9uEd38oO09z2qjj3d3AX/ulgvKWIoPWbu9qJE5LMeRMZ/bGoM
SIU4n/qGkf3y6wGEanWVuwzy2JShhxxnM9Cv3xcP6U/N6NAB/rMitj+Sa2N7zwBh
L6cNoCZwNhjVRuc4CnUQWzgZuPlD+LC/lvV8yCDLEkliX/Mec4kyoN9GUOk4f6bJ
MikO5+gycQAe/H8TVX4eJB652tKOqB52GuNYCw0JCZd/hW5hnc1NpsTnBIDjlvoO
q/jcjqH5NXjWjmjsNspPmjTz+M7neNrtyf7iZXwSOki+QMoGUXXO4OiX6+nKV99D
C6ReCG89eWNiBePvFUk/1YrDwhE6wrvVqZkAvyUG4Qb6Wdult4sDhBpje6CqgAWk
0pjcjM7q8/ayaIDejrYSv8NJhLK5tLsBMiW2/5his8ELayYx0i1gbdLcCgtfgDcn
bqbhatJZ5OBCuMgXSza1lqMEIgdyTzMb446hMto8tyZ/HrM9ZghVNfUX33iIKq/j
bhBMMapTBc4Vi1AaRV4yFKqb7dQpPhiugLM5BAXBjniMTfFXmH+gcvXZn5Q3oORN
DyB021n0pCoXUhSCTMFh711dZeRuZHruv1ShjjZuimYMtuinEJY9D4MKOUPAX7ae
n7BrC/xAV8Lp6pTSn8PoHz7cMjFfTeeK5jv+0ciHcZ4Grxb8SizuHsIqO/ZlM8s1
6IvYgNlZ6SBW2BMzJEUSpUlpuGZe5tc0qwCZLyGGzQ8Es2lycwC1zvH3zg5aFPhO
wppCSODbJwwC1y+ktnNwpCzCUR3kQMNFTklLpopY+dqAo93+U+J3vvZ07jNOGvjt
2yondMQ8W8WBx0FPJ0hzyjtZ7ISYqum1L2Iuz5RklGOXEMapDNZ8eCI7zspMfAPy
Lu4UtCyllXMkLvz+3IoC4Sf8VosLmrqr9NVHiFx5gMKhkukuRj0CSP+RttgMSkWL
H5mEajbxXURf5gyI7zHB9Ya6vYquctAG51qEXedQdb2BHfMjjsTzIcsVbh1v5oem
Dvb5A23TKv7P/A5BNAEbFgby4yqYEmPZ8BKupSZeOSOkfXQ6NC6LBkwEoPo2aRXF
n2p6RKEQfVf1/kAl9OJu5FpK5lKMoDeWJ2RszRcBHY/ySrdDw1YTmro4bfYEcJMi
EKx9kecZOxYhASLC3ATdVgPsUCM/WQAVy1UCIQqTJoQoZRxX+taa7TxHZlWDOWe4
Qzcvtbla4cFKhqxM2XLAYY1WI4a+sn6qM6kVrBc72iZk36JsnZ8EmSGOSPyW01Vg
LhAeYtcil2hgZAt3S1yq1DG+FLuLOkgOaYgMhsJAC30ASNbx4y7ixVOw8LzVuAjf
XB/sUOZCjIjQFaSaSPr/1y2O0N7nbl3m4QTfBtd2BViUdmO6Kgdpl4NaQWI0i5iX
dGpOWotudGlqrSgUcCF73LVtv9oTkPa7SPTJDpcoKB5KI+MfSaqstr6M7dfRKOop
iFrPqpp31H2qTZ2IKYDF90KqtWSMuwM0Dmq2Qj86OwjkoTFSWrr9aoGmirHWZcbY
nHtVx6I+/ubw+cmI90Zv7Sf6DWUQOcdkwn5nXnEGD7uKKYp3lJOajMDw43LFtT7y
ywpnYX1PnqIwqdyAQ201nOQ/Uh6cgwKSJCgmxOq9YIhk2HZf2znAR91qcSQjWbQc
JHzBl2e6DaS+hdsd+fZQkEWVVj42oQuh6cBTE8YOqw3NTQQjxFY2C7E1OeYEMdk8
j+b9vQC1BK7wuCsmB1+Homx517+nuSiYV8mZ+51uQHQPYVMKPVZ2kJSG1MZUUWjd
kt69GDfCqr28f706lQrzuwSFx7C6N8koGqVn5WzzMVW1LnyJCtMB4vr2JUg2M9Jh
tE6/fRZPPvdrdYv+26q/flxkbD7A+/W/pROkkf+sQ8rwCQ8k1OB/+2oRjNDF0h9t
3QZxpkusScG8FvqPUcaGiKE45xBPQrqYQwTk4sLsjNkh91qE4YOjIuplgKmAeOE7
N/8RCFsIg58wMjMLwBO/3sj9OYdxRramyydYLAy7rp1CZqjhv4qPU1u+KmAVxitQ
gAHh+r4Nt7m5qKBIUlkAfFLXaKb+bdOqlQBVJLS2gJ+MjCmwgGyZUNgr3ieUpCGZ
suDJaT5sNChioI0lD7ACO75Cf8c4FQY4DU9h5Yc6Vkk8ZVpO9mkkX9JA/cIld7QW
u4+flZ7xw1smQfVM6Tr+hy6BzIS05FhpodL/yKYXF/C6iSJuclh6QRrDHFUrFrTW
UD99sxux39UcinIFhlhvRgN1eV0c4CHYq9qXIcvqv+OiUDP7U6uDqF8ffPZKX0Mi
tg5qnJxqNxhs9VuaAJCKYFA/N2IYMH7tWDAV18khFXj2iHItcN56XLwGIGdoaL29
DtNcIlb1CQD5TEJTnOoo/jKMWr104e/3Om7Xf233WJqDCeZTD1nx4jud6pFfoEb1
KRQFghpKMYWfmEK8FBsLcg73KqtZ0z+OMQldTl8lcgF+GLxEn3YX0YRWFHgAkchv
95/Y2jfN686fDDrsghr1zGTQ3XYBFGbU+R4GjCKZmXuVpZa3FaxMPwHVV8y7dbEH
EL2bVaKwBGxRwVa5pPt/tbzgC9urz7N0xSDRKOaCJHu/eynN9rsImZ1csgCcuIiS
ULrzY0tKsbfub1H+/KQrjTYDvB/+El/9OHj2foWhyunXZ+LIaJwqselhH1gfVltT
3LqtEN5aEytw5PqGwJclcr4J0v2zKslww57OwsCVIGqyOdsfNlOO9QKaNwL7EmdX
fSQEeoJdgOYV7jeFSobH8R1+VEJc0vt8sEGrXaJBu8n0NKyyJSXCaWgHBs2m/o/C
3Fp1qLm3K+8Q0FuZZtC0N1ma7dZHkRtkXdKoepjg2zB1ziKVcJrmV7nMA44s3C+q
hXHKCAVqLSqkhG5+7cwjUU+sIEb+/wuvJCwVtsLP2AAj6g0tymgAprZmeKpJs33l
QBEcJn+9IKKu32Vm4oI/z/NDAqk8HT5uXbpquxkRDv0HIWxeXoKUJ7eDnHbmNBsB
ynF3mf48imWprHdF3Vxkah1zABKCT2dUpzwmmI1GvVzbxwRC09olJvDkyyVmcii+
XOj7pt+zg4oH5dV3WClSY+IefoLHSUUPoO8szVwqL08/XvivU8rOw+WlGub0VC3P
iXrR9Hsoi6lLpXPNcVkRMuRFMdxi7PqRvxFS8STJaogBHtxSV8id69rPz4qUDp4q
7lXa2hRsAnp4ACgZJ0ZR/3EQOHSRncg/9W3SL0bFfnY8RijeV4Ct2IMtR1u4cX/8
1/bwufQHYgqITkdu0ORJr43uWBC7GDhZRzxNyZOagbi4er7oYMa7BlkvJuVZ+toO
dxKbBDXzheykTJRezavsDPXCd+bWXlQ8UdcNcDOp7j2pMRoZmEoY0i33oE8yX+CS
+fozyJRNNL6mfvAZL48RRywwxXdHy/rkV9TTyVdaXQhUIPYha/1SECRL6GVbZrRd
oc6DJmFTLozXqNSILHHJ58ApE1wF7ob5Ht8J3892VEu3gTYwibWqBCQjzjvaEXsK
iLIiY0V0kGlHlD3a6cFhI5MtGR5EUzQ64vTACSX/cPBb7QI42R0kV+n04m043vz9
zoOTAuQLrDASXIPhCNyXJd1FZQrrnlNns9RzdTogiLCci2mBEEtkJOQhFjM+TBP4
5CjExp3Ea0+5HL4Fusm3ptMZnlb/dECUqWdsr6SEjXHFlLguUWOwT0AsYrxYkflI
xeJ1dP+UAIdAlGXseGcE+wMRDckQ/opKRjj217C244kY2ceBY9id7KQ2eBH+w0lg
EW0rv2iHrCAFz52JJiy8V7W2Yj4hYE3Ch1CNyLHzX0Rj4kHpvqRfs18iQ1ZMGHFe
NPa7Re/LhdanHtws+UFKxSFgaV5D/hUX0QA708+JttivArjaZrNDyivli1uLHwMD
Le+lCBtjSPysYExOe1zAvlZyLinUw/NRKLrT8luO8Y7A3jGENNAMm5GX+3NRSe6O
3hk0w5Yc3BuQOzeOH6sBiikKgtpswFbPj84P2ykmfOuhlS1vFukX4MT+jy8nHx7m
rUoBsHcj+bYLYFsVlCep02CjXK0dEfEywXefT8Rqpd62J1Hy5HCJDLoVoEbNn6gB
LUVujxRLlPllHh9oW0rLG87dEoCziu46x1Aq4PDAuhtJC6wgB6Ze7RovIZvCN4Ba
+n82An2B6VvVS9QsoOEr+s9xg+7E6taGgZ0nQpx+P+9xOMQcw3bYTNUl1QYgGYdi
K7MXCi1A1nLQ0GHE/hxRcfVUQrELzK2UO7Iv2Jubo3nLGpL9cG6F6vh1654tfNJ9
XqnWHZYbBufRfLEfNHX3gBCBxylVY4vGnZ6oJu8fgPTV9/cN2aFVDNPOMmu4y1Rb
GAEdGotFw7M7nnYJf1YI6LX81qX0Nzp2Cowup7jvrudU5PIqUNmYfuzpA+cXuyVY
Bgy8HnF4aUgIMjHGiZcIEvJdBVqDKxDFGb9f02vYjQ7YhUhq+y1GdBFLpjRatRTy
E4j/FYt2RvPdalDCTwpk1tSr11YpZP5I52L4wQtO9RFiSO3aiEAR1jmNo9Jb2dg/
gFhfVr69+/ta+PVBO/JjWnbZ77SBMCaPY42x84CmKWoxdq5SN3IX+KBUgIWs4ZEu
cvxw9+2fMpl146utUHhVIDtPUF3dHVYT7E+eN3D3NXJRBTHV0IBocFoi0N84cDMS
tv8mQ8p0GmKR4jro4wEZwENM0FO+xyVmKkyeQ6/CV/vvIc51iCddW731OStwgLeJ
FR7mt5OXQ61gUjMt+ny3kCt+G78503xVRWdORgcyaPlOf3evF6NTHt+79sg8jN3Z
MmDXrKytlUr93OswNRMOjppjqpT3N/vrfeUEVX/sNlbXFMpnG350SGHfdgh58/uU
p08H4tJuSdz7aVEGy5jBq6m8umby498bHtW5Aj4UVg4xpVupKHGwJbyw8ZkgjAhw
MAzTWBdhi3k9ejFD4eF14K+XIVmhYNpdHErapwfBJgC15QuoKgFNwzFuxbhQGDk5
rwk32HJttQV0aCBuTFRnqBE1FEEL0QLSaP6oLaRteFZdRE8RFDvW1jy2mjVbY6zK
GOVZoDRPzC2ZdWf9Z27p3HLoNDARvZJqqAG1ISIafwXVOY6u/0/jCF64MXAJX5M2
P6D6XUSpYEGwv1Deh+CKYR7X2mIyUjvK3wcITWGej7w4mjwOqOHQL9GywwuyMrqu
Ale/IDHNwB4+XzlZ+DuDMmmeXvARbR4l+gXeIdR4Car64Lyd2YXA3LUfNM9KrBsx
DJMPpdAubLtMabI9LTIwvVRPwm1aBsTOm1PI/TYpKT1Bswnrus09jF2d6TbYCyYU
ECKUzC69xQjrI6hHt4L2CM0f/rua577x0XJbftnPxNuUpzDJgM+BWKJPVbBjBy9E
UOkI6+Xx2qHmJFkxO28j3WpRjnl2fttjalXLLtmqf+p7zRSh3kastxUty+4kObF5
W+0j1CvLaz+bPxyK+6wTB5++dVCxTAxkgo4Z7ucalP+sllqFYQdwTz4A8TSz0tA6
1+0DGBFmjcvW/ZJk0LYDp9PwoLNLstFPctyGbSNtF1Hxe+8o0gRD3tkus0TTIbAd
Oj/e2c3CTwAqzBEKIwfaACv7wCFKd8G+knFqSZiiNL43OhfVAFYAk3CgLOEu6Dtb
9berJQUlihnVuamhgLnLG82mUFtefxwq7EPKh57Y50Wi4pHlNb3/elkeTGZmhIMO
Cl3TClH25uGapWtIto1aAj+Gih4YEy6TaWDXU7NpQYiET4qir4ROfosOhNqzP0Z7
mqW2b0Jn5oV2NbNXy1lIoSPhvSnlZ6UW8UMe/TBA1a+Vv2ws+BR7mLZPcL93q9wu
anke/9QQ2jiFEoGy2cIu3uvJG2jM1Y4m+A0vLKgOGhfgduISMbuBVu+q5BPT5l7d
39cWB5LpDIOBsi1V8OQ85pLI34PRRs4ISLmvxhYi+81fja3LCZi9i4dLKrzH5N+j
1EgCxFLV/NKIT5yjqQIdDRCkjYDbWA+Ralb6be0nPaK9SbbSHpc1aAv3Og3/vU5e
YsTFHnONjVbSiJZdawH6X61aIsJniwS5xfavdkoEuHmy7fhaPE4PPqaSVmJATnQY
CjMghv7mFGzaHSyXXO+hDrR9Ye48fjFFkWQ6qvUG2VBWe6Sym/97/qhc9cpF/FXY
21jQ6K1thS87rgbbg3ryXEq6j1IfOEKSwqZHGTrCtd5kzyK5f4Sw0Ln/UAexoWgJ
8CPCrnc8sSMdQg8xS8+CJyzcQTxjNJskAih5c7KI5jakQuPztqxiJWLEQ+gOgWoz
xGOJhJ2PrTMQNchw8lQLjYScmImkS416j7fKPMHGLlIUMQcPLV/ExKRa2lHFj5K+
sU6Q8nYz1NniP1Wg93Eq9y1bVZ3b8v7/BVM1Vrg7YzIRcwSP3XtuE2URaW0e67mX
qrbyjNRVew5vzNYTinJ/sm8KJ2CXXpLjY64m3h0b4+TdfhtuQflbZXJ8EK6aa3QI
WGaqIP4m28BAw34bJJYqBQXAMZtMTcfve+FhEwDN0pfhfT08kWft9EUCtQOrybee
1XdyL1bcjLnf6dPx9wV/0rEHcAhwnAAO6qyxCflWLL/anhqCuFpKS3TJJZKQH8YO
gt9+LfQp91ZFQj1fwgosFdyACLJJ3M5s0MiIGrSJ7nHVArJZBrsDljALtnHugul1
iUGv2UWN3X3dDuHC88FpBgTFZKKNJMMeZgMpQxZWioGhDls3jRC85vCzEK+iBoD6
EqXYOYplXAWZzaPqybjbA/wZCGfW7y9qhJ9pKMiX3EwHtBP0u6XKSG0a0cm5I0v7
+wCZXc6hDn/bhls3oXvBJXIh8EGaDcr9plQkQO8wHoc59NrpSekINYKBJ81AvxeS
DGq0bRCS/mp6MUBqhpfSTOTuC3xDo9Eylnk6NG4xcWMe2qBuBjZdLBUYJIvkz6M+
+9OTCR2W+0+WpD1hn5mlweXPOzCxgLoWCU8kxNR6lm/F/cKlBoNG8a2Dld/3svPO
ACvxNkA7bu0rc411onZCCP+CPGxQj7ksWWhBmwk6co8hRdOVzeY1k0rT1kJ7uaX8
SM26J2PVQNJBHWsuWiqJVEgg/HFJYMb6UgF+qhD1mBhL9O1DhWMwe4ICOHGEi7V1
+FJvIr4brSCJUJRDzby1kEbMsI1Ivpkp8PNuIcgFtBDQRbGYUgLXkt24tnRZBN5K
j7ycDaGb7bjkSFNmM7Pk14+0E2hKGW0p+LINs7D1XQsz01YqyMIs3aV1wjz4vKN7
wVIa0oBD4hY8FyN6P3s6qcv6ItCJN6vuEkD4JFtOp/dTyJKpFEFn+D5RiGUUDhoP
xulDc0/n1w4bmdawrlTswN1QwbjsO4YxGoosTSFWV423oX+SmJ8pdw/kB8h1LIb2
IvU6UNYVBNOtFU+tog1GYv337Qn4ZXRZoAddX+dbt8Q+ucOp01ALFiY4KcALlxZO
/tlYbZ8m4YtZM2I/jqbMbvgT1+eVcZ1wXbx7kkW+q+3bUL0IOmoRt87e2o/ORIOc
InAC60DVqWcybMg3rYZ/atloW0ihnJl0lu819C2LR+MxjCPlI0M7BogKXsEJdKs8
E5aKfWnPfXmhHkRlcHR9cIlqQR0sixHHdy8TGcrD6XmDFxln68c6Ehmzaa3+yaKC
hdjuV2eYftZt9BtOdALB9B5OpEwiQUobm7Vj47+Bj49G6oqEOtj2q+a3rwJfjnbo
Kbjdnznpht4DQ2vpKE935PZ4oj7I3DBsuCa8ACW93TZs7rf8oC1HbidU+N+Hco1e
H6M02kRJW1gQhhef29FaYuK4emOw4NPCwnqDKIvN4maTizIHZeLEI97Cz9k3AJPM
DMS9kQxanXxUzUMK7P5Ye1N53pkoHa37gT+/2S/JDcOfmUKJCP2vJsf2I6iU7WSF
h1gct5hz/IFgC6+j51QFjF34zTJsgbHB/KvAwccgBvYMz/4Dl4yFbzaBaTxqpCpb
wB4eeEMtx+cxc55MStm7wox/8cADAy5/6aElF3QMYqDK01boyssxHnI0B7f9BM6M
r3cwyhIAAVjpqfGYt9LedmfrUu45GQQjNyW7G5p9NpnWcYksmjmgw/FMSbDugXZp
35CjlCi84m0p02PB4D1nSNIEB6aIv5cNimvk9M2iZyoof2zKKM3h6f81rMyCH6xy
GHEW7vJliLHSAr42XCY7EynhVo5fXT5+u5b0Dgep+Oj/KYU2kC8UMQUel/POnpJc
sOrlGCZq8lEwGzfoIYfa65fU/WjENMmk9UPYOr0rI1C64Up5yld3s4FK1lMidC8n
00QwZ3Kzv3eqLg63YOBKWSnALjFaGaliJkLrQJItIsCVCiCEd3RiHbOqOnPbpA9G
YO2wABTqCRrLdKg6yIL54/0ZOjrqw1oOqKPCwebG6jA/wKzdN8YBuUEiY7DUT2T+
TTqZQ8IdTVPBqNs8AjUnrJ0KVrzSD3oxcF3W5eQEi3vySjJCAWi8kGIsGtl+iiu2
Q9KZ2j/6GXc6apDFbgLa8zFAAIG1EPYBb0/cTl2en0Z3kT+J8tnojg3vMoITe57N
kgLpJsKLFGKM/kfJ01WMblEx9CB6TkzMSMjNC/LMi24XcuYb+O8HE3ixNY+uoTOZ
DIyuAv8E/kxOpfN9NZxZmpzDQfNdA7FeRNjeiVezifyPpVLTW0F1FALtmtL1sWyo
ExZKDBkQvGk0cLVIlKt8Gx3Z9ApVE6rAdiW9ARn7TNOj6gECbjfoCnVBPR/3WtD7
Wvjro5f6T+G8Y9l9AK/ZFLPY+MsYnz/dL77d723Q0PUg6PnNjL74jkxDSDt8Zbbm
RL/ZIgK+nQEfrzUOjfyuM38dC86dYzrk/d35awxvMi4uwNiTeEdZpGBvf1FPFoV0
J9Gnwgf9SziaHgM4+H/EOixnW9qZBL8Kv+WV+7X4HEVzX4bWfcmTMccCr5haXLpq
QSbc93qNKKjVgV6R725ntjs4SE5ZyUs+F8m2UkALqdcy/9f8iVxJwfc4dn477EBK
01G3QTx0sbig0xy7Z8fBiHZCA4YMolQ7p6WHyoYk6EQNcC1lK4Pbg2JixIjke5rI
EA5PJLOBn5ikrqRIA3Mq5KpM+TPS3gn5sEyhAceKpauiiIzMzWttVK6Vqf5sSXfZ
uevvycr19EtSQi9E97aYvy1P2p9TLoNbz8yWcWIa5v4+V1KKTuoNBXWIo4zLZXYu
j6nTYYd91q3cJ01KL0r6LAE6FGX7sgAp4mCT/H4c4P3yeVtcYNcLvGvGsaA/TjzC
DJHyqYP/W7SLFN5blVHY0MSjpEB3fayKC5zj0eLrYFXLeBISRrx6otSlFlqCVV0t
shE6XvSS1iwzQ5fS4zx7EuayH6t+BsLLZ/40lOoyjM03rFgcZwnOhEAy3EjNeWnW
GYti+Vly3NmsUyV6eTKL1GDd35oqFaL/iErRbAYC/avSj0IDNcAJTCRnxC+m+WaA
08Li7+/9QEx89KiMciIxRbDtMw7M3MI2048Y1/QSlDlVbWK22sBLuTnE3RR+ikT1
ltmUdWuVIgwyT/+09fLZDE36llYep18zpfmOMl2jBPwGQ4DbIvtqMKDDtyM7yZZq
a0knmX7ftZXvYwbXRPLJevYkjju5+jW/FkdJuG3pO5h3eacoMJ7xIKOHfwRaY7HO
etx4UQboQL3OIaDEYnzRYoUEi2Vk2qBSwzI86JBldHloWiYqH//IADJwmKKLJ3Vk
ZAKdGKc4YVK7CJ2mAg4x9OdqMmVIeXuTATYm9SgKEAf9/uLE45+utY/QdarFzSID
Avfab4OGfleX3Ru8ygUV4PJwH9TfSxjN4LIWq6zhOIKWIeLmIDcRpe1wyr8PErht
eMktFQcMl0qbtNgUGsGu8SWGay3WjTwtLhRrLS16oEpz1kJdbY5vAGQOg3YWZjeN
YLoRCR8qX0UMoR020lzsUcAQALbnT5DLWa+/4nslfwkE/q9py68sFfdUD+jQ/Yhz
mmPSlg13cmB/Myu68la5NbYYfRkb8pvBfjeQUSS+GyqZ2vJBlh5tHpdf2USRM1JK
P+jDTeYe00RqzzzKRLWX2UUb4r8mS7wywOX30obOvzPj5UJyrt7ThSkg2JInLYLE
EEBpMgcY0ayGK9AT8/BLBQx2sK9lAyQ0KE+tL4FrvmzRPppJK/iZHa7LvihHY4F1
3tSDxZPCPHNAFl+8R+Y+biNh2qfWEoW5YoKDCLL+YfgkVhDJNMahkxzzdKpklTtG
wtAP+OSzNBPfJzTGIDQXsnO4rk46iz9VcP+NCNk1ETuulnUoANFSpSZrbFwGZdQg
SVlaF1aBoqXVMAOccEbGjHMU49gianz1WNtPa/krSMUtPtWX4+y5l9tyaYZoWHON
aZcXhg9h7kskA7zmDdNRX+RKaRiCIvVs7DDbl8+3fdQAT0oXRjTqfPqyvMD89gqJ
SURIPntcg4RL7zFWl6taMyM4bbg2OGQvgWi7Z1Aug0hPFKhx5LmWsRGaW3CrWrC5
WOuU8ZfoldSn0ZrhehmHlrovT84UuRKfYrWLq/mg3j9fiCMv6+pMNIalUKgqLdGQ
EZWfuwfmEEW/nGQQSlMO1yi1SZu4dn9Gys5XBE0PhXzkrdZ6Si5xG9EkO8IQ+rVj
uiZhz3zbqt5589aEs108oxDGMWz1L4gd4bWV90MFT7IbfPYSgsMJ0OVUMy0pBOoi
JQZL20EVpJrc1IMdeGVoHMBci9RSC4pCz8bORb2sdmFwEtQBN4iodGsYCbCAyC/l
6ofvyPwxd2mwcvwYLIcxt/Vytii6ycrU192V4XDqA3QXBk4sCFB6qGpQCJrQMDUA
0IYJjZK+TGjWIUqH5gTphkrhX2upVQYCvU4182/ETzDfYwtVi8DyVxGkOAZEd/9X
AlPrBowvjMV2ZBA7bFe3kfvWMKH1niuBEkWykdnEM7zsA1oa/esyvvn+IWTz8ujf
0CH1bLrMxioiUTp1PnLZd7sfFltJXw3qwW2fGcYqBdZ2bJnOfrqET276+H5dIRkb
aske6LiCj1FH4ZexPfafn/nOV4whGFoE1pzOOFvJr4ZZgh5ArhQMW7Lyam4hCAsl
4PS+SI3hnENQ/cwhX+YIk62xWvJ78KWwhSoK5VrhAvey0jNT/dVV95LFvzFIYzCw
4t4Mn+hCSdyP+l8onfAe6cqkiGCjcNgxcTJtYz3919lMtIa4rtYBbExlo4R9YAao
6i+rb0x6kQTiUeaLIfqVTrxEzOrMHoNAfT7qdw0OiQP/68ED6/PHPUdaxwe9D2tk
1Ki+8nluNx5bOMRyMevGMfWY583vcTc8QYjA2DjYtzpduAzoS1YXKb7Mlk0GYATU
NkMA++zQ5f0WyiF2oCAI9ECd88G7UuAVquDtaQYeQvih3135BZ30HyjlyzAdaxKQ
bzG8uh4zc+/M5vTrNMf0dCwd5E09TEi24pcDGWFryaab691ljmhHKlw6VsPYM7G3
JFLbayPMSBMDoqQMZUE0POLJ5ShvH3wBgFb7O3UEQxt3kwl4v2VWpOcLN0UlstVT
ePKCkb5v41N8B6bn+pnSW0XlIrrq327d7mWru58w/2TmKyt68fKdi53zeqMshQw3
GoGj8rMH3SK/2wtLUubSMdVGwaVH37I+DMh89rt3/bQb8XTv3jzkeuWVvqukhnfw
xPkWsSnljPMTEL0DFnFJNr5ld5DMTt+hgbLOPmYgoBM812O6QeM4eg9bL/cF+GjK
agUBEhCY6GnSNFcup7f5fpHN1cw/wBKs9k1DunHHPk4lyrQSVSy6diOGw0jPRC7i
oCcwchOUWhuliLZUxbf35zf61cJp7k+P4+6o4AbQb+CR9C5VgQ9IXWi5ZQCzNnQQ
oPzrPArFqzCoTpyKaIlMEJQGdNfxfKdvWG8uaiOrZksrofd3EPYC2JKGMt0CZdal
PsXjMmMdFd4ep8aeFN7X0ln/6Q/sh8nfMLcsLP6gy/R1AH177LLSOwYmxEb8Y2E3
7xiRZpzCQUy3qVh1LF3vPcmYEH9JpKfzV8IQKn5m2loknDsnFEvRyL7mT0HIRxTm
91EQIG1mxAB/+fVjxLKMYk7hhobFVJbk9JKiIhyvW7XKqTSECFZdAfiTrMxOZqnv
MERQWIGoZ/9FbMj10dErw/z8bya6CuiyWeN6ycU/sMF3uNP59ROaYLLxdZZ1FFCe
JfcSLRDUm1Zi7s1qoXP8AqFnNqexI67HcHUDeMove2KANRpOdu0IniwdqV8xRclA
rhocs16gJx5SNZKgQlZpUPRobdcbxKayYNo2dBLhcSGwKF5t5GYC3kMEY2VcGwB+
5et4MiVNhIQlNqtfAvvtxBhiDO8I4x85oAYmvTtUxbAwepUbOm2iu5ToILQPi7C5
RmFeycbjXA1V+qsgNA9M/ZowAOu3nviJE+3aErMBs3JoFbMon5HEhKHPMOtb2+1X
GTu45qjRuS9081FUCiwQ8f+irtIQ4Ln7AjR0gWw4N9ejE4zhVnEeAyAG8bf2v1iC
L7US6v98T66OByZUBET/RoEH7x1O4eYvktHFTuzWG98a0dVx4MxdYxzhDHOf6W+b
RwLHI2VJ9/xQdGyYXSHdFdFCWjuSsfa7NvXMIxLpfQJcyC6HVzw+7d0NrEBBYOkQ
VHYNOf/UK0w4oEj91jUekNQxgRCjqzWwyOMsr2tbewMP2eyJ3vnvIKW6YzwBYXNu
gcVyfKkOwxPTNgO4xxRkLLVqyZznJHcLRJtB1tVMXd+L1xyyUSODMNDOkbjtDRyj
ZeCiM7TD3C6fy378DoXs5wyEHs7BwUnpazWiGHq5WYLZMC/IPDtfKMiD8y39I1o9
DHHQuPtGxhj5MWtk8s53DqpxUMuHT3kJpXBs+f6p07xjR379dGTB1GM8eYbTiTZS
nAbC6bG4JvdiZBQLrZambUlesdU+G4yGPoTE5eU5FSlWiPlQhTaxD2vA1x0gA9i+
w+aKx6M2ZtOkQHZjisces4alOs0bwpS5p6RHRUwk0mPqyuyBaHx12180NZN7OPtI
6386SKM+z6jHfVouUvBwavH7S4ynUtZpTgqkT3SMTYVKhySjkt3sgNuRwE8JeygW
GU9Y+cihO6oCIvwnxcU8gPPK42zJgbGQQbFW+zdNf5wZBmyImqJPs+FT81SiAr1L
fJbT5t3cKUppKgp++SRPK2x6y34liT+VxGxSmd01b3OucF39T8+lE+Zjf/PfDlBF
IJIn9dj0zUA6eFl38yjujwW4ww69tko5fqPbRIxmYi3203kQ4JFN/fE9Vfsi+lYp
QEJKXolz+XxSyd5RsAmeuVlv6eSz6e82b+hZi3flKbZaFstVbe8OzMTdEv1zVQ5P
IRPvy7IOJFMAg8cywuU7z9Q50mCyzYMEpmsEJkgEkYaZbffLzzskuBeRyk0SP5sP
PcKz3FLhlzJcWbK+r3DnC3O+MzHgvYPDstlwfSLcB+RhbVTdBOt8XPxPRviC6qD2
2QBXyw/UffjA4+8Z1h3FgNXO0OAAeUOpV+7E44qGsZvaGt9gJjdYEz8qd+wLu4Td
p3zCR8wkux+V+FBUIOPsGdrmQljgF+GwJ5tR+XGeK+tYLQ7PhKhnnR+gNQHGnQBz
Ho7XRtAIxyQBo+Nr/ZT3MjrXGWHo/dcjqFar0xaUuxpMlLSETT7+e8y0Wg1WCWAg
5j2CIyBptLLEdkN/ZWiExyOpCYBSTw4wg27/C8fOfBPLHtY9TKDyH+4ICBaBLrPm
8K+Rql1OCJNJxl+NQ9UWKcfLdfm4r1kNcMjud+SiRCDcDqaSmGl2E9oXKni2Mvtg
IZCN/Ubk069XE+N27qiWCFPOtD5lwDrb43o4fNWQPk1y5skdxreH79T7ukFUJLPa
R8fMvkinWeMsenUFaau1v3t1ncSpPD/huGsRA3k+VCuOiotQhufNfz8MBJ344U4M
Zf60Q8IyW2z1sz7EYV97O+Pf+rPhHfZC/bEDQ3Ykq6v8N5DzLeWrFHkKjbSjfLzF
HpTpvojXZNeJPekMmsucOS80aZ+4VnGO6V1f0wh5A98KuuNMzg+YaOjEVu6iC8kE
PIxK4PdL6V4F/E7Wl0KreVO0Yl4B2/ItXUOjlYcYOIblhvdLE654j8ABFsgtKyXy
M2NcipY6OR8UQxauS4WIrI7u6QA3XSvVJuPJ56ngRO+3Zym0JqcdQ54TwqQN5Hv5
CATkqkEX0epvGFmlAIKxHQ2FeLgD8mLMP1BCsFnTzof6fNA7tfhAM2qTsW1btB+I
EAf3Q55r0mYjQm6mF39ZdkYItEd2I9QOg0lMplyHc1PwEJWABaKHQML7k4zpEhZy
4jF9nnhSR8hrsQsEsffgIb1ruLoO/d+FmNE+DkT+Na86FzyN2Wv2nGYMy0SJoTFb
U+M+Azujt7HFo4zzbiTim2kCuOFB9ohFhG9wbmL71A99FKWXruws+f6ELlCftY+5
YsaDm295ew6HhsJ1fhw8y1tDSaeyoD6SMpxwhlMO7JcBTqYjM4yYjrWp/rn/xKbc
9zyOEuWY13gYvVCJY4QMBg3vT612eseIZ/74+ALy37veIEIUd5++IBxMZln6QQK+
MRb1lFeIknhkktyqnGXolqjY6w18m9Da41iHZZrfsIjY6BUF0+m0/kacEE26+YyY
E6n5RU2qgsQW6mnVL3oxF00+cbetX5LpsOykadOYnX42X+rVCW1XphCUy0rL2P6+
8vm048t2gaHJQ/PQNmxamzLH9996at2jayoRvMwGfBuN2zMjoeDaRQyCqaZPSRCA
70izY5q2yIFmRu/5C2sV1BaRG4hEmmbcPG3P0kGe/MFMGPSlANu4XWoDQ6ZlPqVR
d+fRstLNtVBWpFSROx9Q7d24tak0lU+myY+sPfhSBaWZVZOlIzN6mYMcbnkmzS0M
pSFuF9izhzX0ysknuphE9g+cLY6UIg9EtVxrcGfQYnLLAZspThPcyzgXMct+Or35
vOrGzu4Gy+vdCc4svtc7wuRehy3V6e38EuYk+dbcwT31xeYedUq878+VRdHvA2Fk
/LrGGqK7JIR0NyDHmYOcWbG38LH547eN1SZAxqUEaKGf73IwiGqXWwxhDvrQF/yb
v9kAzIIwFeMKbSjbcC/Spjl4rOFHIMHwNkbO1cU2EfRDU27h5cOvysrINX6TqT1y
MqHO4CIQDc82Qx9IJw6gyfPksFCUu/CFtQtL9kzmGTsasSI3jDT4vWVEeshptUTN
Od1dizrPucT7SWyUZCF1a10CV8NEzfMUw8nCVsW90RlQmJMZTEtVLvtYRvV35qD1
6pZfTp4Ji8pbWjbPlFce0ljib4Zo96BDEp+HYsik7d/rekT+sRBFw+kd8ACF+TTW
VbgShpwxcm+c2lVqQQhD8jSq7nycov0ascnbiXWs2xqysxd7xxyCXLKxiFCa/Bfk
yE2ILLx2M3VDBMYCFaoElh8mp6E+gifP0aJgT7VZAYxpvBh4NSB3bR5FOwNQx46P
PAFOfoxHpL74i4onIc+BjrPDbMQ8dGqfR+PBU1psMpYrLCdEO2GPO0YRsNxD6Pvb
/MfPkJLo3m96B8qQpuvHydgJHD9wlE8PWYJ1prCWtEldU9BDyrxUqvl5Jr7mUHkb
wCZsLK44qfW1Gr1AJ01MxByG5A4OVyqFO1AMFx+hwLLi6WFha3Y7TMhw4SlfGGec
PZ4DQhqroz3GasOGSvodP9AqcsA7TnxnhdPM++jJ4q1fN4Wo/D2x/daUs3MoTA57
ix+toKOSOrLgexcPJcjt5tDbccrhTB3iut1NfrVJxyv1abXa1wjcb7CE8UCXgJ+u
rVq8S1wf7TJMOrKtstY6K5GZzmjke7QRZp4wkkaC0K2ffJPrV3nfPpIkrk4reT8O
Wt3VtJvXxYMin1+4dYWP2i8EtrmSYi2tr6/ccOpjM9bPV0Z+pHU43BsCM9C5HX8N
UcmdJIBvusPN6tW2q1ewGL+Pmv2JyPO6Xz2sFQmHTd7CxPLPE7Tk2uPN3P4HO8Xr
RvGaYYQmbX+p+L7OeAbdzUkx9NgV1BApvUTy3ikpqaKL8XGMV9mnd0QtZXG3+prS
zWSWI5x35v+NoUaaUwB91dw2Qnv3em6ofe66RbR2MEVKlcyxYdrbfJxKCf2tSu1B
nV1C5ejGCHkdzQMoI/BoSKO2YKNssFUXOAJenmTFWq9E+9pIq+rP0KKE+mubhaqV
0cg2nDLRRYduROt1YOWI7bo1DMyj6qQOKGiMC9kLb0z59IskbSt7gVrzyJRabE5E
9Cfcj/zrSAwA2IosjsQTt6dg1F45JzajJAwhb5t0tKJgkIZ3v7ufkATumjNggqD9
/h/Z747uFhIKXda9958oVkUgOH8aD4GNARc6Q5aRN7jaT0bK6/txPyuiT8NeCfSB
FaOBTJdAUThzWJ/wk/jSGSOhn9rGyjbEujoiWv179KItZN8yziCuLVov1lEnnV0/
fZFWpO0ujEEWiJFf9CvQN9Hw0U0jB8S9+Tf8TOQ+72F712DN1/oK0CGV8ovuSPse
yKP2sbs2zZ3uIfqVcO7DLBcVbSBfQvFlXPt/7+0CcDkhzVlUI6UscOLcDhV8rhZm
Qrstz3EvVxd8W3FTRnJeJXSZ4pPVABVmK2KXH53N/MWP0T5dnNymNx452UHH+MCS
yr0+JN6Dbt6jVQxy1cw6TfCBSywn3aKOOy56FoyzXnsafr0rMBiqNqAc4SisFOeN
V6nuMPh0DXs8GqHb9I3IRigwhG+mkFb67xtQmH1F+dE1WXVjtHNRyjkW/KSVZLPi
I3aB7rEzwujQ4e7RIUndvjW7ozSzBYODBs6CZiwwIbUvddxgmeAIYGfNdLZE2H+S
gVk8vZkL9bQSDfeS0jwKNkm+WOCO+D3jBlQZxyWOQefQwSP5IDplxfvIKCHgJlxI
MnAMq/BJpyr63WMlO9RMpT6YVvJ1cGgey3kqmndSuiZvflA1kmkQ/Cj98Z0rtHB4
ewEqcIwWg4bysTgN3HONG8EUhGu27sCES8Z5tRMvn7p3tCIbn+INzQX3eDEz4I55
K0LQ4b24k+XYh2qW2QBUoQxIC8wRF8Mhik0QZG+6MRECKu3U9urwTAWNcKz6ekDi
TQ76BcquVZslDRLVDPesm5R7drr6207IeEGlhHTrooXZ3XvcGzhOvcSEHORESLW/
aVwHeO+gngGRF143RUgopxN+ukKOTCwIGVmdd6vokTYrqe78zmUvIx5PB9a8euQ/
HD3IUTDXG7Wm/La0rfSKU/1kh8CW5bFwj1ex/F0enFnH/jd4KeHzGzDVVF0Kz1Dj
LKCLZWq41LLEOWk9eJHdaSumBlbwZFQJv/9ETm2nLhPbseToF5WNM4TDpfeQGYgo
ce8byYT1AxMs4JkC/Jka8NgxYf9PPM0bDc+L5x+TMR7rS7hryZBWIcqtzI7vOJN2
9DeLiARou6bMgVUGP4ghxLUMWXzsKtyXnqtya3XW++e9hi8Hcj53Is39Z7wPlE15
hisqlygx/t0Motu32n/JVZ6kbVheCK4IqFWJczSsIcXlywFK9L5LkoQWq6LDHAUl
SNpVKqolkNXjpaJ3OVgHaEMMjhn0ew3ppQJZZburz46fWV3jmflBoyyUB7ZfvBR5
E3HhnrhHfWadaX6tpHaM5w8G0gGJk33C36bjGftZd9iHcjCbjnXze95yjBMayFvR
koY1i3eUWA2Qa8QEaLnBQPvu1A6y7vk47kwS2T5xafRudhcupMJfb2NWkDfLIhpd
R0lL5zQL3yC4PkfCmJ9njIodX4e+Ia7kyWvbF/rh1r2VHPCvry/D+VLf8KlFOI0J
LlqHENGegryqSSkPddll7s3Np7+4JRqqVdNZnadkq5U03+MKJVIwHV0u/twxrfJ5
BWYvMbAdi1+mtNGcbWfnEG+WKgamaYrOXSBHljEJuM4maDokXPq7h/Xw1m/CkEI8
3/zX163s2t/1kvyR1dswAVDk8K6ar3Fx9qS+z1lV9k7Re+p3CVx01sY2ao4QshnF
9fO4Ss/IKQwpP+yW/wSXnl9jU36o2oeUQfuPE7zsG4iU6/4NuW5O82ycsEAXZVPK
rWFWdIoBI2MYmiqMgKAqXWiyImU53DN3LrVP3TcsRxwWb35RtNAU5emQFZX5a8VU
bdo+lx247lOyE/L9VgiQvxxFqp/uOD9jJNBs60JEzjToE/ud4PmHd5FirB8eTUEj
agjCK/GPhV9EkHIkbzHtZtndEA3/ffJOndM5IrEhuMdCtnxcvVdVgGcHhxlUSv+V
3NrpaDsh3ytl55FoVUDwljKTECFRymrkUnIIddOZ/zMP+bYtQA1C4fU2c1Gu/Hea
H+PDP4f8jeG60A7PWmy/HslUTScqWZ025+J8IUVDIyqS1Et3hGQMnz1W/N8KPPLP
aqV/nO2RwkMdhMa51J25QHBMDl52GI4mfl1ZyXACsdrzvKHzOIvds1DEe3oxs+dx
QMhkXSPdtvbwDAopTRI5sAwThwgDdSUY/cKCD16eZt8cs/FqcdX2hVNSBS9Wb4H8
oT6tqGUnTtvMBIiJCGtLOAexaPCPxUYbFsR9zD8wryP8HWrYAQeJ4xrnx9PWKIGI
gBTeT2gqV2/mtyUsBZaczKrfuBQg6A3PU1NncynJDmbtqlVo9FQct8gVSUql4zVA
tl+7thL85+Q4ajM3gykJzQ2SQi3XF5ox9wc8LPFwy4BU62EfztjlUC32mj/187jC
PfaXPiGD2U8HHLNxbe7V120keM/MMY2vrzmBDFy2oalV+NCTyCU7ARCLHwdECPB6
YP3dCd2UARTiAtlicO5xCybKlxOEIIMkZhTjgv4coHJcWIxjFE9hik9+Uqc8jfjs
aeK0DamGLKD+0duTRdEK5J9cjV/rBI2qalncS0cDG5DV868CMde8ZEeJBDLJSrAL
G2AHB7y0M68+bz/tOiWE5KdBm/R21hP7Sc6I8Bgya4DHkMJ7jdSgUGQwdVi0yYls
sTszrA4ZUq80rDfQ1qf2RMU7sKC9sILMOL7YHc+GZJBzjoMV5CPdyQ2V0Ji9nh3R
BBo71OPyWEV3qddCGuHcqLk5P00e3a2b7j8qSeS4oWUvUvyMBLoDFrOgsTDHVkNp
1GdN6VjbL9Y6YdqgGMsIDBDt5PsCUjqDYaDPzynZA304MVeF2GwChPEX+ywuQDug
TaWglTL9Oq96A39wqDqbelNrRJkHXI/QA3jfDG3irure4J8Qrs43tMmLb92EPdzd
yog63mIP1MIn+E/yWAjMaPxIIVGciHHs28epXPO0i/+ToA1ITJRzxYERGlRnU0eE
wGpCIMqup1vGBH3tCq1SFffE644EdiUsEo4Q6EiuyBZgHzF5u765SI2Gu9Z7MEwT
GS62S00U4fD2g1ydL8fwxrJ3Jy1W1WPS1vFG4pmRnH1MJcyp462AbDGddR8GU4yS
75Z8h6WGXOf5kIwFapfpAbSj8Qtubh5v4oaIwJVFlkMzexPBJ2HHJhj6kjxgOeo7
ySMiYOlCm3Gxer/c0U86UDkSyJHWSGn/o3uz4SWCR37I5rQ613U15YQ+XMJEIo5L
Mh77RaCjZFr3bKLK+pwqx+qZbj3AbNCxHRNlCVAbuZlByEHgfDM1DB1NesEDUXD8
0AS37d2FX0NkhUcSLt6Ne/RL5VY1a0TCoFoYDihQLVcwZ5mue/d2hR+vPF+aMVDz
U36DlurCkGVv6ijwPaOXosPMex7eMxCnimN9CKbidZdJ4AoPZ8nMMw/nbWORNgDZ
cMEGLMF6WpROwWs6bxRp9EaaAZGt24NDrzr1lvwRDM4YhRLd7I3ilt6CqgZLa20Y
Hm3i1baUf6h+3oeRXNfwtPS0fYSzO/Reu85GbRYLFqQ3/cYfYuBb4hlYlgjJCsD9
WYFNtpX/2oruDntotRC2bMaHE4Onsd+4a5B0yNTcPZ/f824JDUbIEc3HZDX10TEb
62GfVU0rpecxFnrUO88FgeHVToXYinK6k4nF5h7fZbH7/IQtP/g2QEJDTh/czE1F
Zdm2OCivinlyFBY3l+7LPixaujAogkMttz3E23D8uN/oOTeHY4DDAZy8BWmB6h6G
yio4Ulbd5tgeacpcSkdaVP2WzrTich0WDCUR2uZZ53KWf/9Kv5XfTSs5qwHMBVaB
Zb+8RJ0d63cAgxavvu+k7i+dNpfYl2gpBV7FVGJJNkYtHxp52fnJN86y7qJk3fBH
Vhy3VUbmv/Uw3bXyX0rWuEFwweEmYQEbkcI/LMwogALfJ0t9XIDJeNWsWImrxsF/
fEzJ2sNyxNLxoYm5LcCWIWj47T/8K9+3VhvJW+z2z7G0IWSNDEdComNKwifnJc0P
CaRrqcBPEr01WR+UbLcSPsjo149jSSwwKsdvO5MVL1SNtyeCvuLDWJ7WpJZnyiOi
rl3yJZyxvoFZZcFHnqnpdyk4YXrmpZ3WxWSumPm/pNFNizLt0pP/YkL49Z7kkHmZ
bAvyNJUJKZQUdsR7Yg/JYjfOE5hB+8xwX+sICJ9BS1AQQF2+mmLl97xOlqb5qpFs
oNhu+nkJ124UE5rAOmLDS1qjffGC/xdXwaOmTXNeGL8H6NFzNFcf554CXnk3udoN
13jexQJH/YpAhsUcqG2enSbWWrvHpuzppFuLC9/sVxI+z7cCMcR/unANye1441lu
1E+adXhNMwF9t6xtS5lnpMhgmLhbxWyMq5Jd1VKJesUXYwkqq5KZcOjiTnmIuOIe
oBTvb+R2BMW2s+sEwXTtrNfxzGFN6n9h9fZipyxnjxAEGbfROLsgZK98xmwgMlIX
3ijaHmNAN4139nOqjAlTYVGR3I8LkWPlS5xeEyTV2MqmXtPSzw9rvBFgaJCiDiAO
/6FH2edgBFH6YBOyrNs0G/SOCLHzES/IK+iLyjdKNzAmABMl3RUGGky0OGRUmwp8
OsyP+DwqQgwosgKJLW9ZkLgEKIKvj5D3rkQrXiu4ckmzbjX4Fks/xzLb5raQqvO0
O1gpKtLzWFu4vyAw47fAjRF7QaYuLpmXqBAieu3304EvLJ5+G671V+yRV3/vlP+8
jXAoWIeaeaDMnMBc6gFbcGCDX/CpK1XEPmPqOWjw5cTGDAjBvYMFQZuzzr4c6vcf
tfmytdOYnzCrG/nF6S8t9tGxFMnttAxoayxOEdKDVBfmDX/PyeHEmBZ0cGZOx5Vq
X6IuS5moxOads2a7E8BUcfXiVAp6VMJFxBBiaxyG8JajUt1NyaPGOiYdypSTE1r+
imchgas1h64iu21X6nmxAj3Fi4szdIi69QmlcNnvAw9eys4OxTt6A3fQxXKnUlS0
SRbafV2XL05eb60cfOHKsmWm6jwIDFzb9koDdmCqrzxGJjruBv6q33qQJB58Sruk
Z3rWXrr+iTOoeLh9gdiv+rbKnmJEWyp2fcG7Lz52qUSdmATQQ0EWj2xqhCNe9YD0
9SCfahILwIjhIJ6c1xLqI1EfYEQpwpo6yKW51hytqdngJm6ReKGnoyCWtd6keN8M
PPMLgrBCTmOL/n4+AoYwD2Wf8qOdqNJZy72oOz8ZqUEHlMlweEVQmVIrt02R8ebo
WtgB1gqGT3rTkXYZOwkZckPNv2dM73C40OJMQSg0CQD09q0YnuL3OR+XOsfRDjSe
ggPvAgLh3L9EpKT7uxg75pJ7VOvfDN3UmR+skrxELSJkDCFiCwWWEL/zH2s9p0yP
B0Xbd6/R++4bkw12LABprqzF0RnBDu0varEYB8FNlS15Kzx6jGgUg4wIIozXqcaC
Ht8CBRX/uBFmw20nrm5e2oeumFoe7YX28mHtgd8pHGWhjaJIcQRV4xUE2GhEjlO7
J54NaAPkIFr9uu+TvznAF+K1Kyi9jvkYPTBRM7p6l5d0XBfs98YH5n2XMN/cvrWG
rvdTKtzmhs+wdvZoCs0nPzVNNWYTv8JZEmmSuF8aY97HOKud1pXnGCFqDFyQaocd
7K65mXQYYC/V3L3Hyrldb1hm4paYf+Sr1Tkg5XldzLT+7BnwArx76WMaoLOFEcCo
/2KGnyT05bEqG+GodnwxJsQvcVZVzdrgJXYhO1yYXbW2ihajd9Cl2uL+0EsxfCCl
CrMXrksEhHctKYYW7jhVS+DIidzs3g+lD3stVYVyMHszrudSs4Edb5Z49/8s+RgK
tS24C4F0D089GAQB8a20MMr2H0rsHybBT8L5tT+qZrdkfAzHcMc10yEr4+fgPc6c
1SGCW2lE0tiG3Yc1TiExnWzYEZk45BoZtt8RgT7vhAw1GIq7Zb6rpfdz8c5iPQsb
dqX6Dgol98X/QdOWsgwmz+sl2Vw9V4xaOtlpgXrg8QqnF9ymlZy3IE73pvx+2Sbc
QwZzMoipfnWjRAolOZUgIhbmy4SwmeA/Rns/+S63BqAEIH4Sm4EbI3wGfU12ZlHf
93lmzv/D/TN74Tfl6PsmIgbUUrHrPcLOGKG6Qe3famTHX3Lm1Kq5FA29fBvmZe2l
cBebI3plIY/ieGNoWcA0GbnougS8Ls7n6m9VQk9atpqvBfWJpRBjktRAJ2/vg5os
aWAjrDqmpJ44ZojOkKa8ZRqLL14OZeOd3x9Gt8YDSj1Mz5MEIpGpRVO9QbVY+1Et
8fmKnVyIJlzXPgwYMmzpeKAoBiBw6/JPoYzWC38ZJRCr+S5OpeV4Fkv8ogGbjo38
vJAkRUpGzbChQId1dnv5ZuUWUeKe/OwLDiyl91hy8TGQYZKsE4zTP3zuJbR2mdlo
0UUKuxduDIsOs6gXh+SIAh5P33XiVRxE8GMUGuHcUsCxCHvhPHBwTG6FUz9tbvxU
2oRvtpyPpsifPYO1EwrihyHS8cYcvDpyq17j3zdVfBAs+Toq2UlGM1eye26JTx4o
oiIxx5Y+4Wf1Ze9F6Z+QjRMoVYE4IIBEa62O6rzxZKcn7gfSe/egPEAPH8kRIAdl
NGmHBFBkZOyelBTO1DAqQrJJhyJqHgbRcUIPaNV0tOAu+/HdX+48aIpyFV4F1Cs2
bq9H/4jf/NQ/zWmR/iOGRJiQc0x2GO47NENqMwOUxZLhQrdEyJaLGutnItRl/oLw
pVG0g7XazcMy32+Cs68dwYZ2qJR0x8xurjz7wql28aVe40fBRIo4PE4dU5NHgnuM
8BeY77KVYavJyX4x5TvxPlxcOkhtiZpIwCky7/iu6bjpDXPM7b00rRDCmQs0Z4SQ
m+i7lDBKYVS+y7vjit3YvpP42jHVKXx63SrzW9UoCSljmOo7J5mc2cec3tpBx02M
iTn6ObjHGaWcQ20Q3KJWag3iw1QqozwByEDnEh/u6Zy+ZbyJSx45Kq+PRuWvUXRN
DffRd545tR5JMn5dbiJm/GNCmCHsTahBgA18dPuRIYC2JPpu1WpFTz2+47Pjf72P
To3Ttb7QL9Yql3OvoGxKupDLpigKaUfbqqncGKrYK5gRmG2VsNlCs+JbtmPPKG7F
u2skUtMLUDb8ReDASeG0CTVeL9jFGdGng2isgjy/WE2URlSIsl9NN6HyfixS6LDi
R1bavCxF85S6Y/NNrSDdnX8Cz13OdKoMd87IwDw5aODoDYr0O3XNQiNwAeZTWAzO
MafkmD2/4ckGzppnkodwB4N5k5VEEH0/9wy+csFJpgMhvavSOeXsjtl/+KEwFic9
96pWb/0EYRvm/T2SBn5nnazScB+5iFp6Ne9VO6g1z+nuPQKE50MABmgVRWOSvjq1
lxiymBnVjqTCNHkBbXS//z6CJ4IzgcnyWbDYT68n7EnJLtjkFpjHJRyIS4jt3nr1
zVNASQSxXNDJm/LhWXcsnEVX7bnqCt7n6YOYDJUBPQ8J+xCALGVFwpvWLtGBs8GB
yx+f0yYetGlXpxGzAvDjc2Pjznt/d0hZT01O8HC5Mt0djeLe8DEBbxYwTqZjdmw/
w0tgeYFtM2+EUDQbsmQoPFV0k4UjXz9aq22Eukyfl1fxw2YauOGhecc6XwlDZ+Q6
skV+QqH7erEC9X1lgqk/ozLJJRjCkQ34pj0UE6vRyZlKDjwELwNipiMG2wJaAnJu
upaTsN1KtgN83rD8SD/yruhpENZ2TfluYt/P/lfYrz5bE9AZBBgHcW6k5SilbO/B
06NhuwVLA1F1Vu84PXXVLHLwqmemC+CPgN2nWcXRvogoMGsv9FnMfeSdcIMkIt1U
+NSoaXb7Z/GGzzLt2NvcPZtMa1hI8w/bq0dqPZQhpm45GU9JWoqfcU9H5j+vk07a
K+FUz8wy6ZLUvPtc/Z1IsjZcp9l6nG3Sk0WXXA6Y/vWrGVUGGPgq3jPmDy2aDmlL
CUT7RzHvT+EzU4u8R1xVsURH0HGhVHuqGG3TsRWJk/9fgebUsKUiLV2wU2fBxB8s
T0FBwDhrGcKu808nCQP99LgRjL3Fa//UYJnra868G4JL5y09SrfNHhlahdqQnWg9
gI4OdP86IyuYizRtqI5BMGr/Aa0jdnT/sboROBQFdXMYAI3tVK8b278HeDep1E95
ZZpTDj0mxUb1JELqQBfi5oa5v3eTy8nWxH6Jxk5qKV6eQqE/y/DyePctU7GmbZCD
aS2zWX00EW597MdXZcizytXwqeSNkQ/K0mE1YgZBJ1pnf0cTIUVVN7jeJ1cXM/jn
R8jMNnqxeElPW2pi9nTQYSNR61bYf/wmAL7on+NuA612XRBZsBFYRpAU497+L1aA
Siy9pyYDxKC33F5SF3x6UFH63v5vBJIq2ukrCyQ+2C4ZjYLeI3FeviuQftqaM1bY
sJvpSncWmJRgmxaZD6YK+clOh+RRXR1QansCdRoq8oN3oMj63kKd6uwi6QC4oE1o
ybgLGDSfHW0X9dct82Ri8/wytnqMU4y8A5Vgr7qf34DW1qpVhYcEyc2BQb8pSSJn
sR+Y5IWNpzJz7OD/MWksh//MEgfB3Nu1SMkJNS+g0Hj0K9KGoSVLR99P5kqFzYcX
9f8tsK+PMNTxrXdNY8Slh4a/oFLome85sQnivRRbcq4DKaidXCaEN+zKdHXaN+fg
zdmvTbnbfsuFViPg34PB0jwcWovDGheYy6uicMzexLBk1sxAVtGauVlIpOIL+DRQ
GXiJ6sm76zyL/Lrmiw5ysELAeBgu75k9JGzhr5T4ago238GPFTZ4r1ypsWtKSz6/
Sq8FfG8XXfiQfSgbV7DNKtWyCa/pNasxme/j1RFlZnhia1zpL1GVOPGFhDW646ax
xGKpU3L7BMw9DvWDxIVvfFXU7/hatDcIDI9DXMORRFf5IHDeH8vgYBV1NMtsk5iQ
RL6xOSl893kc+KyGHDi+2rgwbF7NxIblAZii9k6+49pXsHsWobp60sn7a+jq6uS+
vzvVq+jJ6fCa3SAh8shmGlPHcecAg4LEL3Zfruaugpy5+dDWprOX+igTmkg6ZQPb
ScbJ04KwBtUzvaK1lJaU1QjqjuGprQExSqsqJkWZOHc90bbPhYp8ykh8PWCkHl83
S5OIk64wmuczN+A3+jHfyc2JkLD3og+ScOPdO5gMkVSvxX+D/xbacwjWlN7SLoeS
VS8J+Do74yKQtIi7bsYHaW094THJs1Y1yTziRgahL83RBqpj1HNc6KA/6aMG0H4K
mOJBZHv6Wo/MRlSqo1Vt9YKjXa3J3FlPsm4XO8Pi+xxglXJsVkJUKoVWKYxLMuDF
LRQCTCxKG9dtFdMmJ+X8do3tiZcVpNsXI8nDCPu4CCraPBLCrIEKrh3wsyywz4Eq
UyToDDq5kYz2Gym3y7C1EGwneSFY3Q6/224DVGPbdvb0IVMTC/J4b3Gbc2BcQPaC
D5NW/H2C5hV2EK6q5XhQo2k0lg875iTwr/sPCHL2cVL0CyOjDJZ44bXB6FUd37SW
RcFH2pZP0DM01sIbUA4bYlagcMMLzSU8kH5TmMspjoh2fAIdF0550v6DDKuhn6tt
ahZ2PYDNVMjN6oODbxKyffBT+g5pYBUM3ECsv5xVT6K7e19ikaeeV7let8qhpQZW
vZJqccfkJAdowQ2YQ/d1C/HjCmUADbeAPC4x+TzQFH4f7cFECXMCLZe6QkxbMlHR
YwsFhZ8elZx2CJ2NUJ4vuqaGtRWR8WB47xbOBWTSi2Co79xZAX01TUzp1uxznP8D
iQBqHn3zxbQBU4V+i+7M7v7kRDT45l2MdteAvmxSo0FeDQRZ+YSx7swfyBjXSoNI
3M8L4R+5/P1h9nWKY3lgYR8zF5KUPOpjwVFvY36akSQOSjvNguFyypx8vb1HguWh
YZDnJIqh1ZzqoBlSfsZIhG19Rk57Q1O9Wk6IyQg1f4GN4CHyObyN+hyvA8vmQqbD
1lU+8GN712hSir343pIwdVO1j4PWreYpZ3hyLmWES6yYGkEv/hgjA8st6rolYgFX
YJ1+S/hCQMKh1ygWQ1SLQpKzCogbreDdcTJbTxYbek/5VAZs6YngKMALzrN02LZy
EJz+ySk1SnKCHkJ0SsBidX9/15KyoviqHnkCgDvfmCscbA4mkJLg4q02zVF4GjIv
TRx/ZUEYc8C054BaA4P8BJYnWHxl1Lddjh18jCXJ+9YjQDK1V0UCZVgJHGSuMM6y
yFxcxsgCvQ4oOrBk/Dqkzi1jPy2Ol77wLxKB4YOzwyyUJ7qh84t22pg6+SYd7OI2
dbMqKq9u6o7olQU4iHNYWcy5ZToLyxS6dAon46kgyQcEM9x72+DWUZgmhCuPOgUJ
3SQY15RT6DhH1clSg+/nClHuzGub+xjfpPLfAwZOPzq/t5GO5oYt9IbZ+8U7Y0qo
h3GBtiGHGnzAUl3A6BAMnrF+8g45eKevOOnl8WsrVH++w0iDvzKIy/CwK05b9Pcy
VVjPNKboGT/ZKHjEt5nRzQUY5owHdCr5NhJO233wyC7rDSkfLV89iy1iPHoI4h8t
wwpvin4DrLllpIB6mWGO6ecfywV25M887Ysdn1eiWsYcPTMSzr6Nj0kURpzQUtfb
Hg3bzWOB+rTqTNDA+/ywlsAiQ/0DGYGb4P5TGquQkPweR7k/UZ0vrmwn28Ratoyk
bR0RpCr5Wy8TqzrBaJZT9E0mUomMPBMYcRUFI89ph37eiyBksNJR9hR8swgj0tdL
52nYsj1PoQxyuw/Enw8nirUSmJ3I6jSKTYMyyzF8wmhZzOkfBh5TpfZPQWTV82lR
yLh2EyRfb6XsUbNFYBsZynLBGGj5mryNQ03KlZJaDc2zfL0ft842IaP2H00qsL3K
1SsYvxUdiQVIBB8roaZgtkEJmG+4l/9KJhApvG2838sWmd/tSliNjwnKRxbqJGlx
8sIKX0SKqDj31AhnO4w/LuxhcNfe97qP7+ztWmrq/NGNzY8t6aHFGM4iQh7l1I7K
vchhCxw6lEMu84KiQmkGIMomBF+NMbTctNJVn8WnQB4pA9dFeYd3N3/1Ew9MuV0k
8htkPFP2Ukk7KiN6rvV/B9Kn6OUrlYPVhVg9OgODQqMqGUELbL45xfs7I7xrMGHD
tuYG8AP7fsG9stNpB7nuUBCJe4GRI+kAKQmM/Ay0BcG2DJXzGoJN/E0zbItr9+EJ
2UYQEFg/V/EJANJYAY0XPmji+tVItfYrO/FECoZbG5su+/6/cWu6UnDdGZ2WM4N2
7j/JLT32SVJvqfnkhbP+jFBNPUZcmbkcLIvl/HQRIAHlARq3LsKBt7zWWky1g8D7
4+kQLgXTUD7BFhyed7ZIl1hd6jdozyoCO6xvcLFyofJbjSndltQ5bt91s0sR9gfA
xq8+dFVKS9kPOp9JtiiVMX1VBFSTex+Jv/P7zvVISIYDs2cApJ0oAbb+octucyGg
2+l9TkkIOG9pyj8E+VS2EarLZG5+i13rX19xV6LmFj+pTTDWf89rumdNhO2eL8eg
7DKDYqBBzWaRyAwmYVUZ4ajI/m9GOq3HvqWgunjmcpw2pteFWE+jooBX9492KxJu
ULjHBnNEFKZ4gEeyZsnR+HzOFY7Ib1Lh2VWiyoL3pUCwxF50GT/BBsvvDjwlp6av
FfuC7u/hQt3Mtf0G7dVbH4rn5y6JpGgtcMcTLTsJXXqum3KtzztHY5HT5bXi/KdN
IRjaCGbdtdiYO408iAUVCThRG++ylMDG9tYiepB5Cm6zVUiRb3x+QPQ3GtfPWgNu
0+3Can/5RFk2F2hkKFkm4sA3tXDCq+SOALshY17u/0Ic1yJTCfh7gKHl1tYieiSY
1XOJBTdLUE+UiGmBPQCAScCwjUSQPDeNF1cWd6o++dK3hvjDyJ6ZX/hl4+Go/vkg
N44c8T6YM6YXKAJvuEeLWMCvtXxoYU3V9SUZJfYvm4slEplierMiNsHab6GBsaoA
cmW6S7/aQCcGN3DBGHlTt3opE5oi3trYxpOOWJTLLuizDFQx/v0mYqAZFHyR8BKR
jz6YOuPSSZQt9uPWfnFeD2vUFmSFw0n76mmoIKjSxpvgni6EIIvB2kIgUYMMGBTv
mRJNVcO7nzUEYgyLdSxr2sZezfkDP0IrsZ/V95YkRgWiDbARjh7IboPK4NNxG5ZF
W3HBNxYoUCpjlnK/gItBbfU6cOMBjaHEwz12p+D4vh6l0dICZU7/xkLQpsgHlcXp
39fEqXxxraOx6Q2YJXyfdbZgFoscibIEEjBZ8/ULs8BKPFuW9hvX3iHlAxBV883Z
A7uwbM7cWdC1fETY8xBFwdUk+zeGMd3I7m92In70LH4SDB9l/60ieyzX4vCgs3Hw
/sSeqLywcxxMDzZp/eKsWXUMTwW0uS5b/n0HsXhMDLcXkL9AwZrLCX0kQe94wnU9
ftwa6rJa84itpsfgJ4gw7pvbt0Vw5okJ1bhmMi8pAgaLu7ZqNYJPhwsXtDJ/cnLd
UjXvipolFmBngoxldeuoJdXxZ6pZ5bvaNZIHCKwC3AR+P7wEtPdsinE/vcHAaU+G
YV6JVUXmqD0mXT70F+wO7oxdHKtGfBh5zKSa0EHDYsz/mKqkm0biOOpKcFicL3dG
2L6ppACCLIg/GgmtnzJ5vw7kuuN+eOPgwoKVtojcWvv2Bf0JSM0tw/dZTdWHcS6z
MK+tdATgPkzK6zbwkb46ykTurfgNrW31tiI93D4cr6xintOgxqfg/TNq6ste0AO8
v50PLcbkgIShRfNsgta+CEzteDoHn2mJwFhG3UUzy2IuY1uLc2mP6SCzdJSB6d/R
AVOE1VPPCVuWAQ7yMdZX0GPNitRa81TPEyp8P3M1lSl7fw0IxkUj6YHngoXtWCks
2yamR52DjrVY/ftavSALmLfsT++W/D5zwfx1reIuBia8EKwj4z+okXSJPPLzf9iJ
4MA4Wa1E90E7eLeycgGdBEWyNnqmlDigFbNH4EDM5o3CPDVdqPU5lXrpYLfpRoS/
Hzc98JfWQagVW9jkEs+jEtsdUy1XAl/l7TWAkRMP8EWN+vryug/GZxfTqkQRVvYD
+CFYzeJkNZ6uzJ4gmXOZWlrNvipVgcYqtW4/Wlw4rolVKIcPnNsI707/xLTV2ryR
pQXBPtPZ48NCbWEIAbDdYD2oguSVy03B1A/pCP14Z0bDagyzOppUT7EjhdhhgPwZ
a05a9oVCv15jkTXc+sqfQ3K/uhB1TGNNNfnTvvQR39hwuXOo21piTSJQ3taNGSCu
6yXlC12hnhCDtZ/dpR2I94Irc15Uu9F0zrWo5bTtRG6Puf7fJ5ZTGXY+8GjhB8o1
Q2wVVnZHU2nVx1s8UayHUelMXEaMpA0ORWhVYnIzDcwxybFsx/vKwEH742feKB6d
lFq4G1xBjEriGER5ClHA8ohE0FNED7ZxnXY0aU84wt1Rx98UtKXaeVbxIGObyQyl
g2vBGF+4RHKZNt5PjkGr+L3GXCEh1AaKM42t0j8ufIhZOmLOLcArrVKpwOY3MfD0
vK4rWvP3nuIhINWu+tOCXdetTPN9qzt0dyHdMul6ARP7lvyobruJWXZm0Wof5d1n
n1cfSGDa8FOWTXaulGUuW/pzNjPrwuPCfXIgxlWdkM8ZPoiTekWhk4x82jv36YyX
651CblZYwJPMZqmF0Y5Barq1+QwcSnxZDChvv1M/E4tuv5MBJuUh5hYOUtc1x4fr
uaaYNJJFUY9MOidfM4nKylFRyd8Vbd7fW1JdRLhv+O/CHtwYyim8eCmU1erjBxFD
wwf0oMYw7G3LpKzPwfXvgcyDnp8SAnLBsEtGiNqpdq3TJ7FwtIDGz/YBs84+MXhS
vo8EuHbln/4UvXqT6OUmPQSXYKYIiYFqReQSYpXWgXC8qqJVdcu/+Y5bGbbjjWii
80cWHXO/66U25+pATpnZqjFF5p9pJ4cpFn4hz3VUeq1zlzlHMBzpH5AUXVgv9Uk4
R8rGl3vFYGAuYhitYqASpLSN+1RhMnt39W7O0E7+kommbckEhosFH7mgb/PIKaHy
sLCps3lTFl4JbM1606/lkHs2Py7XVH6TaQnFWY/7qk7F22/u866JWRP5BOzXEvxI
3dl+humvDOUA9jFqD7IIwFNOVXlS3H0BjzEzJulIPTFprJxOFxK/1xOld/96Gy4m
AZr8ZglgojjZLsuKayh1x6KT+HFRSnwJozIx9XW9NVEzAVd0L8RNn5oZ2KnIpgCO
/Do/zN+psRbJXg4jLOBPyqqkOCwDTdqQfJ8V/YzTw1D494jVhkpyg2MxvmMd0Edy
qGDqmZhGPyD+R2fz0oF2pTPDUnAU1CsMaiNCana605FV0msftHxv6W+2Ci/vTswp
CUePQQiiuut80IJoNUIO6f4EfWPT2IPknNzPUi/fEwO+X3ti1Q5sRDtPN47pkMIn
mHI58c+1BF5jgLiVx8yGfbiCw0Rnf2+Xacr8ZvWfg0mHLrwtZNxJT5yGn7u35Uyb
Cn4gWK+ztyO4yFmmLjiOV0i1+x/JXkKpjfVCcegSkuZ0U+fsupnc4pSRfhYuAQJb
PuHYxPVCBK1i6P3oFSPHwIB52n6GEqKxCXKkTyFLKTSbVVKsXksu/fDatksBYY5F
3SGa88+1bRRCxTs9UkU6IIkB/iD0DN3x+WDIgrguF8p+Ftvq97ff+wy0UjebQnHO
Ol1t3G7XnGizoSUWD//b381aWTW7XlI/PaEW6uI0UYYo6N/OzIhmu+y4+qv5nlY7
cH8arT6r3CuU9FpH8oI7rQviJvJ7J2kw14nQjpnT3G+8CSEbgj8MysvhHpHsh58H
9AioWMNMhWpuQ4IifTQ1YB7rXVPcsg2Dz+PCQn29qRP+NIcJivXfM2IwEzGG1k/i
t+hy3almyC3tO+YVn6c6554aEADqYXx+mqr70wBeeJTkQt2YQL4fiUaP2qojhq1Q
uWq5BabdqNAKI8TpcRzTb+9tZHbzkuvcjZTy04vyqNuhmCpM5uGvZ6wts3i9N8Ba
jemCjxUmCeKV5HDNn3oQgrMSXY6Gy875rPramkXSIbLnq6O1vNASJpQfPNMSPZGM
5PWU+Ii/284BdKL22PBa0pPTlynTfuuxAHkWGh1syB2d1DSYfWs9t32+iankFX/9
x/phzKpFHnMIaa5m4grpNE0fRM0XCFvJ75C/51+N2e7zdr26HwewDnOwf7SpXDxz
XviWjo30UutKjWCjWj4NXhJZRRzIpLkhlibewT2KtDPkdMyhAstWSoTSa8bSxS1k
QBrj0q3gBtye61VJzo+96d+cCAd3g754Qa6O8UgLeWONpZY3VtOkAiJu1LT7ekE/
eoqgjo0tX58T81gAWyix41gcuSPwSgMorivGnz9I4a9G9UqJQEkPJmZ2nfzRLog4
bmu2B3Sbutx3Gt0iHBmWIVPkc77yexToWldlInxdCQoPjV/h3qh8a1b/vnFnwjsB
5x2qqk33R0agaOlh5NcPAoEOz1o1X0ETUdLD3A7IbBlk1iH20v4KjZmIJOGijMtW
Hr8A8LnOJ7mdX6iSwi/3sTzrxXuPC9mMg517xyBNWp2u2jb+KqBS/G1gUUFwH71i
wUI1uTg09QDlMuFluGxVXXkkYyqOemkMOckW/ancgt0Yb+T6kn3yUsZtr1HvyOyX
FbjMiYyeoiPyr5wjdOFnNQuW9ZEZuc2YLEoYpvDPwRn2DBM+fNpMmKVD/kmtUjVd
RCHXSlGnytRzztO7jWC5pu3EcIuvCF2yNG0o8BBL9blkRGk6JbE2a5IqpjduGlZL
hZvcOr0Mj4vYYRST17Uf05LM91fUj4UEj1fKrGwNubdNTvSAaVGLUij3OONbKt1J
lJBkvX0C6aAPJgx6XCt/iKqbFJrNLSiOmQRSuIucdq2ZKRdXWmRWLluP+I93vPmt
4nMmgBoNvb1jWubj7KKPxVv2qvhpd2vaSqCk/6b6S53Wa7eBjDjmBJq3JuXz4XYA
38Cg8nWx4lftJF0xWjYoJmmXavofzTAGD9KSmet+xMrarIFpGDUddQ1+ylYny4Dj
wJu2Sh+CU6apTJK9oamNJEws1DHWUZiYsca3vGHdimvWHN3yIxZO7eSGLsTZNXCw
FnhboDkDaMFXnKBmg2JBhZGWFTTJIS0D1mfm1vfNZBwxaveyhrmLokW+ZAFNt89r
0Ij8Gwq2W6ApdrcbUoSokZ0Mz17i3r8rBYtexpjsp6bYBnKhV3rROCTgrLIQ5NNa
Ss7GatH9QGfSyrpaU5kDBIqKGlK5/wmmZnOlcMiHCemQFXD8NCopglx9X4uxl3VS
dXrggVv4n/VimwOACvwPaWXW2mRInYsT8OB99/edS7MiBtmCIi+Z6SFWh2/q8D6s
C0ca3ixH7MhsGCvBpTLbRmvbI0XFXaZz3uG8GimSUEsfcqDxijXCa3KtO201eldM
I09gJFm8v52TyVmlBdCWPCsgMbRsOVF5XnyQk/gdSMqqBqy5koqSA82tM79E9ZgC
w4e83sXSwQ87CyjJz6uW5NTPUgKxAZvnimHiJLv9+dt7yuiwE56zfy9DKumko4Ok
TILcP2sqFreV32+lYNgRBaDD6smqh/TYPSaAdd7yPMrtHm7FgzyKRe+/i+5pOAOo
k58281Vd50CPSN6buvHaFbtirdqGaxW/1hiWTYChckxWbOMKtaM+VHg8wm8c/jGW
qgboMRR2POHQOKJIN/KUn43tEpuegrrpAILMFg/fwDDQDxW4Jpbp9Ms5awKNMyqJ
97lnVgqhLhQkLzOXwfwCPK6e2N2Akqu7bUkQiVS/jH+BTR3xaV3bYJnOPwx65090
pO2I8XTg3Xo7MkCtk/W+ui0tWMk9f08qSr9czfDwPgPyI6+jsJ3Z4uEHIf8TStGw
wFgg/tis+CcM0eMJIq/wI4e9w2Bc4g9ZvgPb4Xlswu315DdNBjoevAdELz2f3ZYE
HE2501Hctcva/jbHUBMbPYd4TApLUvF1uCjo6bW3RPyIDtMi2/rpxczyGwPh9zk/
PCxO0+Ayh9Q4TrF+E7MgcSCAOI6RilMt+/iNjoEOzJ0Fd7bgQu9K2pwNfU64f9SN
L7wOy54Vu4GwfxseZgNCm3ctFcT+psdClwxgkGuQLe/94xL4i8LxYxLDRxv/DRu1
NBWWSHaE/dKlgR/WTcv1SP2hnFf49jwWhPjhAU4SSDIzuQjWbI/V1CEleSMaQgVH
BMbqVMreRtOMhzS74g+R1F/yQUQXK8ccpeKuephogwJenE+GSw4+K67oEc1VKV2P
vzMCSKtpjPGBLTessrWuWssVcaddnoNlbsEAk0FawPy4K65fhlIt1gcQE5SKkrsM
Q47CQdD3rmsTXD1yQX/QiJe9/LDqwcaGY2I64+wrUVbWs4FIWPYdU19cawwno+oh
JFJ7zMDGca3WWUAIDLsztYKtWiADWMgpPqLYOtXvEhLA58I0b++Dxq+1B18kaeQy
k/VoWGFh4MBypk3ACMdYmYMxu9tYJnQnU/C6u41LLVRo/kP6mH+Mrat1Qm2+U5iM
SJ6nTZX35pkF3OPBufHYNBYFEerYIiWtL6ZuRhATTGuXsYAmiMJkPhg4djOUzdpp
3Ow1mNOO2G8RMhOB9Zux7xJqTkMz87d0K4DdHNkq8BX+odf5sq0plRB2pnO0Ikgv
x9bH3ogqjcstf8ypb1lOIA3/4cQHy2EmyU+MKq+YD54qpgRkmfdzIKA6Ze+vOLhk
EI/Bgitk2rql48tMQGhMEs2nlvSXW8N9CE+3CRm79m3TE5Bk6LfbYm+DngpR2VLI
07lO+VftJhx1XS8mmJZ3CKTZxxBuiqw5WgxWfI72YCGDgJYln6OaqHkxRCDj43tp
FVoisHhqk9dUDopMHbtiZzQLk4laCJYNU6AJNxzIxLzt4kdjfOoaxFGkPsda8Hay
jdVM/wUv1DOO64hUP6mZOyrS6yGpk1RMTwoRg/ebt7P6TBJu/6T+KsobKKjf2Mwg
Mj7Wsiw91WMzHK7QqLagyM1qOn2JsT3LkLr9F4U23AQcl9tLb5D9pNmeV3RHSOiM
3Nm3c5nrrl2TVYgo9n7rGzw4bRVzrdcK5HhuDcYLQ1IYM2eMEUjxy9mpVtcBsLmH
EuS7ZMZj6Qjf6I6LfNUCkcFcCTF4QErYmX8cwIbEUvy1sveEZPVMqjL1vZI1/yzL
5ftK3qpL1GLT4azzJn12tTbqYLGmQiA90Sk591ko5lROldSUewFq80O8uik34Pxd
oGW4RZ1l8TOqZz5UIJVNzW/e++PsfEGxWmgm+23TSHHY+87sUNjAVfmKx7zvcD9I
wUHjx4yc9cdVvx1WoBM8+7TqONYgU3M3ClBXX73zqwAJh7vXIOk51U35s6jtXyaj
0UKGaoy3l1qKH+MTWUBfzEG/dvoZFXcYLcEvXz5QKiT90W1E7HKMMbPrBAHTrveR
vHEMkqwhQno2Z87UqnZB2BF19dP033v73KmFwRScqJm8T4+VuWGGV5S6H1jvJtwV
0yzSMyCzhW7o33nclzDYIAOdIbnhGiMrmV2VedvqlJYK4tqzM4xIkYJxkpRUk9sL
XzHpIh/lkhqn/CR49e9iKwSg+Vu2An3532tT1+U67j2iC7yjY8LA6erQ5UWWD91k
jahUirwtMtx1iooQ7lkqJi4YUweI5mNynEtl2D2caRQn2dTggN0oEsI5QAIUosHg
tlNI9XCKhwIYyJhpi7gZtEKZ9qRXWaJVIob5idmGT3NWAdJksV/UUmZCwAaJNCt5
Uny6dqzV7G4syQIsdC+YJ1R91qpJ6Meg5xjmebtMPVzQa5IwNjMSbQJOaHDpAu2c
dXYPuL4YzPPGtcK2NshsooQm/e+LCDDItt8/ZtZAH9NE3S+yot8/6dgYu7IeGtaC
d23qLd5ibKSi8JIqNmoSQz759zRdbzM47hCLvRCb3CsZ/O7Gd/QrEwLZ+qXawoKm
0RkLlgF87B3EtLQiyLePtZzB3Hi2x0SsxkA+u18sz4cYty1lJzR8sTRnkLzhptHD
m4FSc4DOp6XMMCVDOFKEJj9bISKGDqbBBi18/EgktuMTTNlWNWgIgcuvdah+cvx0
1vEFRKuPOyzpuR38B1bWHggG2xg4CxzGpRMu1HrJQG9Ps0SaQqeyLt3HwZFyJpot
7dp1McfECM+A2JMQIaiKir+63YSdeQmh4qaCnymdkNycJnzwkQuIMSoLHm6CvtMV
DZ9DQKgHp8qGojz3gZJPYdF8ozb4mvBzUjFKSY7HxvoTF6Q8kwRRPwgit/cU1lln
jOXbZHjPc5UQ8q3vo3yLYpi/lJo64VcYRdZdDpkTt8o3j4J9L+MaFUrdOD28UM+W
JrVL8njnRcmVi+TWfXyZiohEnwaXj76jzXc2GAnCglJK9KHPORT20uyWMGz8QGBn
fwc/8U9d4tgjIKxzv6Iz/Klk3kG3nh7NA4kLaapBFXkxI1JEtsX4MLgoJoGwi4o4
ACU5A5/r6+hANHVFfBIlx1tIkxTJyALCI3MKiq6SpAyov2i8sKCzfUBYceMNs80A
pvFFXjbh+Coo2z0b36Z3ltzjOV5QnQYwGf866AYowiExf7fMMFKjMXk6+KQmHJ0D
E7IMX+yzDz53St0BUMv8VEBy/4yCQVzht9oWy7CqrrsplvWINowOcEHsn6a8Wjb1
PgfVw+xq2yxvEMiAn3iSLOXLqWJGPCrQ402eePnvLCA649r0hpkhgoezZ19/hAx9
7AkJyHE671d27J9qknRRKD1KsLh9msIIkhTaLaRgrzgKtsDgtisZjnDngpa72jNu
u80suiLZlNrLmR540TIMYKGYWkaEEAaWm22O24ZAJLP2bATK0bacskmwislDPpPs
FXMnRMlmWeYlHnZSABGy0Nf5Vz4aCnZbfc94d4eyqifXoTOIogtoJHkr9LkSSgR5
8Ht/e25u1CtCrIvwPyeBFpVofCRCBO45eIvsGmrjR8v22VP0pQzRZbSqJ5L+n/4d
jEJd0mRNb5QrO+JYC0iNLJR3U8nuQcGq3bty76lZLmBPsLRootvWOo/pCiTP3RBy
rD+7kqvyCAGGUDw48jYFmW341zGv1QfusYC77Bwh8SbPVrC7VGJTkMc+e2ywX/y+
pVjtLvjIyOPN8xTZ712CZxd58s6DGw3392nzzI1uuREolnnJeEk4hnxU/P2+X92i
9yNytA2XHZUA8G0fTyRZP3xoUbhSSd+RaJ0DFjEly1kBWN9Uk1pRhXxTyi6//H2J
IaHcPczkF6nAjd3fKahO7m8gKCHXivKE9aZvap5cFWz1kQNwfDONVnIGWrzyD+DL
9xbJ5D1qLOVr0eTYJzpa/lUKy1veZ4reHcgl3ztvrEjFJBFmpv2pJGFJKnaub3w8
MpEnyQIk3fmtnvCYG8WE6Cojg6/wuFFgmIhZXmqP6QTMqKsnR65ZGR4iaMFjiX3N
4lAd7D/6Qa6RcJ/seGJHhg3wSgssN6+Sd6PYruv5RSZ+7BWUS1buvfkBXDhsrYud
LHvdlqBFTNfedMsi+9c7uMmoaaZKf+rJd0WlLUvyf/W1ycSHZPWreFFB+K/rQSFP
7cSlGBUIOkfN/pbDyxJ59U3t94WLbG0Ww9eZI2keF+DJHi5p2+/QjWqS4jy2tEH3
AU6vo5VZWw65iGEiYvPvrGg0TLLN5N6QdPvK8g5txfnlzYTlTjnxfRW+G6uCB7q+
XZHrPBALgAe1/Bwr8gm4mzS5btydhDZeaIn8qp8y1/KVijJnsA/NVp5dy+cl0J5j
7iD12zkDBgYYS/XTveM4cevFWuxO8gYL2IqyVZfWQHjuK7wOEaLtvjpfcKL8bVsd
vAgmF8zsDVikuDNX5Hus+tSmVYG/fSl9JGA6ULOjAy1FgNdH1MhMEkquZswnSPSs
hIlqzZFySQsES/u5931fYkGLVGXUan4C6EA5PIX53sYPR2pmQeKmvddjRGD4oIt5
bZATtjdy7h0i77QuxZJCWIlNSD8L/ois0xW53xPx+9JF6lfdykbOjEndQdnJRZaz
6j9jCG+zCyaFLb4dyDgDt04mV3UcdhtKxcG0gvjVrfGRpAfq6ctCWO4Bw5Tyx9mW
IhqoMB09Xq2He/MwAt9YNY0AV4ZpQeuhYKszJ8OZBwHOgK5Mqdz5U3rLWlVkWhG2
kNQ7oCwXg+9Gra8k6ME0JL4COZazU7YgGrXN+TPloS9l1D3sNA31zUuLIVdpBguX
ITYBMt9CpZu8WdvDbZVW5xPg3F3f28a5LYfuOxBIS2AlKLEXSvvJU/+HTDXR5Jno
5cA29raZ5fP8fx1nHz+CQvG3witlfLdRvMtG3AYrr+DeIw3OowEithD1pd/eHPID
aosgHjxcu0u0XTfhA46wqxdqbCQrsZUEgltwS1+JPLx7nS/Zteix1EM5SVKlR9yb
HbTUSKAdN/+PDwU41fteChkSBbi8HtRNp4AlwFmFdlg4ny17tUOsXfTPL3Kta/tA
aM3a4KnNOPnkJkN0JbgY2gGtYS01B7KbfhfI0JGSvMCBrh54TadS7C/Dhuh5WPTr
jcTuGuRUDC70+A4wkx6W+j+7XDqHEcllxjsGVLqLwCK4fOO/IlXX07HYx/5onquG
mGXVSIUCo5euYOgWNz5UHnrgj0geIILHtrWapp3G3u8ojtpP6KXTtFiaJ5n1J7HE
yrsIbRHN5BblHpSl9CNaRdRwYFssE3Tgpop5wMmzKnAcykYU8wohDetIFFrIYGT1
iUDLOVEPqyOluqXwFZWNgNW9WJH+7UaWN7XZP3pne7KPyk8cJlojVwW7SX52FcMj
zMBju8ZmRmgw3RiTYCuwk4q4tgJ0qjOGjbPgL/OC35huYo2BTAruS578afOhEcQ0
+fHvZO9WR2x+6zFKJzMrmbRo+hQJoPx3sj+WX5GcoEeZYwBOAu5TdqMFw3dsFSrJ
ExepDURx+tcBWmitg/ZGcPtU9lLTMYK0oTlnQKW8+MRKTh6Po+kAnXGmvFC6w1l8
jIJPo8oVvbMOwCTbN7il/5u3ADZAgagPEhrjoKbeAancNuSaxbZfNZIalZS1dlDM
Nc0gCCla+IO+1NlIqVyrqZqkNIlu5A6y+4FBOJXZjNNDDCFj673/TdqGaF1YRpuK
LIsZ+Q7jooC26r9EnLX2XDFq80kQrtReXUiRFEsBniTggK7LIHRfynNAFAjlo1Yk
3s445W5XxJtH3N73zsAyhEOWzKqBtdxshXStiXzmNdlUz6l95Sr9FeLuOhIdep4M
6Gw0Rmk6btJLKf4I1DFDboK4/8E0loJ+pgx5C59Z14dFsS+THWLzEukqbQFAqql5
G5+rr+AHsTT0VKctDOiRVUy4YZzbblIVnNniByltxYTRvedzdgPE9N7WmWiyo1Uk
53435JPuXVNPiyviK90BiCqBe+UDe0f9ocb7n/mp33tozYX+YTVenn1YK0yb2HZa
SJ0euX+cFEMbi2PYCem26ApGcEGrViPv8D35BJAXqEba2Ynp4u8bPiH3QHVt3nLd
0Vsi8W2a1QgaTBBMAUATs+mSNk0tIwymr1trgc2jGjrKWizK/VO2v41QGNYNLkp0
zVczXfLi+Al/XrvhkOkHZ713T0hYBAtyRiwoTUfBeXbTwU/iI3Gcscyagb3PZqgM
56iTtiuiVsNSMFHtP5paXe8P/ryRkIhryyhgzYr0UZ81TeVcdAeSz3AUmG4kRJ53
kucEcYdy4AjT6fCBGdXUfxoZRYrhGL01h1jYcU29vUSgmi6wduKBnO5boTH2XvRY
UH3Qjus4FLzD5NoVedo2sJtyONk0VRcm2wRgT/M8WYNroCd/E6eQBWkm2OoDnWET
wnKJwEnVgcvmgJ22hIoRixbT9dZm+W0XJqc0meztb5CtkPSQLzt7lLXm0Z9ZRpm5
n7/3BxeTcj2xK1MOtyrO1JshKKR8812z/FTe/vllz08zJqkOxbkYZSex1Fhu76ke
nx/PKEEDYIYtr8BbhUouacCdG3xOszjLn4iTsn/UvhMQBT6EQYjs57KjycwAkIUn
vVTFbkCfo81qqiWSRlQZ/9XEBJcqhyluLtDCaJAb7pKHeHfmCHfDKL4vxUSMZHz1
2Njv4089YcsHYXE4yYQYdeMIqxMoMocuteXC45e6Z8plNzzhocX96v4lOW68M2wj
3/rZfjsNNXqdRWTbGu0IFCO7H07oiCrJzF00wwfFbh9NxFcHmrKFsBmP70Vs5Nrp
asZGSrqMQKBchXuWpJI/zKVswgP07turKMwHVu1S4Z6lT0M/UO3bmyvjaoN0wQPi
+dpgyfGsaIXnTE2pcGWhaZIl4CrUbdut/V75BdTb84FwISAloFvBWsEwT4FfC6mW
34AthqWJ0AO0o8xv8pr3kcPM7Fl9aUr6vz6lxM3uNajVOGjpbI6zTY5fk6duGx/6
AXewMnNvSUEKdOG+bHrPipDShH0OqK0w295IDtYcBeg9NOkaV3XUcFws8Ar8twGb
HMxcDcdTGvRkx7fnb5nzoerEdoNYCOhKV6tR3th8CtItfUgtQRxeczbyHRDWMFdM
2j70nSzhX5O9dZd6qPSm5tyVilCjD9I5cCWkIl1MpzB4IUQU7zSPH2EGsCrPTaFb
GQ+yg9pAMt17L+MX+DQ+zytvE95ywG/NXvjOGgzk9k4+8McGcG0/WkNEmf+81rN9
DE5vohQ7qx4ObfSMcMa2dqfZyqFQiwvGxXJiAHWiePkGRHhjv8QHxeDMDpQwOx7Y
pwzg6wBetAO83Bep1V7UlgFwdqJ+0ESIxIqvSjlNkOsda9tyAgDKRJvKsb6dFXRB
0TbAMea8hgGnzdzIA9VWDuqgy9+OJj6oGDWPTVWkSRZHkbF6YhAID4iXIfUODXuW
BS07WadYQhBHGAwSMnUi35vWQ4AR2kSJ0UKM7cZ7FPT78t10P61a+bZ9lVvixcKt
mGeiARfFE3nSvcIwFETHnLHLQTejA124sK5iLRoftqitTkJ9n5GtFCB88j9pZgA3
Qle1TXMuuNji8aXRjLUFV9m3YUKHur4IHPCb/J80EgJs/BZAoTHxWBiYRum35rkq
ihiYni1rLQG5/ROr55438uoWJkhv4rrnabJbpF0cvcO1fY0FcZC/NbY+vP4nn60T
UHMMNk2kJSeaI9VgcCSYm5mD9M5Q2f6/VEsa9B5Rr3hpj276syTDNyRyU/bOH99z
fPEsCEgCCEKD1KagML0/m8TezB6YG8iuaGP7vulV3yD926cQOYmjOTiLjypAbkcd
ngBkLSWG+JlQp8fRmCQCatk0I7G/WZ+Sx0LvThF5DTPtF7A+2K6/xBMJtdoxR8yD
g3vPV+CJNyVEgwGnSFz1z8j3F5PmZS/zs+5rUwh37x22jKQXVRkVnmn1lr+h4Cqq
5VdbBStq3+e0iLlyJdQDiE5L6QZ6caRwmDORJwxAIjAFLAn6dpv0yt0EsDAXZx/P
eud2hGKbnUZpruUlXvwM24KGinpChWcprxuu0GgScuCmaqEJwtszPsRSMSyzpNnS
1FcEn+LQXvfW/+3eNajKQgySEI/8MKwxqiAOLcv6J1PB5AM87j2lDQvM+tn6u85Q
iT3LZILd1sCgozMMdrqTtZO7XCwLCTfZ017udNrudk+U9wy/dw0lKKLO6LBgx6Hl
Sw41BfZzvcqJzKRgoTIxHC6GDSANQdAmo7tr6zOekYfPXjnfy9F+1ewThxg8wUCf
MJgiZ0OdCgPF5rNGZQhKS6bndV3mayWUKwaLb3iL8GXydGd0pz4eJJDW1yYQajvM
gZRG4nHcV3NKMUTwbcgbBsGU3AgJyV/Y2wDg+5mt7ARFwWDQEXMoNMr+Z703V4A+
vtE70z4/RWCqjkXI4PnaQnUXwUgoD8hpecaqIdGoej99mmrEQBs2w75TqE7Tz1MO
/hQq4O+fz10tVBOGk/UVw3UgzkgWylSGQHEQJPFTwRT0ENcuSHbEQmywiR0Nze3G
paCqIuoBEOKbBw4IS2vh0iouEf7iTtUC46IY/b0+7mVjIscuDwYZLs3ywsueuQaz
XdM4Bs1K+erhrqP9RnNsQ/Ml8HyJvSIVCIOEKrgkCWJelxqPo37OVmGEQl6J46qb
ndZzixLVFniSfRArAr6YiKqb9Ae8/qOOso5QmRo3MhyUGFdb/Pew8+le/E6SeFGm
sWPBLpZCBEH1h1ONiyOIGR6S1zc63+9L99Wwte1+RjLMqlp8EoHk/vnghJ6sapmN
gqKjkagOJ3mkPPR0ex0H9SfriD7tqVfwc0iBtuS/m6V9exb43DwjzJYL95gAFj02
gW76jwnTJ1ZfoK8tK7YuPDNFGYKJOA9SU0uP/XkHXuUttdAeuOUPR2WhrpI6tqaR
8mXc7jrnIjkXanUJjqedlfsmkFvLhQtQTSwHB1pkG/QU6vJ3VsOMXbQWcNJ151MI
X62WHaAk+et5YoNEBAnp4gg7dHXq6VSFXYvKPrexObQr7avgT3VlMRmYdhVVYBqD
ryG4cr9wB/Ov+6IV9xXbm7/WOCed/f7QpGR8FNxkznaaQcSfEV+bfeUCyzh//t8C
ZqhFt/fUkomtdq+nnjDFBSPId6YhYLPfeJkXO/XxkIHmGLO0YvW25YRG/B0hX1nL
BToQM2qU5Ro6KyDA52ASUzCBuLcdX2KsBhnSbksCGlulRgSz1iod8YW4Vjc/+Bvo
t/osHLt0gAhE6G5+F6O1Ize7OnJ08PYAskYefe1Z5xETA6XKwOEMicIYIhndzfCE
OSBf48/Db26HV2wokC99zIp4IQKTxDrz9CZ2FHklYUFmEkSigksue9m0a2xP0g0Y
rpWkrzvlrbRiiQ6DA+P1UIjXUM/8FOnIQ7iUkRDXCAnSHpY6XRrLfXmlaUKeFfo/
+rry916SsRVqRD83wsdyVg7XQ2+CJJmXi3BRfrQtj4bLDKy3R1lFwHIo4M3I0Q86
R6Z9LE2IlCC8b55V51RzUCp01Ibq+I0L6hrWC/LbhPg441dMg5PN/pOrtu+YiJ6l
pn0tq+ci0FLdSF0lMKvbTJnlnLUwSEW9fLb6Doz/YQ0RY5NkXQLPZsuRXfKNYXgx
VBcQ2mCoYfWbSBf+0x2iEY6mK5Eb/blgmRfNF0se1JvqbgVPcy+jZ+rhPKpWu5PU
Jwjx9UTW9MgOhWvj1+OBasEsNetucvJ4CpZOQ07mjG/o7+GrAoUnGzxk5aFCeKxK
jWOv6QpvIFELe2R+H4O8sR6b0acyad/Xe/HkzNiP+OTTDntpNMBnB9jOEsjwMr+e
PrU3/+VGJQHc1Of/R3EUyIeL0Q82n9GTnPEHMtKPb2SxgfoA+UY7XRcA9q5wor6h
S4HEa83xdmG36e92L0rcZpN5toeM6Nhzp7JqNvMi6WC8YIPLqwEzrHaHvOj2rDip
C4dCXs6PFB4A1E3Ewn0jzJXcs5Glk9EooB0HrKM7ggMY/IFmsW7mF3DmOXGI370N
oOA/asqJciquR0jFJkU1cXiaYdiRxJ0VK59ZfVEi7bFspAN7w68DiG0ROGVPbFGa
2kXviGBMcFII4Al2Zs+eQLjRtShR2WuWRhMFWzhilxJyOwm9S+05cvOOAv89/U/B
/m5siWSn2/jslWQriv41asXS9LurWyiKkr5FJDX5Waic34cW54kSt6HdeLizJpFN
OnQgvQHYnsQHQSDS404753gcR04CbGFBhUU1ScXFW+6DfiahQNt7A1+vEqBhtbwH
sO6iPGtMUyPU/48RItpkzZ8gXm426vyO4J2ScQS2AVcAXsz9l5zOk2wu3OkIbXzH
l7LTC0ZQlgU1fDZwsWc7zGguaKqvH3pDhMe2tsa/1+kGOEbC5aqEBfGPRHbWJyLO
OoS1CRF7kvSnDx7aPo95AYFMotV4anW2ObIThic+FchIgu8lYjuGRTvKwzIwS9zB
OrJ6Q3Sq0aXyZZW3zVBMwEiaAUSKXeuecLA6na2fUeAhzWWMGqzU87cfytYcGgxR
Tz/1HGQY08JOhnnhdX6/OjFmk3yYFyap/aKZCSFoS2seHSHNL+eCEvNRUAgGkIiV
vK9kFoWDm5j/CP8xmyGEoUtJMpO0Gas3SEA4xPzPD06Plt3/dlQliZF2JT9HJznt
ie1s7yua367z+PhkT6/T4bBjoWinR+UZ+RSPA0+GWCu0VImNg/lI89zkmSOmDuAO
49TaENoRZUbepi/cltU+hqAWp2yVh0cl9H0UrRUgeDcjuJcz2kQrvDzXTH+RYLOf
S2Q8QACFN0T3Fb7fM2+HWN57XhVjk48ZCowgxOHnBPjHunfT4FhaBabqD8rqwLhb
ml66/d/65WauyTQ1fRFCzusD5UHBPUyik/moZZqMuiskjZeQnsJaNJpdpuO5+97i
XIumpFcrYE6wtMncVOLFVtw9S5MolmBLYbOuR3K/jlDtdj1vS4sAi6tAkpJgipBt
jc0rdB3N63dJAbSphqsKUxtC49SnVK8qStZBrlRhv8JXA4CNHniMZUbXDWlP56OD
raT72FNNB9TB9vIkqdMmJgURJC+Ypcr6VVAwvBD3nKQd0xECQaN8OOEGvM/OevBz
KLN1tYR7+ynjZKERBga6R0e9EAtc7vbIOkIVUR7ARRX2vjYB7fZPTuz00BnSw9Ev
+d/WQ88qR5+aPE1wJKK0pT4D5ss8GhTD2ym2Y5j9vsYYLre8AALCfw/p50qcoutE
mPl12+hVrMXVsNfQuc8OU9p18GqzVRpYh7WmUubDSgccqEmh5yL8o3YEfG/1sFIe
VDwG2ajGolR7r1CAN38+7JHbl/vBZ9nqp/fCdxaeLxl7KW0WCvFnkLOdcimsttya
Q1zWrcmfNInw3dTMCowjQJ16nfD/yp12qU2L540G3W8A+iVAne5LUsZSqhIhu1Ch
ShNiHSgIC9VfivZlPxW8XpSWLy1mzqCRlf/Y6swDV5xIIfUSp+4co8NHUU3uVLvF
BVpq9e02rPGI1kG5eRUIRMs8nj7YPbXHs4jGx7Us+i01jyPfBDDUcxwiAppTeUwU
hBDzIrgubr31SjksN/jSPC0AHa1hHuNV+L2QdPbACh/DdlhLL2vSr8AgWb0vULsW
/8nZd3cNA2E/VgT0rikLLKRBXeOwpTjYgUFmtI7Rs0v6sVX8jdjMDDVebW3IGmzd
xMckBb37Syvm/I25vEszyvQrLMS1dllhKMbrhfVzbPkx/dC9Nsp/1wmKiGaicVt5
ULFSui4TyWdYbav7PtoXnCMpvS2dXT5qSboYV5BZK5Emy/D12Ncie7uwf/1ZvGvv
WkBLSTBOFC3jS0tZ3tRugAsoZ3QgIMkd6PCoMpl/3kg3PPFgGdO3PnrpgBjhA5Zj
DDjOxaDy7ISQaiLw7u0CJRrhHM/eBcK09Btr4barxm7Pclj6JXpSweImYG+hCQ+k
rWjvIncOjTACAYFZK6YmdU5w7hmy6E93jYll2Q7e4n4G4/OFMKDAt79pOTh11ETM
Y/1FjPmVZ3gQkAxpbBbgQiMEY7DklwVAJoYHPCzzgDQY4STIyyyryQKVtOzAVe8T
faHyGomUHRI4oq5gvj7AMEikwzp/y7nR4/1P5byTdenKIX4CNLA1iFWiPf8SQv8x
TrLsZct5UOVBQGBtSD13/f3xVYGsqAYdZuS4xc9yukx90glrJ4XflZmKqYlgzQaH
IAhetqEWst2gMuRvmDEzwl23ys6rYJ1tWM3bobUoI1LaTXZ7/qiH+BKkuxXjyGbd
Gi/qGTyDyyq1xNSi6CxupbkSJA+QAj+Ss1T+AyRPvPHyoegwj/9oMZyxntxLCqhX
sqgnhh3XR7Jl9pljLBm4kfZdhFsMv+2x0u6paiCzxWaaoSOLR85IRi3B/2zyvRPC
ZG4Mo6/ejzj5YPjTHaCCugonLvC1LGcbWGImDM45xs4tTZW0/iwkFMooHnvNnC4I
MTA+Kj1yk/atMK2ZRIOfnNzXMcg6BSVwz/hycR1BB+RKsL/6x/rogLfhe0DXGttO
TKXmE/zAoWWiXFselfGgTDQhZjm6oCbXkOXoChTc+CoXfa3j81p9kW6sFpeDhyld
i5qgC4C6s7eh1gomrxFzkKYyNvsCShNykOJVUgY7+JvePEQk7Fu0sQO8pnj2dJ8g
wwC1Qc8LWScpmyQXmlDy6IhcB3YZuUY/fiaVak9S8H1DmkKMwzL16L18XIi+xZzF
MJlxI40Hx6B39EzvnsM8NF/18Cpn0sEwEhZ2cI3/Z7WXzwEn8kQXI5+Jb8lenBYj
mJocbg5DXLhR+AY297M8g+qHCHdxG+x21LKusN8tOI2Yw1wnX3Jg94TeoyoUEnW3
Vkq2g6Gl9F2Hg6Qjoa/D+nGzhKuPcsglhiWDcHqVvocZH3jl+dKhN0X23NqHUaC+
K2hmVbZjZEdiLf6b1zeaXKNjyXA+2rcyUzOo7Nt43NHHkOSsSRG4QDrPw7Kd2fdT
3BB7eK9N7+h3GBEUJiSlubTLZ6RGf6PECanQBm93yuU8s4T11Js8vCEj0eH1bUzf
/AB/IDrHZzAr8ItHC+YwPIe4l30V2HBaR+/eIYmQDeWiExxoZkdR8ou2murnuqxb
bMt3KJ3Cz9pAyH6L+jHhI8tTtm444MMGh4FHMCW3FYdRHDgZnd6fQcNIg8croX7q
CyawbV8d9uNhc7o3llKbTT2jpY/YghYZbS0pfWFxDYQlnSw4fNqY2exj7gU4ln9U
u9WSS3OqIFC0lTBV5jxzbH0NN+Mk0nGh+g+hPJ0ZeP6jnvJ3iLgNge2Av8uxLfFq
h4F7j2foS+NBjXL8yBrMTRH851J1eHSFQPZXcqI3j60rywRGMvYWT0NudKpjggXi
PSn/QcqrSPWB7ZKcMx4gXFOgOGptq5+/01XA0+ixpkZWF6Eyih9akl7iOK7sZq/a
Y6bhFhseLx05DZgovt1kmK4yxeVg5mLNZQqMRSEMwm9+ySZb5cPhboqVO4qn8loR
OZZoHEQ38zwK/72vnxe/GBNMc/GY1k9fbv3zREMkx80/ePuc6oHUeIaH9/OZfYro
LLC3YarfS9Pi62CLJls99OmcEgFljixEjK9yx6geiwcWHh1pFNXLNyPwFjIXD2ZW
h29yRR92RbYjLgh5tspI+ZltYROiqwtMMFU8OueTn6oFbOCutspxg6vgiwfRLeT7
vUBt52opEHo1kjGHhHufECuu04CyAWDXppOVmlwtL7+hWDdLz7HEKbpvcVWIjFO/
jyYMqVbucgHrbdZ+22sssK+ujMQjoLSxMKzLMQ7yEfau97CYSKoGbRlBwt0qdln/
Y9ERxxmFEFpHN4Bb+twQvaJDTLEliHBztHtwg/IRlEdtlayGLJjlaK/X4lNnMmTu
qb3qUizWtznygM6QRLcTu7QnFyT11hxQduZ3w9wEhrtW/3sQ8lWm6swUsrXAms0/
CzsFdekJQdCW8uMqc/3zToPzAX0cc7nvjoJhiwI9G5PP2hdqwpeWlpwb26aBPYhu
PqjcxAhPWLmCp9u1+Quh0IlfreB8AukB/uYLLqKY2pm8O3jVQKnQkEsMHaYRoC+h
sGbFtU8/7N2u6toZBgNttlMU0NRdUb5Ixdo8m4Fx8c/eyDffSXvF+w3C+OmeBFa3
mdbMk2w3QufoYqMVOi/9rr/g3yu7m46w30TrC9+2Guv43XvbZXUPAhogCaf3PVEt
ESl5rJKlokKOYd0QO7u83hsXzsar4MISSm7+ovXgoGYKOCMJLPmaOZTESc6TSJyj
ZnRSuPSfh4cNyf3EjPyLIPrG9+F+DR/PxlggcQrT8H0J0tgb2UUzxRJGEQipFoQ2
k6tjFuWTEcHZR3Yi4IMD7y03DLr+OlbVXtukCbN+5Q/KikxAITiL08rZVaZAZ1SF
csWTO3LCwdyQ5VE1ZlXZm1LSoI/ILER2TIGFFtrQaR/6tB0EVum4rU2LvWPimhdF
IR7kSL3IfeIqOiFwz0XJhzooi5zUzw7sFeU0ZvoslHvltyRLvbrA4IPq7HXDLzDs
6iF1zQ1Zcwe10N+uVSzSspyaws19569+0oZSLFQHKxQ6wiVkCf/mUpxnlEH/AurG
ehU4KR2+Al3LTSJ1DHKjFhYM1BAh9DyrM9+13jq3nV2fRhu/Gl6pH/5LRhEclP4b
gP6e2BitK9I0L79shmpY7fkydAkpx0J0XX+q+BJSa7f/fdV4TE5ku0PKm7Qe4p9p
r/ojH724o+5YBbaOcvYxc+Y/0ukVCK6xYCXMSSm6O8ZUGaYIsZmLul5JoyJBvGu+
rlon0xoQ2T54WmuUDkMJEkrIVdtg2dHuJWN+kj7z9iwn/K6/4PEPGtCBEGVF8pTr
NIoU4MbWuqaVXdEMfJyfXUJnmvUpbxUbfLTJHM1QWFEq24Luey9Hd8e0jiLdCEwG
Vz15oY8Sc1txLJZwyISiCa8sq7ErCZbcOCNn/USO1doWmcoHj5GGqGIuLN61NZd7
hnJKgO/6Ls2lTGydCBVQkBauwjXdilmz/TQe3s4TYNj0+IDF47PRvZwHp/q6gd6Z
fSZxFanoyIW4KudT0bACsaMVA5PGeeli2qTvJSTCSoV/ZWBuQQmEHILaYHj0y/PM
De/xR7DxRmnwIXNonJl81Bla7YcpCMpPdWNqY2QugpWRDSEyxuMpFjJlaYFdjb90
FRzcMddfhU0Qu/dVB4MfURIgFcTTHF753xKan9u907oB3s3wK9uoN1/0os/3jWxg
XhDqNSM7CJRmVp8Fulmyj911ihNM3XFfV5M2r9uz6zv/soTETU5uA2CD7CjqhmBB
+uwNnexlgw4KX2F3AZYwNsZFyTz8iG7yrMYLbCDYCqMkahI+yWcPt77jNdT1ngAh
xjehVhJsq5dPmirAYtNTFHaktBW5/AssWYWG0a7imx8/ZH0ZrYmYJlIaOnlg8y38
WBwX3aUaZoOcnaFr9xButK0L2Wi64nUBqL2q8zPu6YNe3YvkJIRonhvJfbq8MZEv
RofdXooxgi/HKO5QddIzzu0RviAuDVlDKLisHRlxJdin8/9KSVTRQEJXHd8ubdIK
QNjCdX1iXcfBFRYF3DdzxTmRtHPk/GkzFsFykHY/Q5GxF2xo73yc29Ova2g7bxk5
zbEoe2k86MVTqBJKZ3blLz8t5CeNpPaqepvvNDdpQ2jnFwllOwgVSlzdNLretJzU
s11jALi/MuYHF4ZU5bL+7gR8QrFlkqR0p4iPPjjoFIIw+LXNINB974OWe3at1Df+
dA6fm7wGJ5a9hwLC0rfFR8X9vAtBAW/miFfcnxTgW2blBjk64wSPysDBMDTEeHwH
Wwh4EGH7iXcPCRHYFUfnoqAlOynm+M/PWiYqdQTtwU/EFE2ysgkU60d1qtLcQLts
bJZKHzkV8AgQgmpMmIbkTZ4uQx+MW0fMyyA+uOgGaeq5/N4k6xp57aHPqcV1LI98
7XI6f7RPerrEQvxnNLTrUtIXAU9FyIY8F+YIhzW+0FxNLtlEtg5KLaWZwja00Ok+
kXXUMHT0is25Y/4b9y1Ow1PeqD+f2I/Y+nqxci2RSXTrNxENmqun89IjPCG5ldlX
hNKAwlGsGkAispwwCVvOyKidGsy5CfW/i5FdkK7dqb3/x5YvuuSE+AaTHvdAt7Zv
JblLYGoYqsaXF5TLdLm+ZtP7u+T53B1z5g5WjWD29ga+ABwt19VnC6/Rl+sia+DT
dTFs5kOEHTll4kDH0cQSHbjwTgEy9CnQhUqNUibEXWSQd2VRu9XAWVdZs+5S2DiH
Q8N2C9Qf20iYfmayD1lHa95dfh1IQVO9I/OLdtsjijNeAo7gWf7qW7jEsMKpesVa
q9GA6Izo+w7DdGP8X+X0Ic1jug4HfsprAm6MOHA7mZXSQTbqyEvrvasHfihZQXRX
mtuYeK9EG+E656WbhGtr4t8V1+vqP7JLT9LEmDsECVrPmtM8R1XJ3BQkFahsccuf
ccbWFCKCMnugI9baqISa4VUqqgu3DDOLyO4a2XfeJGflr8WbVTcr8PNxymDjfhig
jfugnQQPDUnTB7OB8Eu7ZUnFBXm5F4344lh6taeQo5aYY/HYeieUBsR+UJH6++8/
V3E5lD0EsFCHKTl4P1kX8XWbSoPAxeTO52eTbcipHCQmUuaQkWJ9uVpMW5diJRSI
d25ZGiQ/cUgjKK8Xl1eYArFBp2vFrnNti+SS16ADjLcwiTiIwVVlb9Ebq8nuZ5om
E8vmabELJ25GdD6lHwvuDswHcmeGWE0T8QTN07w9QVdte3/hT049Wz+9ZRxBdSpQ
27KV6QrvH/xDoQ5TNwPWYn2leYfFjX+9N8T+B67l1pBIsZ4GhTVAM6VZH4UMANRf
ux6JOMWIXLsTmSlQzwjaHycEVW/CfRqzmU7RH+c7M30dhJKpiH6QTxqkhK2E8otz
416LVO9T+4t6LSQxegK3cuUgOduzEJWRybAtbnBQb3bo2BqB9FPQRgaeCtYVEhM1
K/V7dDoGk/EGCEFzGSV6nnbDAksALbGui2zlfzen0bS4HPtFGPIbABHAW5dYLnQp
388+DxoE3FkNHuB229dSoFiMP8pyiolaViD6BWJuMIr1bPL3KcN/8nWcZchpu01f
wRqL5+JjpQJ6n4DAmr0iUjAxPJzxZcitTj93n1hErDhMLwdt+HVJF1w/uGkHffSX
yM4+Ja8fhSuom7bgBYPayade8ynr+4PvUIaaJcIoaR8Exd+Z4za5mI+dfEObUwdO
WVV9rCks4n0lQU5XW+jDo3VtUQOF/rX7sqJHDLvCA7aBUjEpULu/kKM+BdBUr4O4
Fmw5tibdVklrutBMuxAs46UQW16BOwTqf7ARKn9rSEqpQyA3acXv9xDfUBPUuBys
6iGeDBCSb4iAA3QsdodYThP3ZndZwvmAmndsFZ0ra086Xl1cDyv90Lj/igUbU2Si
e+Jq+KdsDsi66p42rx+c7Nj+ujvdHZo1rNknF91UHy84G/i2VI109uIWnpmIBiQP
YFnJ0Afe0jaOtGI1nQrm+6Fi3WbmuLQiXlJ54W/aA301b5/awOAQsf/0leZQMWOE
KwxCuNgUqtBe5yKW8Lf/Byt2B4u/QNtc8BcAu/bTNxEnM+yFhzxCuVgSYp4H2Kji
RkFDJqEW4jWZVvOoKFvocFNgaWHvNkJhO912M6ig7sFSfn5xERW01VUxg3UwdkAr
7+a+25WXnRsaI6233JE7BIPpfOTGp0bqoj9a/lvqxkk/Eos/y9L9mKQWcPe28Jcq
Ac5zj3Ez7x46udGMrZlgB3ftdiCoIASYpFukml896NAiRDp/v3z5xj1cFun7QK8y
i+WQQ+ZIxVCSY9ypd7TIRZP4eA1n4u7nr8pJYBszrhM7yC1fu24PyFtdVOZ4A1Bf
IhWQJnbOSpV/lseVZk2/hGP4HoL9nPWcG+YXkGjOJFTLgHarK/RoTjyjODMHIZMY
qiAdb8OK5mpJJGM0lLo8yogxdgEiatO2rSdN8U2catafXmgOPcieCgGL+wNBiNr6
buVBjGAM3RhkjV8j/igLMvMYF8CmflHmCNyvfCRK9EjyW7nit9/2YqUfeSNLTdsC
ioCZTZtjJt06a3P3ICrg5PFvqSwSiLQjQC1zyplaf99VMAXQwLiW5FBUZL4kEYGR
0RjSCLzime4ip7hF+HuCEf6OKR3/KKRVY32iiLE0TiOYK2R+EqopgWCBNUPF8IaB
bNTcd6Uq1cmAKWGwFYYLkkpp9mVcd9M7cb3KDT1dygqlThDRuA1x4JfEG0qTuXaJ
tIN1plsBmviIAcO3GX4XE5UWpdwkGwrREKRSMiEyVn/Jrwefbbdsx1uHMw6DY4na
FHoJuxFpAPKRHEdmbK3SCi3m5zfHPHp7uOA7wG8ds3zlUTWDjzhux2A0nEvW/2NX
wHnonkPZ0T89i5AIyTUxpmGWRWVuLfzd7Fr7yw37frDmjiL91H1faDO6dnw8oKRs
1dH8I0KKchUJMI7/SWyR4mUoQAMT+1Adk5MQmalwyhjRg9x+KslIO9/V1v2Qlgd/
dbc7RqK2cNmUjbsa1cwQjkl6cbvgdoJJ1e8YOBxsUGiH6JcPqYGlNthi/tsceV/e
991uWzX41XH+Wh3v6BEtplqdTBVsLktkBBQo4ke42GLAbt+SP2J6bpEvYkutO4T+
/X8SZlL5PaIH9m+GDLrHxIo8rjeCG0bRJreT465Ja4YJyuv1JiJIfNVun2yN9NZ1
hU4OF7FCIZBqM+h8wes97f8NAfATOEyBxkRNRmPelniReLDk+XK8NFG4NOODx82Q
ytSmLxS6/4k+tGZIChKXpw/YTCyA8p8WLqXxe0T5ANLt/quApXLE3H8JcXjIkYwF
ci5Ac51X8SqMiWGkilHD/7PQRz3lXEsaZ7F0VEBnpBsvAB6V5Tq7Za6lMT3FNg4X
Huj0EQVeP/0TJ3kekyAVhDCDEm3PJyyag2y64Qi1/X/G56rJZQ7Q/Klc/t9E79lj
AMNCd+nkxeAX0ybSIZ8o5J2Szgy++G1hAEu3GJT4gz3gzjaMeXsoaq8hKTa0CdwI
h/dma5oyqYcXgOjUqeS2uBPyh4LFONDpzD3J5SpUMyN8J5QCwItQlgtgx0qhoYG+
tzz8I/EIxH2T1d7NwE2Gz+KkgrCAXthRWPtKwwghvLqapGw1o/TBlZs1DFnZvbZG
+poVfMgzFnC2jZz7aY0sZLXeCcowpHWtlXoqleJankhF6SmP/XckeQu0dRkS0SaW
oJKxHT/mv4buGTDYsZLUiEQlSf+/ihLnioLXDd3K7qvdfKNiYzazCOoDV8usyu8s
QL9xspri1KYxqJvRTq6glvrZKi/t4vS73oFC/tSgJdCzOuP2vu9Ch9bKwiq0vAP/
14aEUVLZiVLFHY/PCdAKdN9cM2GVuZ17uucp0WKNxSxH5hgJ1rKUVzxkJf/8gMUg
STkeXwlooO0waa0Og1duI4Cuqm2WG0rhJn1tjTHWu2bF0a9mdv23XMFWp4uVyLo+
foz4ZVJR9+c/wE2iW1XjOgssNKVDklsQJkDe4gz3B2HBORVGX3IvH/9F7h0ndZgo
RKkjhX92wKab+mfQgr/uzCIs1lcC71G8DnL2biR7Ty1KL7Bp45oXv4oEx2sjd0Mc
dq3rNYS+lDJwKqSFQwP1UVWD3TO2VwcdDfGld62qsHaD2f+62h7oYrd7Wd+E3f1J
/geh2dXEYlMTAnuc3ZfYoNKj6LYsT9/pLSynsbXd63fqjnk0ZPtNfWsr8232cDy8
QNRav5LkmB9IsIVzwjrtElMH41+9UeT4ALJJspez3SQMIfdabycEguN24n5oolV2
Uc7Kj8JTAEfUgr8eFI4Quh2Zq9vVulgFkcTF4lpe5gb68d7TpKXKMQyqAtJx8fp0
oADKWDt2GvE+MWZjIlJe4WmL3ecFRwHXaPYzgpVZ16hGsltf913v2/aO3oLIeefp
rhbc8aJAQvDZ/oe3rcCCVg25etznB0KAThAK5frHpiEiUjUFg35bzEEbmuUB4lFw
IKGgFfICXlpuDojDLBsguqu/8m0GFzu6TdpRAGUsYep5jCPTxmI1KvbfuiMT8bj9
vJ5HmM94W9tikyQ/i9tZhm2758Y6rapSWChTa3Qt//DecCvTG4lfOP6WGAtSmwH1
6ZcOdDeHdsP9dj5jvOedIXlVfl7LyXUgfq8LNGNZVqvBFMUBuVScQtby0x44zQAh
qrfzCyzhKDeldszZKY4txVadWr+QHYFILewA0i/WHhlfDjGdrYgXoHMcK4ZaZCqf
ZTVAGQNDL7Qz/qIA3izjgbratmX1J81FTzxamUYhqz+RxejE9jPgijy34wA9PNdp
g1T/gUUSABCCo+BVDWjQPGeiDh74Wr8ye5t7NEiUvqQNoj2U2JezNxKNmHpD8Ixb
BOTNdMEwlMzycDbblRYOFo4YPeYe2WdmPasQpRPbwkZwMlYH/DwyWCJrpKjniZhr
NJ7C0SpO8IRr2+xmdR0sVAWHop+NrQRXLdeFLvZhwbK+MoKFlUl0QEssC/u5ll/u
uEV9q8ErBTjJ4XMVfI8gGHVo6NAibeuQhc+Abxz89AKwN+y1StCV8L46hHf0xMi5
AzCX9Mwz9jHpwUhCtHgvhO0iUTXhYMoNpJ5mow2qZPa9zCEnoVBGWCz0LgJepEe0
QY1AfG+52kyAXvKC22cw1eZjgs3pQWp0yTGcLUpFLVNPPcGlE/x0nMGnX8khpE8k
RzbZvWO7a2XtzPqFWL8vRzifDaPcY+64A5oULa85QOAcgzqL5sLV29aX+/FQbv9P
EMiALom+MPX70anaCnzs79Dnza9zRcVwYzqmn5PMjzw62rr3ACmhKcCiHBCXkcjT
CSd6QIje76M9irLjaG9x4aNI7Qwvso/MoiJ1BnGUHQxb8MQd9eWuewuChnpuzPdi
GZXZcURt63rv8WW9qfYyBSQ4o7nTdxiXktlj5mcfoFPvTSKyS8SHjquC6DS2zg0L
mwZd1C1DNEIfh5lmGQAFzmSHW7nV0HzutAda4F+EMYAxVs6Cmp1kT0KRd5Ed1NVS
cRgSa398dhIyUJpQOM7ob2LlCjeNWcLcaghXSckKdSJVpgxc9WllreaoO6L7ILnl
fXQOiLtbrLLdF7aK8J6a9Va0j5ResZpYemdXbRFQqNfr9J6BROHzOagNQJ+yRFs4
1R20idENUhG0Glvsrm1w8Uj8ypd9WFFaMlCP65hdR4f7UXxWqBCRFrCZAo5dIUHe
4bxpCG3JPE3q9Nns/T4ZxrLDuwyy4S3Gi6Uh3WXfy5zK8boe6V/yf6TyOAY45Jlj
rKQrBGAyHXv89L3wbgssjjaTeZYPvIMLzgPZWVZAnoFvypWvs4AB3GrXoepk+iMj
gmUezp553ckU9YCdWdIVHbSHWZNYX6lGgTdJZNdUq9Mc8XzYnKVto9qx4VDF+gOR
ZkDKkADkfWQpxlRyZ/OP92Ojm7jdqKeQUwAfMXyKo2IPkkMYuMJPUaIQSIiy0w/v
8sUwrZK5enIM5fu79p3uB8W0QejTz1Qf4zw5ZhsvvcN0KzvCgnuWkjdJ+t6YVHxo
mS3/7jOE7kSHuQVNUtqlebrF2dY+AjZTIcY7XvWnSmfPKdafF+NCVovMKU/tjfV7
+pr1qCHHR1J3VPtyKqK3DOj5Z86Hq1pRpOoyGvMnbjosAIJFBS+iIPAPYak64c2E
JGZ/fvSX4okznSeDpe4NnmkypjrgKxuGXMrSDntveIoJR+Ydtc2PPFgISfNbRPbV
IovwGjmRJD+PCNIwabvljuyE1GBDCsvDlJbyDyMKhpx9o29/1uIfSh6zwsUk7awV
bNA0sEuVOSmWwTeoZG/1G8o6BDXrwEGQo1sUOKAVtam9rUOey2pvfEswgnrmZu69
sP/xAyp3TAs4BGKziILWYAWJ9hkxJhsWt0gNFW5rVRgwGRinXiU++SQ2kpmgqroE
bxRXfqZvwdhyIuXT0ubU76tB1wfTC8nyrvTEnTbZNP0GjMjkf9pTLzvPGgKN+vCe
ZT/uaW40ke7AUkVmo9bZfHqxGi56OzzNYIM7G91XvfjZqH0FMmss6aIxx0SxhboJ
QStRPJIAeWT7+HrfK0ZVfmQlCQ++cWZWYbMT8AsIMadBuFNxtwAY6OOBmduG2xnd
2gPCO9YoRMoojem9uaBxZgQ6ov89w79IJFp4R4qKjvd+FnhoIjRF9k4hANGf2hSL
EyfX9lzKgEJToeMPiaVXyW/HL28Vq4tLIoAeGym0s5+ooDf6wCCp4j/FRwqTB5uw
DPdOOwhfEZX8ZKCjCHn5Ir3JEt/px3aiWg/Pv+3nqShcEGMOnzILOUMoGtYc4Uy8
b8VKO8I+jEpNqkay9jq0Td4r3RAQS8dz5Ip3s6tkC5IWPZhIQaxMVH1By0fhqYvU
OJbn+hRYg+i7apmVrVVEAJ23atGmHuWj/dE9BmiODoPTuvUM11yHBpPD9PAVr/Xn
41Lvv8pEK7LNPqQXg7KkGd6Ym4zNib6fsbWaCuRGVdieBfsNgz5zom9JM6VReJYV
Ryd2BOTqAh55EW2g7fffjvJWvhfMwv81lJlBzCjQ4FinUBm8jCuajXgTGthGLqiI
d5qphkNGSvxVVazoXMhXolHEaYXcFGb2uvaqlOfdQmdooVCOzorDPlClyCb6iEwH
y3Es15D1ldrNmsnJDVhSAU+jYc6YXGs65eqBX5l2X2SVbuddYbh5DER7f4RtUIXc
M7KWrzuO4OeQ6qAxNRb90MuKNjcAinuIj8GXftrd+jSDu7rXh8Be8D1TySTzYvH+
1wdV4wxpyyNVvWqIBxaeAaGpkSf90Vj55j6V7lfgTpvrrkGOQvGLMsiZzV7AR9BC
mcP5ifc05e7DvFWYne3eGKCHpCYm7EYSK984PL1mHaSGaDpiSr23qvLJyjhTizIi
t5EvHLAJvqQQS9jLYGm899LkhNbV72g3mDTFG7Jt/jaoT2nqZZYeMDxhWqZDQPh9
PAAUEIrKwtvTVdAGejOvPY2t2tdBLdiudZ21LZPpEqywMSZKa4BAxwRtwBtNbGxZ
54eReVKkMo9yq59cCpEEm613OBJG6oIzrxnLdI5Yd8titITKfVSFvqgV7lHAoLFr
8HoiQSxzribHAomOLydsRvElKus2rqpybzsWzM+7FYD86KqCuukDCcV45U9eV+ZH
i+Dac6B0s0xAA3qH5a3R7tLo9HJIxGfyraqFPSdIha2I0RTOIqVPFqZF3WvLa8i4
sLZhzWSZB9Pkf8YQEAObqxd1BkqsKbZH/v4+/7vOpyX0YL2AdLqZhgJVGoadF9o8
+d07ududzMgqeJN/nCMoXquK0H9IWH7TJdoxQEBsT98gL9MGoZvN+VEzDKPfM5h9
/x05b7/gli4UV9ydOIHVEeyTxaqpgkcWi/A1gFGFodQp6TxjJ6IDSJRGvkvAAJr2
5ihyN7fpkbKveQ5cmpDtfQGtPtnnHiKBBHT1oDXnuzZBHeT+VKwnXt0yXcyAWSor
+3hSk+2vZXYCYoGgbIcJEstyIwoJT8iSPl7Vs5aVDntrI/t5CVcrnL0aHuZgBzY0
GWBGNw8dpNKP8HRbLVEAn0VEzoSD3HSvvEv2d2p6ZPSmauGATMKZH3RNmcf3FQax
8nE6JOycCCugQWRjJKsqnBCqjP05b0sP00NDIdjpRlSjkkSNLg2LTvbuDCdgNi5r
tanMsdphEdFMybyGjKCu4BpHCA+KIiIF09KR+YviT4GCaCFeDr63EL6KqAZXx3yq
BhlEOzfBcedop0SgoOROFqLBE3c50VZUXXTnqLfvtvqdn4dUmTStVB21NAOltCmx
z0sp2M4Goxj0xlHp6t9zcDHg4UpB97xJTBvuO1GkToGxmRLCi2knwgTO/v9u7/nM
/kadxKzvtjx/iFTZKV/juMXFFv2FMAu+cQau/gKSGGGdqScGYImOkuoPyQYWnGt9
KkaRjHNjxIl8S2nzGv74tur5qpQvA0PLFVEEedS/D5uALgXJnBJyCi+NbaogBDgp
PdRRs9IgIL0Bt3svbW+MFUbG2DH4wMDylwpI1ZIHXpBF6yT5OAf5iFKmQGiEI11Q
Po2X6ugrgQ7hITz2acnjs2wNe+FX/7P+ER8hRV85ZwmwQF/auENzUeNEm26EgQDZ
iJhpD/1bAER8+sfpchU9YAzKk1Kp2dqkH2Yke/5DK4erxOvnA3HIkKPaSA0NHb+W
mBnecCj1yCDK78j3G7g9wPzbCU7Fzy52glOaXqPMarxx5ZRAkAN1rBlJzPhmHFcR
APYBYvqH/cQPW6MTCFHZjcOCm91K/usYV04/PbTTmc0uIFw+8oSwKjIK63FMs4vL
ry8fsEHQBl2gF4KWqshxmWcDW8VTFzH4jNYV1JD998c4eCffCCX93/aTCBAtYaid
SEa3yP2SSICuPvzPJu/rOVkZzyV7qK0fYy/STA90cnHBxX81ODPGTTttNwk7fbsf
vAYdYhDmQo3qVkqLz26XNrfhte1fnVpOQ+cjUMYDClvDRy0BdoTb1Kvu4OQn2O+D
4uRauYmA4XPGHabXPLeHIAQ60ASbnbdsP/1o5w6nUNleeA8a4Jc2Yk5O0mug/BQv
MpVd3HZsLY3djAeBbSKcx0exnTo4AHUjixPosfQ7cCGMTD2vf1m9fC7jhqNgWBWX
LyrGDlvaQ1Eb5ZdDwZmOpCzUKhL3OtKWMCN9LaKm0htVrQJ3ikwWep8Su0muyI7d
tWiLSxdImk8hXiTAi40WzmZWcwasq23AoUb7I5i3tFwNloH+b92v8Ylmtt7zkwna
QYuc3AgpuazMw6bJGv3sj+Qm3XULFab+7A9cKeM7rfL4ICZosdevsMHbV3czIBi+
MWQbCZ7SCccUQalC3IkGIzXWvYzy5XW95paxQTqxpBjsJr/aupy1ywXCQhDRl8ly
FvzRQk+DYfqPZlZsfTkK/7/jbqTIFmQy/mCvn49twDg/AEykyJ6t+D0/JSCqIkvn
z4sA5abBxmVhCzn1Z6WLpRVNMZ/uH91POR8b7u5GtPWJ9gnf6HdUUf5cxU9viuMp
Wu9pbFrWVaZLBBbX0/PV7qB511WhNL2upLrrWSyNSinBG9olXntrbIiRMz86fn0e
yuh3zHz4yOSWo1zdSVQyypjLeQWeRq3b2fo4y8AgIprMEVBxTwj46q4MsGiWH0aN
e1HoOnpMI/IftpqHCPJqg6UPiZNGlEWh5uVco2Bh9ajvmJKG3xXhBF+borJNSPq1
QcjlxMkVEZE2UpZW+rOw56kmLV3IwKfhKSPFJiOjZSaUSaEIQSqt7HoTBM8vsYJQ
it7lBGcJ1YP+NZj4CCapQArjOY3AKhT2jCYQQNLEjt2/vXxTOynyMPjBjyrbB7BA
dYDOaOuPZFtbzAlIx+SDIEDv3qcOjMop/tZe69IieUgNiBzBuuaYkFMIZZkzAT2e
0jGzuxPVt+G1AWcPIzugqlIjvIZ0Iu8ECKiWu4DGVR0+YkozDbV5CdxWmNmHRuBY
cWqxzs0TBsQSOrqwvGKeR/2SZfCUM/ciflipvYxSdKwzRvnnmChrDJNlneJX1tyb
jiIQFygJS8HTWliyRVxUJusulpY0Lsgr/YQEXJ89XxJUAaLKwOt17lTqaNDGfznB
/TIg4O9wh4LDbuub4cZ9/0NCWa934y+lfMmfMRPyumzIDlxVnrrk8x0Lm5DAA0f7
Hzc2EBA9ilaExofz8Na1ysn7xgaqRwMbCuepNtlePZJRzeAkGbXAsnm8YCTKjpjk
5iqtTsM3sesi3PByXpliHjJAVEGt61Lp4wA+JYeHoha/rj7p4OOl00C2XtFW4IhC
KhEzzx2wE6MvoeeP0Q0vM/aGbE+OBduvdHMHwfqR5iFIpCAsiOO+Kth3Cn2hvkDa
puVUBwQLWJ82H16ZLvdoFeBtZFeQRqcMmA6oane50uC5NZlJw5aYlTxNbbfMfLBc
Lopaq+o/QaHFRcrfnpSaa4faQuw/dKlk2u55w+R889PgBgsrwkdQL5mtSmnJoFZy
KcIPkflSFn5H+TZ6CMSlWaXw7ErD57r7QA/nsW2+axtjE/dUCRL/bmrOvzhOK7+Q
8VuBEBO7U3lblShtFAQwyREqY7vcstpRP2ymQk5PkPLF+GxHQZXs0dDcabj+OeQR
+Tg+f9TaUfG9+tjX3H21IPreWN2mLvq2sl4FUEmsWu3rHafMvAcXor0Qg+mGq5y7
JuWsNPhrLj2jaToEPVXjz1c2j3eikyixDBL/lHOArOG6zPNtfdSEg1Ir17GaYvfm
ZTiK++9K3igSHIGqBgK713DfZTUZL3eZCDam2F+QmmYkSTNW6i3q1YlUHutyulWV
q+vMKK2AcYl1Yr5evB3LZcd2Zha9ZCbsQA8VAs/OrKrdMXU9EaaVGb5PLsKuRxVM
dVN8TMklrYlFhBOz5FmGOgaZT+tlgWG0Cm5YrBOkSVLAfi4TzpiGQFyTUimpR4/f
TYspOv0yY6Xr1qM59zTc53aVYSIGXdaUW9ipELEwEeiMb8TzDoB/QDkglS8mlTD1
MlvTJok2kJCC9mE8M9G5odrADM1imk3m81yDTD+dkmyru9cRkKWsvFe3WeSeXIHC
zmyX38mK46Z27rBN89d6K+uXCjqhzyGuP6mO7f2tmtAzqw7lrdVuNHoBtZA9U463
lTIyTeVZ7o1fWuQ7VjwUgfwWdz2NbS8cp+V5hHnSxOeo331TtJVcarV57wD/HcVz
5rY8F0dllL3lbdZcoDNGz1ca1YfQdISra5BKEWM/rG2tsxSyMnN2ZHko3YsK/EA4
1jBFbFnRwQb+4uVt3eOmCnSJphW3A/Ke+BUoJpM5ggOS9PuyJDNH3beCksvlUHpp
ICQXAPfHKkl9D/IVkPGnhEdQU32Z6qQjbV2bRk1h3754GCOYtAn2qvDq0j6FDLXV
JriWo/uyb4r1M0OOMslXaUmFUt4/ilNu3ElNtJ9V/RopLQwqOyZNHw0QWtB6T0nq
B2/9/b32Eu0hHvQmjjvpP+u3ksDOog0T4k2iNwLZZApbno3s30T3rEE6QkDL381u
4kZOj+o7tLyktrUpHmx7axnzNzeCzYTUdKCXVg/zkBmQqBmITnzTXFVVSHziu8Rg
8/ZZfRPf++PLYbAgB0wdytE+clNJfcTYVMlAkXlDSeuQXzIQuOAVdAkEb+QfCQ2w
Si5pGKT+IpvjA8cxcS8L8jDQ2kPqMEwRyqNPQIV98JNip6Wpbzc84SReKoQWTAiC
8pJD0xAZnM5LoDqPw/1hBkbKCbmqxlv2gHo7cwtsGgm421uOZRhRdJ7VCnRFRhJ6
MLtZQ1jNSK5djOFOs5RXsr2CqKJgKsc4QaPtUZZ6C6vtyCfU1bP4uLIiqlJRUV2e
6wD64ORw+ZrnqtOjvSAOJH7cCs3nRoWFvzCiXWpJQo81IjB+aJuJSbW6wphi6NkZ
rMb1cMv0AXReSG07RxAPzuR9ADxOg5cxCX68queJlbiXCYSiJatqAmfs6sVOXryM
NB2ZZ+AiHsfqlAfMHzI0AyMzPN3qMBboLjuz7XWULnq/Z3sFhBWTkHuKhcMfPKPQ
XqvBGxDqGUAAmmppWeQ//42FGagUjfVcZ+knug1ulHRttiExfY0sf+Hz91Ra/nYK
9HLiNTjk4oF+022sEluBD2AerO9AUZIjlXyl+cNeDeV6IQdo1CmaYlio24cZNUit
zpYAWXjnWheN7FbEA6E8kUi3i9ixktn0H8YjmbNJrj3B81XBHnbUw/2O+Co5EAKX
eaFHYTQlp5t83YvVDK3nZoWTzAIAnvphc8Z95SVLULrIGKCeX/CpQCd58glbM2+W
EeZRVc+usViZXBoa96ZNsmGjR8ZJCfYS+M3TYpttaVyv6MggXQdO6usp/H5ocfl/
OyoTey+WFn0Jn0jygB5lUZ0dlvW/EyoIQs7TsjLESr4GC/6365ilTBeTYZagkpBz
V3t4hUlkJv6q7o4nrGe5MmV5McQA42IMDKPP2Cu6IKDzSYE2KxmUVr7sD3nJrblV
vBXQwTG82b/tCKJmaZlzon4+TNXXUfnPQqsGP5RhQRf8J05jOh31e3w2iJZKSmXk
ElEM1RtczpQe5jzWJubwh95aVJ/FCLUCo0yV/VGcdqzkfiYtXkDiKC/jODAAOlfV
MsYUegEzpll+V/romMDLbLytvmDfm+dLs48M4krXeAPdQ4lklNDCUfiV7mF1Lb32
xrt23euMynTsRRvgy/o7AaYRwiHibqfX2HcRdtE7Ob3GNw9Lmp7tl4jXVhN/gQyA
VQxia986LFncklPa2J37+VLB21Vatw3YVpCVZ5l0yBMD1nEX9mU62Zcv0Kw6KykL
4G/aOLrsBKtm+I3FvtaYLDFZhkwMs1lNV1SB1ShwxxrOHacC9fW9KpPHT50OlK95
hIPFg/iVAhR8+H65ngMB6N+RQCG+o25BGX6OWQOYQ+laJGg0wip6Tnfx5U8MSrbO
dPGDNU0Nt+j+rcbNnvz4ekAh7tKHJXI9efLlN2IWwINSMTrw/2tViGJmm+EWy04B
fdGsP6ZlB77O0UqmCYIBQaDSxu6xi/KtnxQ33SHx2+7TTaAX232MG1CXyaZEvm20
vK8FjvXcyVEB/NbuMX2bUrvTlypLaMDUmNSVc5c3KR5CMuh4YnIPEVnsUE6uyaDG
hjOlI4CRdoCQHu9PO6e1gJklBX5MSQPEdn8Olo4JF1FRaeqMAmlmCxaWGexA5nVF
mqIXYWYu3PWknw4zTLZTldNxoeb4LYD82ZxbQIKk7odefsZ4hCsdyg7nEgdJOyQh
1o3RJBg3OpkPWUc4EK+1ZN2AKbOEAZit01IWgo0iPewtXB+EDxpiOGxygj3m3bxy
IXHZsawJWiBt6X1CyBM8N3v9yodIIJlbYbtoadQmaHQcxCcyRj25EWEB1bOc3krv
WeMpFeNswLJtTvilHHvjW/e40mBQP+WLArjb7gXAw57KSx5g9b+zA529aD33o0PJ
CkBdCuN76A3qtIfcrfT3N489A0SMhhAunkcX5+7X92DO0hL4SYoC6CRuRS/esmJY
7qqG7ePQfzLUexTiW2NqysanySMPo0k5uL2fo8XIocv1rydpXaWirg9kr2l1IwFE
I5WqH4ghndMm28ZG/d7tCdWzdjecpMiQDNnMpyf8HTXBOVySPk+zQY1uQalPb7Bh
FqUe/5S7ARfXcMOhSgZLPuWk1tOrRMdUAn9UgZLdcz70KDYHHqBNICj1LtSZdtCZ
pg9XIVdY+EsKf9D69p184RtkM9ayCLIBLLsNsR/MXJ6z/76a6TXZOYoEfsCZl+Sn
zAgqDn2jHSTa2sgH2OBuO42K3amfmrzV7u0gZDJ49i6oedn6dHhbAVB8cqz4OHhT
FojLm+wxsERCdt2oZ7hTNFAlb9z0QbdDoFdO7h5uLgFlm5fBe7nUxwWDCDu6RPFP
8DjF34+GERY0Zn3mWT/sVa4I0nMzxPM3+DsydI9PLDYI5nT4yoB4cvR6UnMLmV8k
RUbkOMuIxX7W8oE2q88KJ7bWSpOElnuEUOZafDPFK/uBl77m5TiU+9zSMYLkSaJM
yrkTjoiyYRPE2Z3OMXLJ7DeWuwly7ERJEzSxbteyFwovFxzrZSUYWV0puqX+6wte
u8DWD7x50ha04s2VF9D+X0zJ94TTD6NW1VlgEeG/1jerFmOrGx7C3XfifYu+pwG3
//GrCQcLOELHUZEHhc6mvg2/fbnLmBW+qlvoVEWrJch93VYBP+G2BKI1uEaKoD3T
R2gJ556qkqdCmNZEgC+NwPqc0+eZzfYXG+ttwW0FDI8/5pmwnlAqrKvyWsVTrVJg
bOf7MW+vMbqVi1Hme03mR69KEhVSnn88VzaPKQFmht46IjFCAHHI6wqdFvK7Rnce
+EwI3KthdtGc1ocxLesziaqxzVQWGzc4/mCjJAFIUEScwsuJG3hPQDJN5hJDSswt
fDuPHAMm3UEldDfY06jYMXUoleFyyyzJ8AAXxSkIAaYtHz1e801mDccfpXaMXnXC
SsaH+bdqq/iRze0JEAacC93wMG0FCTyLDp/bo66g9ilQURI+RnwrqiWbpFnq+xTA
T24YH4X+1DOXrWEAwiQxBSgmBGbLd+n5rLadtdnw5tzuPUDmi3xC3edRTJQTM397
IPCCDVIjlNhTFazi4AkEFuTs7lCjVunbnMqI/Yikz8nA/M89TKUTHQMvBJdWeghc
z9yf3o7na2UyicsbHUdFiDgmG06XAtOu6mtoSIze2fUD7xVLNQZk5RnHBHWjxHbw
J9a/TK1t7m2BMP5Ei32cyTtNaxlX1Kp5M8IEof8VSc+LVgifp7YNA2qI+3FM7N8G
szxhY0SAMLxpBmK7nFydPJOtnc8L1ho+Cg9UGxBYlDAJ3bu2W0VoaFHNCjM6y3Cs
17dWTZuqdN30UBfGvY7KBRi93Y/VYLwiEIMzlxnUtYvZkENB5Q8XKGHVCP7PoHqX
R4Kuza+5kLJmqnfkwg8q1WtsJFNQLh3GBlN/YyyrPXNhPiq4eOFRQXdzrN0zFIh6
2LD699IVGagzu7lrUDKTed+vsze/3/Xj+El0eGbiPrj0AG8PQNssB/P0uJUf8GiO
kJDIIH8jHDONI9xcSmZVpYy+8D7U+YgoR8bKRt48Qc757O+Yvx16L0CMGRLovTcx
/Pbk2VbjtA/pyJZ88l3bIVNwx/oQYZgW4aNnaYrqSs5FyMPAVsd7PXO75yXBApGO
/KLGHYjD7elaJHC6A8Amt2bK/HmX/ECKatxQ7KkQEi1SSacONtbHDbTEq/I1rcLr
6Q1SQ6jfkQUuExTf58l8yRAX2gvpIuO4z+cU5A3pyESI4fHBR/z9R0bT+pCNFDCs
REvB0szXaVVS62U5S2Ecfs2qd5W9//sde+fzVmOowBVlWL8sTd/+ZE5Cp+QN9Zok
ZwyyrSfnPqfFWat+np8vpKrRfozK+PSyYjWjtFFVbN2kzkXfGuCJmZwfUZe8Y9D5
NPfxtKRehmw5jP5ZOL757OI0K2iCC2f1xrXanYoEJpYH2LVc8inNjdOiFxQtwGi2
xgi809KctYI1BUGXvOECIh+2GTIcXt189I3daT+x35u8+OP0WrMHetRRuwVJVyAK
xSKKmGM+1tF9wgFuU0B1v8PQjl756wxB2UyOMPvXBCrwQXi8+sxGxZ8JVEbXkZb4
R19G2H9RZOZ8JDq7WKFqv/Uiiv3PX8Vq9dlc4hraS6e1v0BvCphhG6KTtmcTLI6L
qhGSwsf0JpYDMMSUqBGCBxlOvOChMaf/TolBB0suAGd6vH3PeLeJ86tnkPNQI7Vj
5Vxp5f9G5xUPL6njJ9qVk3W+1bajloZ0QaCrV/pscAiShGaBNyFIsjDQNz90qork
o/UQEDg51vj3qSnGgBWF5whwdALFmuWJE6Y4biVD7nqyibtmiqlkBUIaQ0LkOtbJ
6pI19FctptBOaf1S3LQACezLPJFtMJy/HL1vPI7opt2EybNmIFcM4Q/IsCXd+9Fk
vDGulC2KsiHtW7OnQBtlmqyE03NHdlMaLON1K03PAZUysc9OXS9/WQJ7slK0Cl8Z
YqNRvrS5KZnbW5pnachDvaRnkysSXW1I+Ji2CvJVm7qLn+36Qq5rxbOZtmn6Ufcu
M2lYm78cfmKSF876cTfYHW9jyW/KT3m1fjYxBnEsB4WjL0nyDiLO0m0B3/lvm2Y7
ORYgbA0NKBSVmZcXk1J/6QUfeEpw4Eq1cU5ceUjrqlCj1I2NK7otSO6SR3qw+Wb2
MagFISB0AoQSM+1VhXUKaBq/qC06Eqb4sJnFfChOIUjH0WTW2HslB80GLx3A82jp
B3Xlyhy01jer60WHNiGM8cCVgcvmFR/j3V7A1H81kvAZJs12leSZXXaz3byUWFAB
tOU5pMmiu5EFUbTHQjS+WWJMdVetnxZpKeLbe9V8LXNf1b6Yr4LRDNfP5BZnbPX/
eAdpiptkAYdMjgNcyPhdURySwEzk4TsYFz6+eu8AAZmZHLLv+zJS4tdARWtCh1Eg
g5KdpuumPPzrDCo2tqxZaMGgYYDiVYCGAYMD/JaWYmz/Fh1tJMQmw11MRniau1Er
zW0OZ9N9PDXCFSIlVK9AjwkimY8Rs5HMxS+X8fC/RCBNRBO85bOBv7q9MsS7t41u
0YTnacCO2P0jKrSYXrNALUlN27uiWds9BNKLIvK+SlUy46mhIXLamMtJvD+CI+Pz
92unY1QRKztq9J8RzKNtdHC/lxerxRlPN2ZN1CJx/KySe07CAzP5WJOrrTjhvheG
BdrhhaU4/rF/JOokiQtSV/Bsz+KWhtV1By9JFD/QoeYjbgXseiKUBaiUjAauuR1a
OmzQZs/MomcExf2UqTWsDQThhojAG3RKPvFhCcR6mUAG0dIgA2vdNPFnfXA7kG+H
Ux/fuIuBoapVHtlZTd+h5EtqFVAXJ7LK6r08hKxW6x7IhK0gltxo9M6e2hgac1lv
NPgVM2UqPUNkkKM5eapHqIcCrcpEKBXJ+yw2mos6nJoBn6U5eeRio0WVsbS5VF8h
eA+uiLNj4AmE6Yjrnxh99kX88nELCD56qOIyh6zW5i9ucHHctQLNi5Jc/RryRwep
v0kMQSzM2eb2JT9WzM9V1UKPokXsAxbsQTssLlTRD4VPawNrF9FL7T8eIKyMpV3E
11FLgtQL8tD+6qGyUihX0UidJwqonMpzdXfFxOn2jU6VUIEvwcQp1WbfZGUFW1bV
gj3awiuFHkliFyo/r2QNO3UtDjGlWG40j8Ura5lwRGC8MDU+XKS7uyR3D46p5eeC
CL4MrbrM9qbT4BrS+jPiiahOswqweFoZh7EHuF9l3iLST0FBvNBOklRgQKbqbsb3
VASEjxf8AR6gq7ZYabufq+R6dJtPHtr8j0JsNAkB1R2GbJsSD6LcC4lgGwhCGcmz
HonY7hzxCYKKGfLVcrFgqrsPVjSopV/F4pzEc19oq3gMXCtrl7jy9ncTqbZfIK4D
rKKLuv+5mSx9y9KLuf43XH/iakrcrbi0Z4o13EyTq+EBd5nFqaqpcehDzUhRHrSk
v7bbMobkbK1xXdQOAnXp3f+OmlSwztcV822gT3DMO0FZALBmcEoKtPiRzu0+1D8o
cRF0rxLTs4HMVEokPWDzvOlvodYS4xXX9XDO+pQl5gcZUzWyUjJ3pWP+UC0wTOFM
v1s14OW15FsbaFyoSv2q/klapt2HAkEKK6vA82lJcHmdu+zsHIP3ybJPLvARHBLA
7X51vniTP4LRxnwsqYVZ2Jx60uDuEAdMiTot1DwIen3bg1SE/QG9XRlGGhGPxVb4
YJtd57edGNDAfDr8CrvwrPqQktOEUhbwKPZL/oRcl0sXG1m80O85n6zWT6Vc+ceB
LQRHiKi/7hChrSMJiZFzdJnwHNj1i/ioFNOIygCo4P1mzjD02UhY3IPsxVm71OH2
/O49jaGXkoiusJxkzwLtdRSz7Ck95uSfy4brYQeeBHH/oXOqKqT9pDU7OQOaM6gB
9SU42P0T4X18VZI71jYiqimxMVORqebmG8z0vU5NQRs22ubIDa0RmUgKI5/exD2R
1Og8S5xnHkHp52gZYH2YcFmvNALAfczoXfYUxqvdtddI4mCXHlo57St9oUN+PdMo
2hVTUTnxMj7jl4N1a/ohbUhsbYd28t636s71LAYd9Mmr+leFKEQ89SFGxFWBy9gx
Vf3kjdcdFS+vGdJ6dAgBuv7s2tTVqs8dWvOv48m6euv6svfPwWr63kVf6xrgrpz6
teGAG1OZDTiQDKoRJZGY2SpdxGgOx5yqmBm12e/GgeHmMFwwNnI9QNlZqUkrTcc3
2yCyw+ieUvpC38R3Z8h5ouVP65VagXzvMIOU2TRm3Ng0v2HkVAoDBgv+75Lkk/PP
ElcsIFkIYy9cCQh9Ni0PB9HpfPKvx+BHn7oXqs0idd2md0n/O5Tu7Xy9DSbg5WrZ
gP6KKSCw2tk+gtCgijpSQt4n7nBlsdPzN7c475y87cFRgmX0g0YHw/sncEo4p02n
mZaSHJ9huiK+8QTfhDPGGC/W4ly3WVRXh42cfv6PbIXn54gSFRCg0xzN19wd8g/b
AVqoNnlGqQLdNL8tW4LNPzZQ2LMUo0ueFe2d96K0zPlqLaJuCIIbbHm3NI+AHWqr
SE/GMTNJvXSI7QE3zycAo6uf5T+STsoHejf6LPnNo8O076cBaH9gn4ECT+g9n5s+
JwNM5DNWT3LOdJzkSa1bXlCKPZsdqW8ci1yEJ+oOOu/oFf36/M8MQo8MDCCkSJwj
Q7d1D09rrtR0/zKnBzuSk/i6iKYAeX/2dVgrhQP2AB5QMeAgzGJeTzUxVSa91GXf
6UcKjps3oXTaOvi17dfdcuoPgEXmEG7kLUqjlFBYG/9FFj8xOr2027Lf15GpXlyn
4RxfEuhf9DsvQwpHDpdtAz4ztvkh+uwcRr8t0UNJUaA49BMT9+DF/qlZmhp/2Jw7
1lp2eKs4uHyaJp/kdZ+DYHfjhBPql+Edl76TnOXujfC+Dy4BA8gPWbyx14s2vrFY
pLf0tHiBcPTZXq02WItJlH+5j/CDQCfTaJeOh62d8vOOlkw6MFd0RDCRav9QfoXx
6Wq0nWgvXduE6s9UgBiYotngMUS5CDS9pXEUc4VHAXjg+pi95fEP+6QubFS42xHE
OtYt3mw1p924Yg3c2yqaIV/srZ7Q4po2PKOG+52DipQA57aEDMQiKt0Jcp6bWI1p
163dhnj94cSPUZL5MbJi7pwCYepeHyHHRKIpu6byQnVJN/UKfcy0cf1i+css0jSm
atbwoqZILoOlC9k/u6pv+O+WgNplMwgn+aXlwt10fCoqJ0ktdGl0mFpPLa5fB0S5
RT7vL3GHnUSPvsxbQ1YJ3ZPEFlMmeKxLnB035nPH8Q3vyXZ1kMxELy5uJKtjLuwT
4XHE3haKGvHgX5exVrBYpHKcEMErX1vNO2728UtDYmDsizXqNGl9IalrU8Wag4oU
E941IQJi+XXy8JuhS5Z6ehr/dIEe1rUGlz3P2o2fjLVR1Fm78WnQPgCAW6ujjT19
e8iQ3NO+X7f3jhnsaXhOxiV0RXEBsJ2cGd/E169jrzCrwJNO7pLNSUDr5QN+YQhM
z7UcRCsJelbv47Mua+xiXh7ybjy3w+anVQI9JBzbQpD3bQUEPXTz0oc2n4h2wbMn
rFPOLlJuZuf3S1pFFoE4QYVevz43EX0x57uAD/RDtQHVK+GnZwe7cuRKEISzrk4/
q0xKio/2tKrui/NUVlNGsGQaQGIm7N17uNdcvTKjWiAFXuYe9MjCtym7xTkllDbq
F9KjcjzaMiapVL1hIEr3cwCR3DnFkizQeNAd1jH13CdViG+FvPlyCr1FWxksoFjK
k4aLp9Eo+UnhyrIXDuMipwG3vOFOZn+dlvODlkfXuB0vhZl4Q8+6J/eHfh6eCciK
kCWIV9yIgQO5qAu1K4dm3FiUmGYbdFd5+90n4yBf6uz0XHFsi4M/ufiEMqEGjty5
XGRENFbZi3SJmNAPr3oqtbk3DljhzOa7VG8rE+f3t3kIvMaHy++6HcNUb6MZ33QZ
BE0TZOvDpqE2j99Y1uE++sRt1QV/Qpxoz4n5CZsDPUKonBDHMkWQMw/kmaZTok5P
dWxrchD7Du/D454DKEmouIVmd+HEKS1Uxq1WX2t0KNBmpg2hKPQWTbG5TvAPyMMO
WjhRelk3qSBapSBNEXmpssiFVynFZp1Ws58oNPXvfcn+ohgvSMaz9iTnaHtWREiO
Dxj8svbT5MPagfqIQT2p4+TchpV43AAiy54uYi+qi+ma1Mpujxw6r69WZISLhKrO
EskG07cbgvOOGQln0JnkHaxCZq+Sw1hzUAQz7os/0hQNoh/0MyeNMYfpA2gIB+Gn
DIY6Ru6/5owowX4fUxBhj3bGOfcF0BscKOOXi/RbUoG6XOZurX6PgM0NxB2v05b3
kwzs+MMe4tJEtz55zb3AZnyOoT7loHlXLkObsAKYG+cl32DtRRugH9kt2QI8dpKV
R+7ibFK/KUfQkRiqfIYQtCb7OY9yJqiKHOR3Xxd0EnqVJfpKY2jDdzPOaTbM2N/H
w6W+icEvKww8lacWpZu6YhloeohTx79PPr+M3jq/dvQyGqnkgmXDID2PbVRB+DtF
6UYVzYuYSCrqspbANf1Be+8ePekQQD21VmH3sY8lbleSfFbE1b63Lgbw/J5CpB5w
I9hy60+OlNFc8nbGYIFMTMJoDzbz/ZufkfQ0G2hdTkOlGrHtS2ZIN2lLwD7E1a95
+TZwZzKyTNoKezAmMngY9x4pAagCjhDawm+y19ux0XMG7PEsUNiVWw+yvTclPCPG
ipLBbSQsFhJQjezsKx5/+T7RYvGPuCsKxv0tldPo8OGgjaN2DKuNPa4l8EhJTIq8
0wd+/d71Hha0Ch/5l/U7FF4XdxiFKgJS3ZKNtTIQqEK/rPCfP3O0nmjJqwf5u8D7
XSiSve0sv/AK/D58KZti/D9x9IGit8gAeT4I3Zp8bSm6e0SUTC3sVnWvPFmH0+Kq
3oVxKh8RgiYeZ9i8oyiM8HU9S6XT2hpQ0/s2dh9nzQCqOOH3+iy3+upkbdVDgqFJ
txMCOA4+f48IGqJPD4Il1fx02LpYH3ki7f9Ksek18VcxmLrIENVEBsDuUginqjrU
2aYC7az+DBZPWtjGhbJCrmf7u54cqowb1TjTR3w3vmnIvefA5fnAyVh5jCohUrRN
uo0NMwMEjCiHMRwYVzKUpC41+JC6BU7gDTUMq7hHjZLtpL5xIyjaKSUzH7VhvH9V
6x1RGmQvjYbhxt+Q19xFUglQnp/ydEGUrgiuDT0vB0Uf37HUFI5KJaUDNB93VAgx
sXnkBAAo4WqTJzxW5/Quu6gZfmNiS9iusJOxPR28LEijF4vStdKICr9ep/ZR4GiK
tOYUTiNyjvR2RyCpYkjUw8JMglsd9dasI30TlcooEAYX5V3jlXPV1S1VoOCdAQsW
4D7Ok2X1MA1XXXOmQhd+aH30SFh7Zj5OkDJVbjGlqtfquKLIPK9PYlfwrklU2OxB
b9t0GtXErL9U9V0Xk6Rxq5pE43wVgWEAgL6d7Md237EEAD2rnJDhmf59VOG2i0Js
RFqQng1L1Spn4Dz7aj/6tTHepJWMAlzq1ncFguSLxVnIQ8bE8G76WxZh079VFyFx
RmpwII3B2z1cdYDRuNTBruR9HgRvp8ieFXzfibNvpakHiI0l5ywVHUL1fpueXohF
KTcuGwZS9HG6Y1lFJ78kH66GUK8WtPsmMyoYM4/M/Rhu+X2ypuAwRN4NmwSXie40
PuCGCiNeDdV72EqU55habomiJzmRli3F50KEh+wLJ6x9UbflDODb7mEjVkDZJwSA
9JumRR5wmqQ3DOK0hyneuhruMgfICzMxUPF8mX1Mqrh3A0FdAS90iYzn8IUYNicl
qnw+miYItRCxM7HUY2ILavXBme25C987OQ//49/TUN6CYODh5ta5uZTmKQR6J/Cs
RlthDhde1xptFuHNSzMqwBGqNAcFA2RlcMMIbO5haWY6/Bv/q2T4vEVi+fTCkRil
bhYNn0fS0C5tOvniIkgQEtgxmo/4AG8pP/7KTkdiBLDdZYfZAKJfrL7SWhAQG+UX
FsMyUKxagRdOULfiz+cddf8FSN3Oh83G5HTLc2GuDXrBqStJtCyKECeOnw7rTJ4h
VZj7SNJmbEcN7VzCjmPhqKMqmLxS+p1cUmMu7JBldGflTvFqQMc6xaWUbp25XgEU
F11LhILHgNpFK+vwaaEzZYvqnJMps/c6V70b2U2AU06qzkmMcqbuw8ukhgIy4hjE
rs0uhyFYwUKQNoZsPBQnq0GsnV2VGZnPIosAomGK/1mayeqIHMTKc9nhgh0IrE91
uyc+/e6rKN+i7C2YaBlTqxRAGei4jk+Vz3/zPA8CmNIRkj5KjHzRYbjPse7L7Btj
ADJRUerbQ6ioEgwqf6L8BQaD6CrAzWcbKRQYKelVi2zF25OZRP6NGWVfaZbB8XZd
uc5Tug6S5zhMl6WWeQXKeS4AgBkjuAUPSWC8R73tHhgF2PMd+x6rEZ88fXHlSY83
gc+rzRwfWvqe2vo7eiD4gpzNFJZGEhk9VsdlwqKDEQsSvdR7ZvAEPLhpZVBJssKR
zvdpgjblyyzJ2oD93/Vi3eZZRPkrj9iqnMmEzEfDj1Q4LOXfVrirnkPFc8tgIbYD
oOiy8ZIlhGAqu4GojuSqhM9NPDm+NogsWXzN0U9zuSpTZAC+9dhmsnCyCvrtRe7a
sOAPizEI2NHGwLieBzFyZH8kFwy4KK9YuxfrT4YJPaq+vVQoPly3Qff7LZPAz3qe
l32JheUuVlxsvRqjI5dg4EG5ShvMBKTx3Mh07bC7wTSWRLmeZVTGmEQb3ornQWea
E1P4oHQYQWvMIqsrT1zYiaHuOWUyorpJvpzSGtZSyakJaTddLupmgN6U63Z16Oe7
HsSnpmMOtImrSyGC69TUX2LOcyLe8Pw/oJ6lT+jnKWdk1glBayYIvWQwCQaOhxDF
KSg12ZjkNpuTG/Dbv4FIoz7LUZWoFLlhG4dkKzuezeGHDUaDGX7bgYteCf2F61mr
b6T/jEwxvr1qg+CrHeaKB1wQk45cbqhU2D5C5AMqdWzQppF2AllpVsYpfHHUdk6H
+LAMFxi+MHecUTQVE8pSK5bzd95WAdVxuCemEXgFpCczFq93/26lT2yXo7+XK+Q5
pWnOh+GiQ+GpSknzmq9BarHJ6RjWtx/jx+0Afq7vbe3ivp8fozHujBy6xg4pqvDM
6TK04LS47LMpvXQUCFdyt0PhEO86GDVJu+TE5ms96tALmHlbvjNgAIQZtFq4uLCX
RaBZTO6oSgT0JAl5SbDLpIzrh/GOONgpazbAxjUFt/L1GgpWoO9XfdcaK3GiUDNt
N+VNHG2xjMxD9D6XyJ10aB38oBBngtXSlycerDgFL7bv0+9Tf8poZo5pYVq1U+Hg
+B18GFNh09rSgAqYmzqF32DMPBUhUuAregWKYpcyAfN/LuRoBaaTHvz1AQNgInQ3
Jhrqu5c53o7BAYYh7tAkeDn6uqRbfA3g6W9+PuAB/oRK6RKAIZy5xPq+mNYUjAkq
ns2A/Y6YAMZs6/HKHlsR0CmWTF/btr9vcsbFfVogkpdOQGCG6NUOa+3/5zG0h6Oy
c1bKuvT504gZ30U2i1ZJRWuPoCisD4tjwoAbdR89c5fpetJnJfnMCi1QVm2fwcfT
cPNo+1QfMkIRyr7wJS4DSUbYkVwoq1NqnEyBz+TP6i98l0KuntQikNCg9VT3Z/XR
pi6kJEW1Hh1bOP0gXqin8fP4kicizc8EFw3tp7DNx6D/jrIXdcOLP8vb1kX2hCNe
BOMFr7hZjSijS9PkceE2lbzrV+Dg++dONtLmyOjqsjOI6hZbdlkm7n8xK9Eihimh
4Tm/v4KKuUTtGvpA/TVyOtOIVCxzdfYwGoz+70pFIA+9yE1teXnSdwo9xS6hWEkK
Lpscx3ZdvMVVH3f369pSh8bs/xezE1IcUN3RSBR1K8FRcEukO3H5j8Jp2QEjHKgs
qxUe70pku8j2IPMhf+NQ9cd4acrmfT/HGmRYOJpN/v5cOjy9surdwHjYLvXS4k1i
yRMy1bx9WwlgAkYx0HuSnPiSo+6GJVWdTFNM+GZ5KWRD1sEEK0emqGXGqWFAAr5F
yRWrZ2UH5t3dM9GpY/PQd4GCe8KfNtf96p9vYbJMol+T0OINs0JNS0nazgK9QoGB
qpJX0oTyNhLknvMS2Ksaxtiu3HQdVkDKhAzT7wVeiV/nDea5e5aJFtvtTgYQx26p
tY7P9LnNzxkC+RV3CfcmWhb0iDpq693mhA7RhFu/5MT5P5cRZnpSR/AWWsmW03dx
XiqP95yDcpzeV/MEDsH5qpr2eNntBFJVpRD0RGRmEqoXM72zVcDZ1sfPbjTSNaGr
BlfmrI6OtUXk/PJHiSemy0/YdQDOan/QRt4T3YSLaAkVsZyJBJrQGrV7baTzrTVx
IXwqBqhDeUZDEPhyFdKDsJPh939kbKAfv+EbCZn6bcV15BeWAX5WOpyzf7cFfBy9
Zc4cBLO7M2Oj8N1/8iVP3THf/FAgHnBkey6RPthXxMQ2U+8XqglvNiOLd4shPwtC
+EP1FJLbzXE61gSAgCU7EMSNmaOy8ti/suQlU6OGCAr+MPx5NF8R/yljzX+3OH9p
R7XQCB1AGg0kZHyA8D6ar+69ZfgBDvhcypo3PrM1GzfxHAJjwVps3yQxoIxNPeoU
VJf4CldGn3UrktGTpxEJRhP3odApidawEHvKdh3cYnXexAiQEtmSz2dUb7ogmP56
hB1RPRkprJ+aa2k1wJ4xd/xplHVNWLNaR4lHwyrQ//L2gwIdvQ3WLj3PHO3c5OZI
wxCADOz8aO/eDiPTO/Bn/xiV1jG92Cgn7iuhdupxYqUh2JFhc71nwWkqczqnd5Mo
N2W+KIzuQyQP/sLVFMhQULGVWaEwdgIB9yGZDMuKO/dmGgqOnQgbo8EQo3BM91Rl
ju+p4gvTBuh4W1H5aH7gvddSaSIJFHyKUfXyku39OFyTj9cIM4MoucAXKDGL0Cjn
3mflRuou0dWVRAb0jtw7vcGY4Q6MAsEgCl77Xmz+422UYzFwtbnRdLscx7sssDKI
Pq+aJny/dWPsZWfh+/KYuCUY24eVJhTRRDiZI1lJYa5RmeJ3zX8zooU5O6RmLAJu
xF/EiDzXgc9XOV+bc22++l3qtTkdQjZPrgbQSho2tdkw5/+lQr/MQJFKX1kCKeRI
bWymLiw5zcrEZ6d9m+BGpjD5H6syFKXW/WQRQEOK/WOSfQzKO/JAQGkg/uEL9cKo
bxIOtDXkj2B1MJu/RJ/2ixa46jPOzdUGW/Am0QWGDYols5BlkLRjONBs3GMTXevH
dJIbKNhgw5BoY+KBSE/b2yPwCoM8PtemmuvRXKS/JDAHcScqJ1f/8W8Tha1Hx6dt
r/35RxZYabbiimjc83gW5XLcv5CCmb6ZgR1U7qiHzhHaeMb2Ejz+7Oj7hR2Q4T2M
MVP047rfHM0LFuyv4CuSVPt/X4Q1kGJG3BmvLHPMp3GVYEZKvCKV2XjuJiJLcB3S
r4/OBSc+Y98bpYEKo5dp91t3sUw2LbSBhqRv1D0psrnD5HBFqfJu5JsoShSMQWYV
JKQ7BISPFxc0Y2O7AQD8TnQ6QLMMd7IeLb5lveS0ktQ+dFPeDcECzTVPvHZLkWky
xiw8O8uXJ5tsdv529eFPdhZuW900OySlSMTPp2z70GjvyruW10Cv/PgkLzY4m3C/
67YojxSJLy18mzz5Vbj0RGY6K6/O4+YcM63BnbZsBTglaTp0ysn+4VUnybUh8fdH
dbFvw8p1VgSFHJZrowh1xn3/snzijTR9X3K0k+Sy2T/lXoFKnweUs7A0G3vtu8Ot
Cj4E5qnG0SA5kZ0g3FyL75h8UsN0guNwViz5rpVMSxfJ+PyxE66SkRBPRbvl5PzR
kIp5Sj0lOyYp7hFPRmaroLVRGmK2TVG6MQ2zWJmOGRwF4LChd4G9xP4t8GwSG0AF
KZ/dM+Bu1WhK4jqeHP2gmTyE9EEYiZIZ0Jhk2uaJBBMO6PL3yhw3fJUSrpoGpsp8
P/58bk+3pSvaroqP3SXIYJ4HdeXUeuLdmc58Rcl7y7reeEuNAz9RHSpCDsAFNMq1
IF/AaNuSqZ9OTVjvpJAHI4rC4KDSVfQF0BE7Uzsy6dgPwRIhKqf0w99o/OIVzh9t
rmb0wFRjv1rV1Ye+iDzR8WXu2dqL4Xi2fUPQiOfVbRWipijJIzkavhR0StiQC8ce
0uphaaPjx2F3acWgcfXdke8AjrRxR/PTQ4v/NdKU63+EEdVPFzCsWniIdkm2Dbxi
8ABmAFWWVMXkjz+7lKpmevF7Lfd5oidMnoYk32wq2C2jubDGiWF8Uc/VlawnvjIg
iqTjGouoVmhqXZzGj2QOtL2Wo+g29emIQ0TrnqwOn9nUqicUOYxGqs1E9S0jKB7k
bjJlcu/GQZG7fFY10kjB17rjiJeq9wYUXZ6GuF2cJre1ExcLhkxudFruijYM64Jw
VNduO98h1Dw83izhfgT7WP35VYASu7nucwccYNyg/ArORVB0tJnXejZCN/KIK/3u
UG7gK9q153BNggHqFu1DVbRruhYOoTfHm0xnIW9faRgxhziBDmg+W3gZIcpHNhGj
/GGNWmN7sESUW5XMnIUMqbrLu8/EIMbEuVJlz+hl+TJjNCjRD1bUQetnkGXrgiOp
FP8eJPbLaaPJhZKNTSaDDR5G2DzB8LJBINfdnK+nWDjtag5gpabbyj7mNA+2r8Iy
eKT4ObBxwirz7kAzGDQ1NnZ9yth38dL2SBxxVTzqkvybWHtRPN/kvgco22gJA8nk
YXry917ArAaC718UY2+CSoopNQko6fmCC9hx55B427Zvh0NFxjNvg00l+1D4ZTUp
xK6er8nftITKgCOoAyvqu9j8PeRMJ1BKanBEJsVkRUGrGuZ1zy/yUF50oZd2qw3e
TjePC562JZ740u2h9cX/OHRQA1mtPTkkbaE4bE787Ovh/S8qyWAgmExRzfITI9QD
5PgdBOmNRaNmWfoO/ZzYETfxRw59V2C+qmcNv7NIl9iJVIzk5fqkJGNmv638sY7S
h7QaOLjhQkPCTcKAJokRwj9AUQQAgaoZITjAm1LCwZkdME1IqKQnKa7b8y4CxWDD
BctT8PEvcqGmc1K4bXgUGFv6K7EmsdWXw+jC4+TjnW3jSLD6nXoG4XFlYUyrfnTv
pNPmGJbb8OBtDS5+HR/2kxm2r17jhsRB1r7trg+e6GO87YxeUXcQpdkCOz6VqcEB
e/W9G1NuicK6fjAWvNScYvgSc90zLlnAf/axmTENb3PCfhs8zzOMkisMMOjANWBi
0yDpJjatJyYx3scjN8MNeudxYt54BmyfrY2v6sqMFPdruTsTDY+XXLUAYtC/tfCD
CePleKPBYinNWFBC5LRmtRfQWxj95dKIMETyJD6cnCu31hZoymEC9ScFyp1SQ4Ay
voD5fFMfN8XgMsw1MwQgB5Ea2WV6ze8RWnAiZQovIYZROscEbWjSlNNXN96NJOmC
c5WZ9bcNXDtga32wTexHwU1+oL/AJwFCzO4xcSWLssusfntXBygMtEUtcpQ3y/5n
+D3okypjwUpBJFS27j7SRLQew40HlSKyOiujC8VEPHSw0cv6QpHBxP6CpHKSaLTE
fFFZS1ZxTHBNWSKTlLLLQU9Huq48BLpEj9J6G2iBOkEi2bBsVwuO/OBorRuBEOeH
rA/x3lzfnZQAR5ZX5eRKKFhL+Hl+R2nT3++Syx5ZDU2pGTCgBh+re1HzgUKftzfk
G5y74rcutgkw/VueOBeBgUy7b9/lp5MT6Y1a01p0DFSDDvTuK2o4UMgRe6zWkXc8
bAxZuxsqhXSDOLMpihqCJn5VNfPJ+IxLemYdCxbIrFd0h/4NtikTtR4EN+OEdTDX
1rVLbAKmnMucQ/MP0mLFGG4Dm2ySzIr7RCoqUr038kskw9P5/vBfFbK6mZMaYLVM
YwQASrPylPZuqXwauNOAb4OidmOz7mOhVUi7xAE6xNlPIFkr5shIyexZxHRtJbGS
cWAAMDn7SKIWxtTThSqSazs9HS6dfawq/kpIG4sHP4j7ZQEotgIcF5F2l8wUPzWG
MB6QHoR8MbVXuB4h0jQQqoxrefwlPXxyi44rOq+lVjnQJw3L0vZanSXDgL+TgCkG
Iq4N00JaZQYLvH6uwoYVw1up5iXAMu0QotuiHKSSzHDSV+AATnJiIcBHXVTfG87J
gYgXFg0zgkevMJiMwsqD75U8WwmDKPIxTG4+4aR26bHpLplht29Sng1XtObA6pU5
/dYEOUHzJJtDIStgsfzDHyFYVMd2YjHNj1W7KJUmDuBJ6YROyNGJYChEveXEij0z
Em3LtBKbETKoqt/XhyVcRoQNU9yEZ7bQDE6Zvmn3Kdv1gAGWKL7vhFBIYu7jkTV8
w1KsIeM/zh+JiK/P9X4qG7xqbo5ju6mBXxQotT4LMYaM5MvQvodwvFjb98FMTxOr
RyTRINqMUA+cJO0tU/znKLeb2eaDfkTj5y8k3Xo5LOpWQsrB6TX6oim1D2GYznlh
AmulmQvnXF53GXgQy/2kfXAlRLNaxn1awRtjDi0TcZR3I26ov5kXWtNcJGlCJiGz
hldo/ohX/ILjtsL9Nr8KzncF9uaDO6g9Mhbwuq3tJz7Cpb26m58TQA8j1SMl1K32
Y9dUy0G4eRxJP1zlWeNWMP53d1SftR1cXrWvwmNSkRLhMeYqFiQUY9nYcdqp83UG
josiPGYLxe/29dgNIWriyaaIfa2RmuV4YNzPA0wOa08MBFR0IV+1ORlm2fvj8oH8
cddQ64jtDSs2A3CLRFR+3BlAArYMB3IjXcGD6jSRci45cbaO3xqcyLb4lFsFCg5S
Yf+V04X4pdb4RWBlou1W6PAPmpDpo37pN+9GxXPGxFxmGj0JCYPl6Sr9ZGJzSy8t
RNh8E/NkZruE+/hWyv/VfatKffi9ZCYVcYnSbBbw+0x0Zt8HZniFi1pv/163tUFc
i1ZpgZuvL6VzKl9j9B7TjQkTm+er1uzUHMeJoQXW/1JwSedRqjUs/ED9t2NzWru8
ylYUZWopP4hAJKBaLIr/aZyCBbVORc5YPhuA2N4jF9Ps3gRpxuddxxkm6eyNKze9
c6Z2rHreLnANrQLeyIPzWSQyDUDmpmjoHmBmj08fuzAf27zlfj5m5rTws3fgv0A4
8wIVG0iQWlI6Of4LukLoQeNfdUMaiGy/Tca1JCuKGh7MmNkraWQUSRM5RZuTfpm6
jzBlVTdBWsBuXjPxzTLErAlIEneS7CUDODSiTF5+IZGT5d2dDPJtVmq7j0rIMass
SQpnWLvd0daShGQ1ELESINaVwQzNLBDETZUrRgdy+psO5M7DIgaFzv5Z+/1do6yi
MQ1UEZINb4u754KKWEba5Sh4n9ACoMhKJeNPMHpwWpskiEH6zgOCmnntM+cSFWjF
mJxjFSpVEBU1CxsNC+NVWkQIHQopt3oPyDZzk9UvIo0rgDaMmKW+1uQdIkO/bmrG
Nk48rMNAqWT+y7u4mdcBxFSbBnrqSWImZYT81F13qYblZnI/1oIbROAUVuGepp3h
E4Z0+TvJj2nmo2G5H2WAVy9CG64SWtPYPLzAW2HW4ewzr+mNnZX6TvBQdrHSCtse
wAT8GXB1UTQkbC/oaaA/hEMUxYCAny3pyxwlgTlhSmmT1xHu7mOUrP6NK78MJmXE
jqSqBqGpkqoNHn2n7Rosdr3+DYUHlJ088P70jDjbjryRkePGUvzBoU0xfJ3VwpoN
Kj8Sg7/NnmOPjxHwILfODdskxlAM1/UJyLXzky6rHshucDv79vHpOGaOK4Ebqw+Z
KSC9TFPLfP7PQntR6QuQSa0F3b/2d0V8WPmslxnAqcm22w2YR7fxaGhk+EnyfeO4
m//zekkhfX6YUmBkBkactkdNEJVNfjvNQVadOZ2WJ/p0VTCgPtXDEdMr+MjKP7tL
RPTEa6FKKcQa16PuyzrULalVhrvSDqKPXoXYDyL8CGTr5yYcxEXnn7K/S6kFIorX
Wv9X8gKScuQ/7lew5Wbmkf5pE3LpsdQppcQZeby+wqjuGc+KhvKXGf4QPghp/WKZ
FSdrtP+4nxmoeP6XHSspuLrbZanj5J8fZWaLJ7FlrnLzOMtDC0+FP8q61vVtwrIV
js/hwF0oZSkO0PFrUCPGC/5b2ghLhqzGeyvUH2uAZzeWsojwr9gfzpax4YBbbR5o
atPNhWRnB2YcmmYLivhX/bmPAW/jMyHBiiPAYdVDTd+Rpwo4AXkvugmBb0YP3pm8
VSiKaL8zsR3qPBQ2x0vJT3oQ+JSo0NZhVPuEpQqjzBRcehEyv9RduwIPA2dGjBr+
0/5E9KQ12HXf5gnf9auGt7OC0JCsIaWM1eSTMDLH4GZN4SZGmk9sqfvHj7i/hcJK
HN7mqz4qQwzCoyPjNU2Oc9tYFVA12ZzbWHCkbr0fabfKOOQKuL8NRM4u1/nlCfsJ
OBu8yi6fIkT/XcgKOgWt9ecT9qrDpJm3NEsBTt9Y5L7sPfdF20XWjPJrc+RjW9gt
1MG8p51trLqTOqGokvaajDZixrfDTkGMnaH7mJxrVQw+qRwMzXzT1d8l8FT23HBX
0qpJLHHSFo7NLoBFY3lezHe6OyXlYZWpS4qrL94kJkxfEAqpHFX4Uv4SHmTFVhZK
gjzVwsqJE2tNkMeF+KUIirR+m4gHYRl41jRL+qpnioMedLvXINjdTWHkBHRcxtDM
l6dAreiAuQj7bQWbODkYzcao24VpL5j4Dm99XlTywpkKJPIhZFNAVDoYu4+4fNya
I571FJommv60KV9pWLa/lQeP42k3vRKns1pOeJXHUXYhrCSWrejjTTN9Jq9ipjhe
M0k0qFUsbTglC39cW/LxB+1uxwfUqopbz8hG5krss6UaMTP9L0AUS55BoxA3tz5V
DyK9VIY2SxHySoZPxAIY4eEZrn514S32VaUikmR0a+qYU7idh1LljsLPpJ2J7+K/
tASENJA5nKnoCF+sFQSE2xVbFtnDHvUx+IsXZRxP0T+Z//dhsPBZOB6NUd7E2Ezh
XAYN1nZhdla6/af0qUqfij8b8LZzcnwxFZClylNlaySGIwegLTjJcLL4BZ7EGMWx
6wQfdMgqGshNgzYNypBBLw3Er6MEaO7ae9jh+kj8koais/rhXdyAwtk5gEBZQN7t
ig9/bZQ6CNdihyay9gxm+cDSnHFcTjOKHzvCAoCK0YOpp5we4aciOmnn9bHLIWkF
q8pnRAcSCLKcJnAzhmtLlQ2NZPo/ItLt0Zh6iG3KsSRbgwsDazdwE9oxC4pcb9/Q
3Bl+pgIDZqnVsTZzFXDolx2F135Xa7Jl2bxs1ZOySX/afJL+ClNk2oAlYdoK4L2A
Hx6924iPaAYXVnMpXWhELU9koWDzCITiIhZELdciVP9LLF0P7CTZyX2165N/KJOd
H+ssKtxgkISD3MSmYVGgR8oQSl05Q3H0IkI2uBbsoKVPFfA6PEnZz9WDIBCBpagn
3C4asZTX6KlCRFwAF8xRLyQ5uC4z80CV/feLHxgyA2eBqFt3e00znkqp2LbcWcx8
ZBFez+ZF2KmLYpQWFGuGfWa2OJ0g/L+JAQqsILD8oihxwwBFYFH38x7zhz3vT+Yy
dT/n7iAu6T2FmsNRDeQVEt14FoyfU2eucUkl5yqNoUf7eahDXLzsxcGD89m34YKa
c2acNEnswKjXMmClyBJSIuFFzvjm2+PsKhBClsCqN1MzVXiv/ZthfaGQ1jKUJgem
RbNhgATuPPpjTbpPc9eR44KCSeJEdxe0rU7VZl4AxH9cy1mamzggalXy8yBxwIa3
ihbTR/6wus1mBbG9McOxkFnopxvp7w+oyT32suB7Bfo2a8hKuQwTliKOhHXkPf1x
uiQkHt5CEtPNcvuOVdzM2XixIPM/IfHAsED2AD/e5PFJJYHNBv1UPkQGNHfvWOGt
EZwoc0mhgNgvpu0CyJx6sHoUdUhCtHgaq6LpJZrPiMqnmPbk3smLdsmJ93YjZosV
IDqMAHN6gCf8ryDHCFNYkDhhgIMAVlCLLsRAvI0BOxAb0mHt07+4M2ThDDCDRXn7
/Ou+yQRvQ87KulEZ+iiIMWFAdKU8nlgf9OOKj1VTNcgPB7jZyo7LP7wxrrweZenI
XRq81S/ts5twaUJQzQyWIT4F4LBSEYJhzydxXODbsVufzcfiMO1A+i0pyIcbWLUw
Ra7OMAJzYYhzgoyfcZmSatRF2dt2udXidJ6C8fqrxKP3Yx5RvmKrczgmyyvkY/zM
XLKQK7RvuS5Zu57vRdgEqixpU9coNiGkOglbyyla4DmV8xnvCEc7gegy1IYRdhQ7
8LwyYNhG4HXuOZsENLdSf+lyuuan1XMJ45bjKhBYHKzxg2HghLxqE3D5CRkfvaaN
/WFGzaMG2jS65EfQo0NwEPh13MwMcA6i+lJyXhdX5mzbjTTLwkMeMgZwTSYoXDDZ
6tNZynRH8DankIiYKUknbmKmMYX6lsG4gbqXNBqydtPnGm7aklGSweW3b2z0vi7K
17h5gvs764/2TrmtNkGBzMsQO/dH7uc00X79D3EaUIitf1d8gUD42lM3cyjl99Jn
p6S2Hk7mK3mGmamIlQ4sAvHpDty33in9Txri2zWKE6Ue9c+/h7+ONTXw1nuY2B03
adjEYZOkaX1Trc9ay3MmQsrlNhPoLq2s2XmdFg59FgrtepKeBmhk5MAeP1LMocyl
Osl+H37VEo1juIOlabv6U+0jAC12C3QnpOGxetfgh8SA+odJCgec+lj9D10xRQzK
ts/X/pfCyzcxWeB67mf4PRBfiHKxbDnB9/QC5vC0mQL8OC2U5LL2LeJDZVc5cRMH
9SHyAFAWQBMeM22pgqf45N2Y+IKPCXEjRhnQ8EmuB1QWJPe6kL+6l2OR2I3oTym/
HZQQe0LDTMTCnp3tY1fBudzjBV1OW+zJGpHpd84aDLXrk4jHKz5BzfNkqHaymnS6
wRDu8YwTARlUjrmnK+rmaM6wvgU9hIehSNXORCQH4IkHZNwtn8ee4mUQ5e5+U7r6
j9B66A6ATHbvAOgkqxRrkNuHtFtIjpTaRUGbbLwl473QHfGlWitfAtuMPGmeb0WY
vja9CmTzmZhA2d37G0nwaCy+/IdkI1w2A2LDL3gOenQAQAmStotmhHXSGGMWHREw
CfPf30obHy7Vvzzk9fw10b9SiC2J8iDM/OyL2Lb7059KHtgacA/Gc2RL5KiQirve
bijVneSIpAS5MifXAzK6biwqe2QFMOK6bSft60Jv/Yl/in6fftpLMvzZjzd02lU5
vvkl9T1DbnMyNv/PTy0dxg5Q73zAoOvQNUK8W8y2OsEKJPfeaPXdFkABc3MZqW8t
GzP2MbCcjtexb+Le0Cd3zHVLfClhkb5Pn3PeRxFGzvbATFijH2x904IEMdqxazv+
1Mrxi4ogPYfEQuVQ+A/PGYWM2nPmvVxbGXrXcBOWXUHlUXg/ALfbsbfctcsNB7HG
BGb//mUodi2j9IiYZ/g4tf5sOh9Gzg/CED13o3Jsa9GoXYJgIK5PYbe9wwjx0tVX
KveE4ayOZADoPgXkfxsSWVIA+jgNm90PbkWAIjdy00tzGGRmMea1uOdegQ/KaVaV
Gf5gXOrHNlo57msLo7PakzeEsXW3jtjTtmD60Dg4Hnkbq2i+WgvbmdMo1AR+KYHU
DZgGX4J17G8gmNGHZzTTHBFC5JNM7xqikbNQXTc3LinZFDncDx0GMY7/TA/Bkx49
AJqY7jzO66kvVJbxUGtDceHaM+K3YdbszwAM8L1eE2KjQa0XmRExE4R9y6bz7Z4+
Yoc9S1XmX2CI48RgHnGhQJfGyiMNcEDE/SXxR1SsoQ7s4n5CS5uhCTD2dHtXG044
A9nfxo6nGgVLfRBTm/idknfp7sX7LuM+G0PsYWfoHbGwGjwJpjmrFXQNpoAMdjGL
p97+c5CrUMtPyGpj42ABUFjyTHN9c+2g4nzWfFl/lpg/2K4/E+So9lvtDEYHllEc
1+/EHAG+WIDgR9rDyxKylYxmqGRmar5BhDK/Z8iyFhWspoN+CzJmSJAOsuH8IZCG
M1rPaeW6BHKc/9Ip9y2ElIQYR0Yj4DuQRHUeOohbqT22KBiEX8OUd9I2Llb7gbFo
+SvwqCGGNKYY3wWhRpeWYFQT35nKtj0UO2ly7hPAXzeIY8U6jVGzCarrQ0qnZ1+O
CWPtlLowinyATvu1KD+Ng8Z5HmAxtPOuWz2CDAu5uyyyRPtQLLR688mDjuGbaTr9
ejXA6Tdj8hIIBxho9VsnANc+j0xXMYRdEqa3Kdj3fg3BsQbiLhPbVNd1FX+RA4lY
gWhqCjQMHfTtyVkluYKkz25hAzQotM9B5gUg258d6Nl2gcxG4WshQ9NXvBnb/YP5
G/h3+rU5lIbi1V+TNs/s9E9GGamVxNZ0X8C6oZQH+ojw41HMOzpE1oissC/UmBEG
X4WDZFDfccuNbKgBx5edlfvGQSF9/xUr2Y266ScdgLgKf0mF/hwZuCVhFK47DUuR
AwieBe5vU15ajUMwKyZa4GOspyTDRdPVgfG2gNjxEN2mmld4/WskAxPEePicAhG5
gvvbcv/wGe8QwpLfLoLoHwhVDDckFLfdHGB7hOzoRRqnXNB2fpCtnhXGqtNnbSt+
sU3KZ+xjTD153sEmtYShG9KOY7IA2/ZAt4OaSD5YrgUC6y13yXXX8HbbRZBR/t0e
UM1jzeJpANH2BJuA5GCObTjBT8Td9pMU/osMZK6u9mPL84XR+UiQQAYxklPvS9Fj
wbyaBsRBYVJlqmTfhYVxzleqeb4s3TqW9BKJXS5aUIBULDY3zqMPnFvyUTRspHd0
3REoz9uUwyJmyOpsajygnrMCy6L7n9S13CQ+pe0Q/BjhwaXGgL2jbFXoM+FX7gxJ
gioILOfmDX4w5Dv2v5/zPdMKhL4xV+jMbdJb9HCRmLMh+hrZuqwe8VqqxFXoTe9U
notWbES3vVvRVfmN0QSgHXj4nV3CtbZGqfGYd2qdz+wb3uVJs+jJ4jNKZmAI/Pn6
v0iZIJvaWUB62Rw39OF4vi5zDdJ7KmTYLkYfLFelHnvQ6eDVOQ02xccBu9Bf++qU
STVDbk31UhMWZRSYAJ2pdt+FI6KfovDQx9mfCtHLVlfwK7EU3n34Z1xiYLcSYE8r
iYB7z78rhp4EL67y5CjE8Pi+3dTmV8VkSeM99QizNJ5yoYE9b6l89kWSKbbwXcuE
EnvwYWreEkteR+sjkcVW/+FLCsbpZ+Yq7cZcWCqr87MZdaY3VxS+UDNhMRe1Me9M
7UQ3XfGrXEq0Uj8DmABdmWcE/Ickvrd/z5CQIz/43tUhx6s7CaBkk0gC3eXzWjNq
94M5WFMUoKEf6rdn0/X5KC8yD0DhDNztaVdUmYOKHRnPh/zgClZ+5UL/98PwOk7H
TLALh8uUq2/iK7mOjf4iiAkVH23hD9PGG/ey9j+W0DcfP7vgzAKZm4vc6N8Wm9Nw
F4zmcyablwQTfRBgcdznh5Li8xy52RKzqquKfM48D6flnGIZSsyT9evWWNToE+gZ
qxsXwu7offrREopX3SPzLQn22JTEvtO5FMoeYs5rot1mLfsijvVI+rjeYG4vnvVo
xusECqv8D5gjrZ5idj+ueGh6VCCr3nuUCYscowGMDK+mvOJmwNAcn/beziZbMoHs
mowFESPU9xB1vbLYWNiNwO7iT182aCzlFIexYbc/p3tPdxoEdBGJRl4B58wwRCBL
ENlvsjIOCCHvaTPSV14W31i6qXwcR0QoEBvk08d/+K456rUl4CbaSgiVekCU7UUq
f0ykIQXKu5MAoiP5O5XorUhtIthWKdE758PM/Wk5/f+57vu1QMEquHN/cGOJjsdB
BB/2j+3cfN7vi2Grmb4worbZiy85BrkEBa7kyyrRLxfoidDsZMq4Vu9eSqZgsO8U
1iftS4h96DVa8e/PKmbO6Yps7O9Q72E6ItXzoPqsO7fbmdXhbw5jTBMeQosYFaoG
FRMRTKJftmv+LjXn4RtcFNqUIDU4A8bgd5x0YtlNyE0i61Ppzr19rAlD1E5Sp6b2
DUCueseGBFa4zds+E0PVYMIifQBJ0TYEauC3/YGx6ZqZqUw/O14d4rJO7TxwL8EU
BNwvXWD6m3aTENG6vWagotBMyWdGa4Xk93Cfnklam4/2YavfxlLCYf2YfHB6wUa1
M3zmnJhXapay6e6rTJ56znGXoZeTFv73oP9wYVViUxD0AHsxyEDG4rbE1j40mkN/
s91P85pOM88V9lL+8c83xkhFxtxQg6KkOuID1IyTkORXiIvjz6mzkS17mYwzd5kl
LqNsMWhgr+WvgmGlp8UVVrHB2gi6fm3en8fLxuyFgqesPsm0uXrcZ/g+pct9NgXg
OVg89vVI9YxxjdRE867cgtv2y3JyzWVZMFqhhzjx+v1IwdGtk/xn5MvNQnkAFFXM
1Y9PuG7gTeOTWubCwPuu2iNbcRrTQ1Wt42w1YERJF4b1Qt7RUIOClHIKD+AAvjFl
YSAG9MdDQsXpgAcZf677UtxzM1TO7HsIgR2vos0gLh6+7PeGj279NDQimNGDVBM6
+KCimo2geQVS+WfHmY1zPABdYu3xKwsmaj7NTBsIpGyAeG2NUN1b2n/HwdY5Nvy5
fL3SEczo5ngBry20YJSKJ+RtKlYPn4CapZeQYUDgpGiIvojRzRnhnEX3k47x1Ydb
YOXZ9TRnTTIBT6myTavyqq7u8snqPL0pixIKDvgxD3ecdwAAPke/rjz2gBQ7q80F
jaBiLIUVkh87lhRZ6XLNMN1M7g2k9twLe7SaWWV+8bcStBoUFFsSWoP4Bpw40GuM
zkEsRZzOJiSUadJG32QUStq0ng/Kxf6xp7IX0z4jDGZy+Vu/j0WXnQbihYm7huRY
Nq2okSm55H/kjX0TqpRPhQtZWKNBrCjAHy9LrQsm+IdTipgmbmyhyer+81taZWBT
xGeWNJP4DJ+XF0L1e/6yITlOPYDNBIAh4ZNoO+Dujl10vI4x549Q1JWTO1dBFFkl
UhYgM8D+3DEaYLdIYIHWE+1Nl7g2Tt3zNghobm661RqfhAG1eB0EGrivjlUmXgr7
dQy+F4ffKg6UgKOywAr6BnaYIgvorHejLiFPzNI76oHzoNYEI7lUUp/YhVNZ6GDw
fbQgu5y3cph23fGSufbpGZ4oCcrRlti45snKPtPmAVgrtmiz1DtGNeM1rnA6vdL+
YMloyElXg0b2GlnLCUiinLq9o5tw+tgQHyTOO1C07HdbkMnVxpAC1zXbbb/7+uxs
1L+zmGGcycILJcInZoLpTNne5+rEq0CVxAy4D1lTDdxKYf2HbjWeUcsi3UpIl2Q5
m0oBcVJPLXbwGn4pINf5g5KNMf1NpEbI9IpnJqvO511ckXqqUCmZUPZd5bu6aup4
z/rU9jcbcM1q8A7Qh0hZE5R0I3qerRy/Wd3e5htCvWpJrBsW4iGiG5r33WF1w4T+
VHlvkUHk/v3FnQWykvpTEEdrX3kphT4VPWhWVcpKtU5X4iOl0XHjXp0L2XDOng7n
af5NSK+BJrDyx64/qEbYloIkuErzyJhM+87q5xOKv3XIp2k866utAaQe8Bp3+Xbz
2wYSYVweSfjaZkl3bfmj9GFUPbnL2Q9PhNcyYmRuX6EAD28vrHag4fQO4Sm68EiB
GUTxj8tnTu0rRMuskMvgl+6xvljiQ6mr8NUeYSYtibZpt+vyWFT2Fv3cUh0Jqy33
CGBR0rQcenwSnA8x52Aj8Yyr+Wcb1FGS4PsOVyESF6MrXtzE3oqV4/hXeUAHsp7G
BfWFQet/6MA8/r+CEQw3F6YnIA3F5NYtQ24phFjlpbIatqe7VL47XeKMJyOoX4II
Z+CXF+XgUW4SSbBSYRzEwBPOAGpphaJTRVfUF556zK43yS93AwSGDgRT3s5JaZEE
MS/DIjqQhhC+smlV2hX4KOwQ1ZL5C/4KVRWz8mkBccMlMbdMHDecSYAgeXdPPLPs
EhO7je/Nes4nd3l5ub7eWhgLiNhop/a47PTjRv06CSSKuF1yqmlvMrdxQ0uG6PQx
ImpW7KAiWqGyBkr818ghMlrWI4FZl6oqslnTdu0yVpNaE4zBsHUVckPpr+NYyri9
0yzQK1BGzPllzNqaj5EipWajARl3atdu6fdYpqRDZzyFe2C0852Frp+zeFLnDEpp
EFZMixVLPzCnKLUO7tPIC5MQ0xvaZIZVleel8If+r99H2iJRLY6pELQ0v1VzO1Ip
QZ3PfuHB0oZfKcK8Hv6K4PH0dWiXUpm6+GJVh7elfIE7wMU6jhiPRUBITYRiO9AK
eQABmDnpFTI15Szj9VOE6ANdeAisu1LVRRT/DV3ZS0b7+pABlFuyynnxpYHMweQd
aCElNnzllgGXr093wKAtGZCzA8SkZvXO+BNnQpp0BZBnfKH5pPG9NmM85+fPW/bA
7C332F7OYSVayn8O7Rxh9iJ5XKdjT3WSzksusmly9pIEmDwn3fLwDpApQ9xq9mRb
niwYhSS8mu3ERkxinLPswHuQiJN6PW2sMYEo/R7ezlhJvquzZbfWeRcPB45rZZpW
Vsf6TlNpzCKIyTbaJ7aCEw+cvTTRvwr8n4tKo7BoWldJzzNWzeYb+Eru/1Um2L8q
DudoJrw6UWawLsoGavdFe3uMvmtnPjeaQXhcmFWMHLoWQfPgWHLNyvV3+oEr7clz
d6SJtokGnz20zMaErZ1cZrgYHsp11qIIe8SzgYOs+uRPd6yTuGPFaPucG/pLDtFY
g96Fgyivck3o+sHrGZtfMNd5hecg30ZZRGvj3txMqHakt+dFTcZtOuZGozFpqdw7
cZCFrOigBh8flPTIkIWnFpmqTb7kv9z80M6MQVdjHK9ZV8vdV9Bb0dyWF9h7v6g5
v8DibYJ94bVc3qFgnN/UTaPG0Gp2lwwiW4aHY9f7wZt25ffOqKa/h1+nU2hqyG1I
8UQcmlsEHSJvwwieCDl5YsjrRjH3kK5H27bDYKBaWUlRAmZLp3PRp1Avh7oTvXvb
A6+0s6rlzc9I4yGRgN5eC6xFUMiN+CVRAb38H+6IfopUJ2+3LOYwy6JeCNKdOT63
f6NZ4eu14Qg3US78WIreWeMahTujU8vFOJ74lce15DTH2cFV9ad6tejQ386+qnt1
GSWuCd879yKe/uhcdPeISNdFJ19gLzni4CrKBg3ubOeNISb9UtIJEDsKhf8ap3lm
KAWAfKx5vsjt4BypZblhXV7BJTyb+/haZs0LDU9XeuhvnLqsPI7QzBaCos/4n/Tg
xmoNUBtUQ9eoT+REkJBM1BH70j2urtWSEnAJQSVSdRACGpqa6LF6DagjBzCLW16e
f0JsCnUEOLDW85PirDzUQCueYJthqIbVsDNvjsfkD1KFcXtRxgudEIw+5G4Q4jwx
4Y/1pJOF42tmWMEISkXE/ABqW70ep0kQCepqT4FjfgJB81JRvTVjpO0HIdyiJN9U
/rUYKASHyoy8cLsEFMEEVHlLrtomkn2FYQcNN+Tkup77PvIl1KYnInDqZS6GT1GA
X4KUXibtcKwOMBYCpqFJOrbYvKTksueN8W+/fnnGFasr9Lwd5MCsFVEm3un+H7T0
LJLFEQo7LXuyeYjw1iuPkDd8hmOihoNOTTGa0L2wOFAkOz23SeQmwwgnp/k7Ez98
RXOPfxQAX7dKxUCPJuH+mnUSKW7DryE5ZnXYIP0eOGjk9YIlI1hBMV4peJZ9vTE5
h9IG+GAh8F18uqNSOZpcedXHPTLwCqzF03OwJeOAfDTjAg/knS3ItstJQckykxTQ
BrqlEsz0xo+kfzLqv891xjW6Bs89cvhDVOBguYNEM0QiTrqRhnDqfHFbWKD3YAn5
liJWi8CNkSRj1SoFVCdTlNpNweiOX8hbR3EQl9qvodPPWPpAzVMW839qyqHmxzn5
r1BL0nJGcAohHCU57OFxLnRh6rGPRM7fPKnwiQ3XpwZoTZVQWtI+NR2bTF1sAN1W
XAMsWGhcaax02mnv8q2SZYD1XewhF5JYNF4ZbkESldvhNVvugij7vfWaFcTEPBTP
SaCn1w0Ungn4WKHWBi/MEbusMznsbGzvD3UyrlIRqyp0Nrc5LjPVerYPPk0QisI+
4t/w1BFAB3GYIb2C7d7o/1f1XcSSeXcnG8O0DPo0M4DeFhkW5P4XxYOoNTa9Em0C
XVtxJHHysV+2WvSoyXUiM3I42CJlfPn/VwJR/uIyQL4CkzaScqc/iKLoJL/bs6UA
ilZKThSMoRay2vEsvg4n2gBRsqSwHkTBpiWf7xVEinol3uZDb/dgZmbfQQkcX6VN
hWvBL6v5JmoWyCPdCofK9n7OcqRCVRcrLJ4nMCXEWfcDVAQ4JRyFDjvUBOxmvWRV
8bVuKjAoRTiuD70mX+8ClhJ29e8+xQeMCjLFTTjOIkRNfi6yD8uhBTu0B694WKIw
DcItQ0awe2gGpeULenAqhgJ6luw0UU7RWqM57vqGqMoqtgz2qojW0ysaHQhjyJl0
Nc4PDMKxbhwABkWe7+sn4mLzHwrovdopSnE6x26O22neFFquIv0/H0QMvJcR7h86
7PJimWEYTb92FyBum6nir5woUboDwuOH13/Ydfl4E3JOsyP3qfj0NM5KzLkqWPB1
LZCHTCiSlIEk2CVVKMNdUXIeXrT+sWDaSCtnldmo8KlACwYojT8dFY6vaUkidz8O
hvkY1ZXPr9RIWkI7kFDAajn5KYdeD3n4GOt9TavxICJAUxOmL/rYsG+6fif2arRS
k5ugW3cPAhTXGf253gqV+6sKRcFrK4xy4XZycPoSpicSlHTlFe6zcImSLX1NpRLf
fitl+JUbZWgAff0RrTmzt7UcMwnjKt3j+PWsjYppR1CP0iO7DnCuxwZOAsTxhKuJ
E+ZAqnTgUEjg9Uq+gt26mD3evzMMXpD+KAAgetO5srvFqlI0ULYh4J7U1ZX0DBMK
atJ61dqg0PyPqEGRR6PLegJyZOvkaZq5Ilm/7gv21lQ4GLlHB5rBXC8MiueztecM
MXwPHQzcVq7sw4JRfQAbIUMOiY9N29+x9aq0MTofyiK9jGAxII7zsh2/dDa7jpSF
9O/QD70XlEHrcj+ebuOv9rZHLFpIMzgvu9gr7hQ2xaEnftD1NmCpmJbhN5s1te26
9Xy+52bg2AFl7LYlTX0bRpbzpNXBXU9j7ADZbzU1NB3gGAifZgxH3elz8FG0PnOU
BnaZrQkOGIKgbqFuvcD52EyMzUBcELhobulB7GsDX0SabXqRu98qZyyYeU99JFcV
N1HPmjUcCa3eIIo0Kjpy1LVlURdvLF3ppxpkAWg8ZkIQHtPOhCRD5gTVyF0mt3Er
7l1LT3rhyecJF+5GkQLsAtJ7HLGbgcuQX9qNj5WaJi44MmDuSlutV4FGZO/f1ZAw
MIpZItEO6z4tM0yXseElRrHmrGYowWrfDkBALgfbcnKwvgMV9hn5al41WztLIVHO
94C2Im71L/T/XAaKSr1ajwjSshnwdJwKtgsC/X2wosnhDajlPYQYnoccjVWHLEi7
HL5ShzCnuEREf+bFI3CB+ClPlDOZbOixu/sD3jhBfhZd14CUe2HJJ3KNM4xu8+W3
7SDBtxF1z+UN9a6Ep5fXnLgg2CgUGjAkEuwd0bFPhyKNZ+2QzB3SICHhVY78hd2O
x6dgMFvOvtUVscAYJnjEZfwVF5QQgsVkztFULEhT+Vf6q5CqhoPobn0AxXAPpKhK
RyTFjAn/sRaEsh9jG0wb0+fZNByctZVzqUkiPS5mEQ+x9SafjGss0rmOsL4jgmLs
IFHTrx2GdhPplRDdCbWuD/Khowt14h6E8fIKQWYaOvbhYFEgGsgzC6/gn+MzuIZJ
TJP+aq97wJKi66tytJ53yYjM4733f8y4GIoTtlnStbuIe8N9uoSqZlg7sN8Idwc8
7pYPKxA7+NQXH8k5Y0H41aYwLqAym+aV/LQhvNO73uZzbJQuVofZICQkfevj9uSw
B10l6rTsPHRuKEK/g5zWR1E/E9DYm8EAXhF/fu3y/jXXU+BkomClFMbsv95hJ7To
8jdZSaENwDD7jVKEyeghFovQt/0MHAyDCd9+ge94YkxsjqjNBUC8TWnIetzvelYR
2Dhahc2YyTaz4akrjGaf8+gUzpyKZlFfaJRymoZl9ELAmOi5zeA/oIWjrOrkmtEw
GcDi2xHW4Np+uME/XL+aSjYEXuFQkacP1UUFDj4fgdEMJ3S1xOMo6KqPRhLj4B5c
kjyHhGZvCz90zE5VQ/Oc6z5rGRDkS5T+bx/bIVKcyxZAbUiA2ZjK7mAlkQ88a7r+
dNaB/JxzCWcJ1Q01vrPgVp0UCRtFpPTTr3mkMbqusgYdKdxS3S3sTkwsD8/BIeXr
/Udv2ibeQxpg2MFuHwiF+1ZbmMlpbh6nap07y/Akr8XkHqsWs200jPZR4VOXvq3m
YpVLYhLVvuYDvIvD6Kh/3uB/EGW5g3gxIcRCY10sR57ej/gN0hEdpdHUkjxhwAKG
GslByg3E3YItlvfqVvwFpG/AJUUatzAz+/+aeJ2j05n58DvKkZMGkM5afXvAmHh7
40GTYqnbST0FdAup4Tj+LqWTYO59+/X78XchtkdDTQMIH8/OwGXDgyavfXjJ+I5i
DyhBJmdcUoZzozhv8KlK68D6wMSJjKOhBIL3F3CJQPIg2h81Hzc2FncPuCdST9Tu
+fClwvRUrItx4P2hu/kvGiZvvfp3N2V0jgkoBjlGWI+bN9uD3/Z/WTwS1f4Ew+AB
lfRcU+Yxc5mQGUECQnaBtgVQqJ58QXg99SdMZFaOnzPkL8W5lwoeIP4SMKrm0SSq
/08dDRlEPzppS3/LiSTNBTJ0OwLohp/98T5421LKazlsYI5MYrNhWzY0VfBCKPJ+
1kO4GxyaT3QwbMcbnltm+ngD0AYI8UQX6n2GhCcFcoGbkPrW1aTGXKs7DrMgOUUp
LbzH/uCUe7lKIpbviMUl5TbD+26bJ6DOlibu4e46sAPc+s+3EypIbss85gSsPR3M
4HdxW4pyIBhRiYUYxdqiflbbgsgrqh7Z78z9R+THpEs+7998ruNgI+ZYCCBRt5MZ
ykde8W9ThHN/bL1i6u2IAhXRcugi8FKGmp86c2TXhcB3/uG+X+v2FHqOEjuvzJuK
IHASQVgp3jcxGI+07jXT6+95JBjBjpPXomSXa4LnUZg2zIC5GgifJFoRr/aE/NMV
rX1TiFeYmmvYxI9t9oB6bJnQ2sVnRbN/hLTAlh4mXLWfHN1ECbP5AQ/wvNbuNft8
3fGXuSaZQ/lPqsoIOZSHkVXJ033ywg11V8fwjezQ+ETTgjLRNrMJa3fN5dCkaQgB
HPZIXSLEsaAStG0BgLHpr215CKNapRi9w2yS6tHLrQ8SsCHXtSjeNPpbjqUaYt2/
9VF1VZgd3RIRgefvlZIYcu/Y+NHhxxD7v4hgYtbDfVtnzCEd85YPYnF5wr38PkM8
F7PIsfeaVdvlRfqBmNeTT8tQg4RCQmEDBnBNBXD0YoODDgiZiBp24dS9toizK1Nb
ETep97RC/JLc7+KXJSMXFOXb5TiVqtmshqG9rQXyslA2/KvxNgh/JHALTrk/6nlS
7PRUiSyuNcBlCQdvKdOL7vlrob4h0Or4O+W3XvPZTvaa5uLpp/s5UrmCVf8vgRBW
bBWs6mEsKklqUkwGIwbvfsSmPlQ7tXUylO3Rme4dtluJb9g/Zvegc6szVWc4Y/N6
omT/rpBg5A78fQbnpQUIyhJuQwA17gqc8lDCsxK2OEW8ZdqU0c+NDrrky7DFCg9w
Win+XWcUUeFfcpJ9ONnsnFQhfUybpqMRVfQomZRjU+qPprZD7gZWdRNX/6t91a1U
Lssq/o4rRUKDrYGuWtx5PyGWj4J+MHB/zNjh+nDtzOmwBJjpr5cbH7+r4i8opsVo
MuUO8C8tDh7gYFN3DtVFK2y4FedzRUn0VOSTyXKHwStFIGz938gJk+/JRWvB1GuK
WirtefrLLHh/mC/Rn9t/KqcmrMcDwYTaxQMPsDmvaTipMyNdE6eUQqcuojjpePbo
gcrnVIlAFv7FsffxqvaNQ+eASCglNRPDjOZkc+Ef9basHfiJ5O9cN/v8jdz4Fvp0
UKmzH0Ko9dYS4I4HADHKYg4iARr/dbxt3RP/eNobe/r6FHqFRl1LHs+hkxO0E5KN
H6IysheR5ck0L6LrKCm7/f+kXHl89abvYbmHC5SuzEVoYwuA/7IIXmhqloCOkLER
rmKW75EYZTAo3n9qpvUAmYtF4YGLYejZjfdYvnkwo1j8tPAjbZGlv+flpVrsbDLb
INp80ujGkbuL8t2j9707jKge/VyezrEO8FZnOm/EuZyIMogFpTPqvv/60pwdwUIp
lO/PreEnWnfMmIIFKm00frFIvuXLH+rpIz+VtRyIHZnQ5n5X4d3+Gf4zN6t6lGbd
2QhwFpr8B8ah2LqOpSWIjmCK253Staj3ihC2gmBvgsL/Rr6szL5uYQ+oCNbTIkVL
ml3t9zsVNSyOrobAbiD6Sa+mEpiUefSqoj2/B2e8np0/3h/zLcU0iR0HhvHifgv2
+bdYbmUmaowc/Eaoh4lXLh2/XeZJd12aMXE7By2pVo+fg3csEmd+tv1m7i+sZhDS
WKjVbRbIEbKujKNkD5RDuH/R/Fh8g4vtMOUkl8wytF5oHgkqYWQEBwnhY+jwMGr7
IubWPrjHPUUZBTvfTbJZkXPwJFdwWmSF3X+KAWd4qZXhLlPkv6KrllZF5M4VgfdJ
foysPdGqOxpfsiTUMNg8ZE4jD2BsHizKU4ZBEmVrSSlzVjsi+dSC2oGdNAFFswXh
EDl/pGX4mNoEunxLOarl+D/xCkQixc3GFBsVrb8siEF0wzvvJYprx0tpvNnDpu8q
XwNc5RmtV4jBfXZGLTOBtbnzkwCo6jihnRZF7i8a4mmlAR2wWQlrgnkb/caH5mAk
gNMy4SEl16jtTG2KC9yVDgtRu4mAb0VJ0fg1Uhvhqyt462cAtdpGz3o75+0HUnGZ
NmecB1naSD1+mcwfZWNyRJIwWqZOjlgzSYKBTIR5QaEVOP75XoSCX2QSe92QntBX
Q1UifDjbBEzdw9rZMAN44I4rlN456NHMY/hdRc4FxLBQPWixgcWcFI9I/G/oDaUU
uywtlPSXrjdI0zVIyOCZVJAbvbm3pXejeZCZ8T+hF3Mo7JKSdeMJODL99kOjQMFS
AEPuZUJDw6rXzy2T8NIs/J+5Dub+O6Ni9PdaCIF8TxPWxfynOMEq0kVIQ37iuHEk
dDYzXrhdxFkBs05iwtP/iI6FFj25tmdvrDO6H+EL2cbjRNHK+f762vf4BgjAJQ0e
DlUz2nDdmKCWWxwDlmE41ZHWFC8i+sMtdK+oerCeldl7LGN0mB1DMAiKNzdkXYyf
T9ex83s1ycCnhXf1UT6q9oid7VCIT12WnTM8C7OwbUIbkODIvZlqNl2W2JwFfqMp
tdHBv0tdiQHGH3Vl5S3cny/k5i6r4lllwqQRQNw8rQnOXpdZlFkY1VvP5ovy1nrZ
9bYnoZUjUqznV375Y6RpH8tzbtonvmDOdzzT8ekMUlvxLgdaC0xQX7KImmMWCQV7
+JOcKrhcJXxH3iqezQKETOlE/MefLJrRAT3Q3Cb2XfIeiwsz1FtPkUo8vCq1ziN+
pN7f6p5+XCvMg0aCpCg03vMdnkZ559BdhRcCm2xHZOBhj2XlytI9nYzUzIyiCxDv
9XfSG35jx70OuLQHCpEC3M/2RQbQZJKaTZSFvp7M5977KwEGSS/xOWlOyGwy+T29
aaMiDGLBw9opKukftTY/23ttfh/Y0pxE1QfOtVkeDmhKkz12Fo7XMWuI5K/wrSiW
RkpkA5sEgr+zh8IgZll2SuBWvcOSEEGj4DoHxeiFNJ53g3eSoSLyI2r2INJCJ7Lm
EovqVJOCj5fju7dxbl044U0mEXLBtNncVNhTAyZe8ZB45gyfpRekEYX1CsE/+7yI
m3ZJbd9uBS/60jUqGJYYxeExLyk/qL5Lfsl10U71ZGvbKdsWSCdJnCq37qMxIMfV
nHP5Y1/pzzNsAUNJdC/3l0lV6Di3jFOV7ZZlpg37chgOQr9o8Zz0jy/2PxpR/MbK
YjOV0TUUeFTLy/ZdYcUEaBmbc71W4X4/8nJK8ye/u1Ai6qhQ3UXOpBDQbOtZ+dgk
L/Cb3gEDGheLWZZGzoDo9l5aosSAtkphz8wFCZQaFH2DVBiSqgQe7QbGeA+LCwcv
UjmHv1EThqlkVlYy2KgY21dq5ISCT29q++oJqTYjR6vB/J/gSK7P5uDfNwFBmFMQ
j4kMX3DY8/JQkUYkHSHK7J6rR1F+bzOdawaKgm0Vr/nojT+iDq06nhMirMBlXBRg
wvcCGSL3QUVBjml9782PtkUIvzz9aUxdV7q8yP/NtI5cio0Y7wh2Xa1yYBh63LK9
HpvbfLwrb6XgO8wopEqUKzOyi4ekK3tjk0ibZK26tT5SRVWppnDOPmd1nx+jpd6L
TCFzj8MkXZNKgePDNaGZHEUxRJmEw8X/A05lgbq1dOnjIzaN651pvB8fGbDbQdhY
3b7OquBNFe8vJBxNNFsYz9Pju0iE3Bew5kS3PE516UuDt3qNHZHXH/zCU04SpCRp
5G3vZiUTQHlKF9TTWGyLlMuG6Aq24ZPYR27tkcN6vHWt3TyOMLqe71UuYXcMUGqJ
YoPpr4Hrex+BSjUDi3z/POYp1tpU0ruYWHW3X7lqhKFuV/4QX2f960rGgbdFTxqq
B8ZQ09Q6jSIZr4knr/T6Z4QZYIitt5urITgdrtgcsl3ZfsM/aVpOU0iwZEZHZCP0
V0vSRG34pbU6TwtXOHXIXx2jsGhF2EKR0nOcwx7fSuloovGQhYs4Chb1f+mJ8uPf
2pRvUROSwxIERU4CyYVaRh81kUHy5qo5XU9FcBtkmqPy26/IzFfdIINtxh+RACDp
KC709fstV0krLzCh5p9jJapBuKZN9yqVtkCpVpZ07stkEnJkZs/XfcJ3qLy70IXQ
cZxIoJ3Kh5VqZ78uh6erYn14qt4uvz2Tcmx4/QWZauLW9NoLLb0YUhqGtAXkDp+W
COjoUFJovfwXHWTUu0VaIsdSSBSMQOcLKEwotY/YA0PKd6VNaPL1UDveu4FCSf/Y
eVQWe653Av2vrB5ukvaV/pEAYayCTEasE1eJvT1Ujf/V+fDO5R3WjJmz41RS7yI8
vel4HMaC66yB4JjI8R5F76hKbV/nZa0LB7SU1d8La/NxObX9VjXJ4c7UFm4dRyeg
dRFT7yJ/dZFr+uWTXbrDEWNKdBuKJj3IzHtlMsamBEAtS8OMFQhbHl2xq0u3zaZ2
sTwqlVc1eeTtxWfWV94YZLePYYkd8/S5p0aXgvHgvBdlju5He5zlnlWZXgnKF/58
xPPEQ9DpOJtWm6m1cJ3DsGX+b5PXR6KKFnMauw+ZxgyjNPcwsybKSqth+YGNVZZd
OjxnMfaxhADh4JiEShYc31ccYZ+gYOHKrTsi0VYVAOEmFSI4772ErBjRsuZ4T4MB
aEO/X4mOM0yfXoDgRWejuUGajpFuW9dAJ8vehM8UhHtjIfpu3c0dpd6LPxWORWP4
J84ciq8YEhV+6ymjMXjnhVv/k5RSwVWpsB3mh51IeodIZ0gmfM2lWDsGTS5Us0Wl
0mzNyeYC7K8w7POjvYqxbTd6hIpU43kHGiURyEBbymEeFGJrrP7jzM90iUWA6Olh
UpRsLOr5fmbC7iR6lbsJTZB3exfMOFZ9qi75Fc/yf30ZkTuJEsRmYnpn0X0G55XA
aksamqXkWMKRFe6oGrKahOYxpIpUr2M6K5D8RrS/GqnUw1z5brbVtGPmzkSUY2VE
+X6pLY+Qo2T5OrLkAT2dg8qVmohmIsG1IlIuRLKaoeNF9gTtIM9sKXQVomK46YRy
XR/BHeQqUme0mM1WEW+UBnoYg91A3Jy8JuoQ4rQGJzYerI/DOTXxzGS8kAbVglVY
MSTqSl85ZFYKTjUCJo4KN7MjWJdhIUxFGvo7v6XUPyEYQmIGazPAKQZi+UjIVLbM
gHjSHIv1iCtJi33N5pdRkuSzKEwHWYAX4oCxF6ZwHhZXNwKD2Ao7lFRFO5tq1dO9
uIXa1qEdv/UNHbE57AeS7RtHVYUQZ8zB7pbcJBH+qpeJISY3neQF7w9eMNQaoWt5
GvmA0BO8/AT/9waqPjRZL/uifc1UTdTK0PkcC94RY9M2m7mN/te1EYD1RSlYgfzG
Mss7MBsF/pRsOXGbUTfhStUsKKsFhemoBr45r1MiFaP2EudpVXHyhcnFI7EeG9Io
zlga/4hGkEkclINLpWCbolTJU9tP8CMd1lNlIPkTukzKvcgGLQObqatnyOmrQ1ZE
hBZC6VmhfdjKIrpKZxrwMl6O4RTIbox8Ex/Edp5agJk15+W0STi2+qGHpkAcNNE3
giR2y0y1i/6gTLD5/f2OYZ9nd8YR1H4Ui8Wws3trNDv1k1Xfw9hRP+z9rhqYB3z5
WpTkBVDhfMuMmZ1x3zx+hDj/rQ7b+VyOur3EJuRo6T3w1hqg8F5IBnG2pE5DB7rP
dISzjY1SRF6cg6IJTcF00rwBZaQjOU0IjsFUV91rnAznu6K6pAO9WzLTe4vBymk8
/ViPgQplsSDRAvxgJXa2xd9f4I1jVcPdkuuhJgLiyVFZRhmJ6iPk71cauGLQg2IJ
fnwrEW4zx3vbfj75c/fHUw5Mh+EBVPMyo6iZz/Iw8zGqMZgawQ7npsFjYzGeo+uE
JK/i1lR6DFJVgga6vFEV4g==
`pragma protect end_protected
