// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MbvFRg5i5/brl29RMYVS4CnRyVE+Zde8bAePJezJc7ar9PeRtSJgb0clv3IJgF1U
HjLoYjwqMDchFnkBDJECF1SYHDz/sHckcDP/o09W20grlwGIx9y+orVB4sKw9Umt
QnpiDKuHMfR0oGS8RDaGeZyymEuM2jPyuZWomhOFXDs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5312)
WmXYUF2LSK7vW99rYTPnrfcw9yDp5E61Aw/AScnhecFvUajkHTMaoA6q4+nrPElu
DaYmJtGpJPcZxmSVSQDnqeSgD33qthMpJpjq/8Jjm+1sp8A2xnFL9NWadeLZYxEY
ihYXRPKo7idFrjbqodKf7b9y4bChE/D9EUUIDQyxnp4xPypsfTgOJRgkxhBfusWM
4ouVub+xOcRMg074bgbFLw7TPSM8F6+JtzHjVmaDxomc/HXp2ygUera41RupL0yg
ZMheGEXR7zd0cvK2JBLn2DGfw/WRVuVfUQ5otsPl2HoMfUbHSVBCrKGfItqn2ZjS
KNW3CKxcIlEuE/BTge3mKN47qE6k7kDxGdkDHmwIoVTgRuFWOrddnN8iBZ2GwwIa
wRLZZ4xx/bIE0TI6vAlcCb27P85GQii9q0Y8v9hItwfkflT6BMdIS40vQBja+yP6
unT8XXn5HZIE2YdYWhrS9MJK7mqUHJ7j2FLfF9Nm1RHx5ZaKmpG9UvxAlZaFUBPM
cVX7i7FKK+ZClR3I5kMJuECqQ/+nC0jVjBmvUWXK0P1YLoj8BkvGVryN3MGm4fhl
5gTuel8BySb0VQPQZRzFGTFGGod83VJ0YuaBdmSAy6Ujp9t9w5hjv0l2glhN/enw
se0EQWLtdd4ELh7rQby04WfDgEaqkiXQF3EE8iAHzWXH70IXwOAaaauVWEyH4uan
+2FdNsBkjgPBZlBGNsTPpDR0jReYLPMhe2URNyIu00vngM3XHDgP8aHkEXS1QROK
4DgTjZyc3qOz0VuXRzW359q0ULPMwXO2JJpg89cMVs1ffLxR38yaruG7r5jMLz+v
pZpj1aNNSxb/I+ByVj28t+IiZxti3rlwHru1YDvlj1XO526hpaiww4MQpa3DGAKU
8J4AQFwP6+qoId+OflMpRA0QuNRpkET8Y8a+srDbg83Ij1a2aULy4PkPb1/1pzq8
1PQoon2ODXUJL0XVTk6YpDdS52vDP0CggLivZDaH9oP7eQMerv/eJGJ2fJbJ4Xgk
ES47knNlp+j/dUuJOuzIyaDvGV8raobVil+rFCUyOCLZWjdTxCY80MWTJmZCbNua
MVaXOK/fXsDz+/ZMor9gUtVsMnpNHDl5TIu3killvqiaNaEQ3+9FZLFYwla/l/4/
cnNwrY+sV+m7u2E5/dFlf89dYN5LhL5uZWvTCp2hyjKW1DMB07V60W57M07+nsG/
lnzC9EaVOEpMWF5HuwQKvgLPo5EA4R0zIpjVTYVB4e4FaWoaq5Y0EF53sDkRmOtr
Mosk2rCLNsrlQ+8XNxqAnk0cXl9g+wDfMAw1lwT68BFt25x8KXrR/M8pjW/QlP/u
a8hYV+iyIXtGkisCjOfwSXbUDGizpm1LJgdoY+HULTa++CiTXaAEWoFAzmgGjP42
G+iFQWy5BmvGrKKNkp4pafpwDDloo3Z8zKz2upy68DJPg1GLp/6dTMXGWyp0gYS2
WZdhaNO7aSVDRBkrnnPkbz0LsAygtA3qsC4AORoda1tNzEic3Y0krdgcHLLey9Vm
g31DEdmDknta78ABPW+Ullosn2H1SdrI4MPT1GeUuQn0PREMmx0q/QZoROrXyxmE
HGj1bC/VS1u9wKpYy/p/5fkS7y3l9d4zuVzqOGO2RXAfChPi0gAAKVRAlvNkanFq
Cp/P4P+tSJ6JL4SFk0GoP7HMQe/c6+KOK9h3Qfxz7Atwl9WQB6E8YPRE3UMqmTcl
KJLBSLpTc+CUOfDUqkGQJ094WTY8j2gwFNrAmFh28XZ1rne7+RaORPOr9bI/Bwt7
5arxA+5l//XEsoGvdJKUuqWbzsaRLFoxYIqEgOqXq5BFbJykRvB7RUv/sYCEK4h3
xXPuiY3yDIqZ7nBBAdszaHhyMaWqZN6VW/M7NITtTqNJ9+aOeNLa01RxM5BakNUY
FKWG8M3+SnfK3JyEHGpPiRo/rD6fai1AlzuKcqJITIGBMQ84tvzl7KoNmfJrcY+e
QWycYY7V2YriDV81r6FSd2eTkr3fP9T03/sHtQzrqAO0Tb4MoyciT/natDl9bXlq
NR4qJyt9AlmveIN/Y1JgMu/rwqcDgEN8mepgkUKCek+ikTeK7TCvkD4NHQEOPCLP
oFMsRO30ojQGHfxnZCHjakJfh5nF7E36dJZabEZFEi/0qEH29YDrWgB2o/oS5czG
zuNvLj2zg6cPsPMvkc7ugxmJ9YxSTarvTbIxm3zZQBoTGZP+u+cf4j9hfK4T0L9f
KQx/HKq6KdeKpa8Thln6fI9RiubCpq9jHOyiMdNPyPjodSe1s2AQLwndOcVe5jsf
4JgxnWLQhDsgiTiE6IttXYSF/N0QnRePI/us8biXHqLgwUkxQzi+uiCU8SzLQ8op
8FZdQvZKPKZdvrzsLCr7iv/e+MYrTTJEAtYESx7Wy9Lvgkvh7ls+w7BsIHeWX3kU
v/Ff0dDfGM/4oz+fni1UPgeOkIlhjALgTnIBTO6BjLAaDk6MSyu+nbq4PpPIWU8k
l7qmBrQ3PndZTXd/iPcas16AIrXWOrIf+Xr96QSVOu7AnmkLto6ADFTkhx1CwUaF
bgw22VWroINVns2pEKkeVSr4E46PTRxWCUdmLStIfbbHOm70JQs2V5KYXsznZtGm
V/Bye/oCOOahc5BNAnf5KAJGzH683egAYbOCaaMD58W9Sk6KqxGos8hWRmF2zA3b
7LnCDAvnR2VTOVWmP3ej/uMklYdHrWRFd9qPga88JuOV5rSJvIc0N72VMdjnqRkZ
ByuCeYzg3E8LOVcptZMg94HTZ/YDzP9pB22aDqsjeeA3JMBB/LXb3ULvLtlxe6s0
x/jBd4bZHc4BKE4t2rQDV+j1bNR1MSeBRonhXK8rntNzD1AT0X8bjdkeZ0haX0ks
Uid7CLFppU8KRTFZYPFWH5su4n51jlqR+2vfmniQrP9Tjeo+5z744jIcuVAHNKtW
EQ2HGba63Zy8g5NxSKCagciXIgPAqZ1RKbBOkeU4TAO8hY9PIV6YDFZhLksj0C6n
znb2uRmyHv7JAnAbewGsQKR9qMfgK3+pssVfBEIxjGaZ33XkiZ3pcwOI67O0fSy/
kInWtk5X+v6A+dvSxKNuONPtrYPdEb+sSZwPdeAijFNonQ2LIsIfQvivSTAVU4Oh
7+lNLrtKvsu8+dxZm3X1aAE8MJVmpmWiMX5h0SyZvBs1Kl2THKTAaqMrLhCGAAv3
NVA6kVukl3aV6gK1lyZVgYqLWTyrEmgwsXuy5VBMPb5E1COZSTROkZJJZ6bFlUac
p4eS4+bpNkxcoTaHiHuoYwM//UFpZR8L6PeyE1ltS+SRpqF550O2eWQYytrSArV9
siuFzy32fzl67eZzfzYgzQVeL/9I4R9rCLeZQvdZa4BZg4Uf4KkL46BmOi57Emx9
eh/8rhsFOMtsRO09Lt7HBJOcCZ2z93EK3emfR6xBwd7GjiYVp+TTYO2Z4ndv+psJ
Gk1Yh2ku7Mku5UeGdFcUbMOk/QDMsAcGl0ak/N0gmI19I91Zos0o2NDhbWZ3N6+u
7VhTKqBd8ap8QcDSHHT1lPf9Vzs4QaRYtyG9DOLBqDB0ACBRZZFDTVFnEAgyB6+g
uuPCG2qOaXYc8bcpcT4KqgAnsHI71gx0QPQc9VIaWxSju1Uh6G3i0McHcypj/a5z
uiOpFslwLUEDZhrqdSRM0WtJ6rA6FnoFcxSLaiU4prgKvCATAl48it83f4v1zX3C
Xts5Sxfe408B+g0W9/MWVIG8pj4d/raiPTQRb8sXC1xg+BoEddPwI1imtgflm15r
3o2Ci6c6BQHi1e87VyAn5/7L0A1Ob3t336qNi9Ul+WZ/P8QACUnjg//fZVXbPSxP
6m47zNheVhGI5qhwj+qAjt7dVlDe1W2KoTIIU0EWkW8C0hiK5szJSIT7nh6ysQ72
oox4lKyAFxbn7gH/Rcd2JIIij2CV5C2rqwEbTtqysTU8WbFCU0pQyK2o0ZpeUTMA
3WskwW3/+IPvuLGG+MKNZ2VaTKcwCrpzQ2pPHg9ODdJSd+fI5HzcYGaMP08Y100j
Z6BDx3jt5eMOwmMZBLBtH/ip5/0gO7rsjFfZ2Wq4furHxA4RT/iHeexDMxNnHxyK
ZuS50L5oq9wAuOq/qnWZuWNH9oZ9LAQbTNha1iqej1KqbkbvIeS/KMMFMGt8yqjK
GJTjPvlvC4t36KGBRXL9BnwVQbBkuJYWMBgfEgX/h4RaiLCpB3F+6bDtmaMsGhJh
+K5h6FGVanr92/w0MAi6+y6bePhwdkE8CGaTr0Gbs4bDFL6FIe98uQjRdypXbBXq
YzeMstFS2A5JJq5SBdMNuNRww8gacW8+epuE7EGO5pIty3H3KT/eQlCtBhdarQYQ
aKjWJcIXcLV71B/UMlcrtADndCmVdlFKBLsIkf3xEDxh8tFzw331tnpNOf8SCJn9
Wa7ilrTnm+YllSbAklmXsiETHNxZykD6acZBmR3aozfE6QjX1hwupQJ740THgVd2
fXdoJ6oaPOTfk20N6OA2N3xwV8faPnDR9+d3UpVoBVG3fWsIlwQZAvViwIJN9Edg
9jiTAEMQlkesJTThjsNzy1rQhcgAzN0j+cO2nhD9t4LRYYb42GdXgMsJ0tFrZuoL
8NSYexTYoJR0N7Z/7ge49xZU2/raz0QwY1puMSW/JjnJkJjOsFJAgTsQAqeQeVwR
ShmL6xH/U3MhPuSyOGdwDvwBJo2d7pkbCgR8tP1TIFd4ysp+7WG10Rw18dOPTPmS
0V3mkw4JXyOBHP1Z1sI8jFPSsCkQkLpvvM8rqQz9QFrns2RX3DT8PZV44jKVvbN4
3E35RkG3f+e83QLiLWVHaxKbJSSE2X6Nt/n+bJprwVgba0XxZYhngvNjD6btT2db
iw/1aXJWeOgSAwc9I7d+r4xxX3ecKGFfdkfAa+hGe1Nev+A9s6RPcbpoDU+wgxs6
5ZQojT5UWjVgW8BtIQH7ejxzx34wf54zoThGxVBwg5/nR4730Zf1hXjwlSoWfZ7G
xEOy/ju08YJdb1zl0ZBpDD0QUnRhccRq0K+pjo2Q5vv3rMo1LQzz21C077tl4koc
wGZH6H/Ygr7Utjt/tA4d8F1k85f+vOxGO7CbbuDpn3/XFL7q4RqZHIcW6nQMKLLR
ifBh2bgPNmv4Tct5o4xNGtQlfgqSE6cM8doc1cewjjNaHFSdMFqCMdhC3cCBzQ2R
Dbun+4BMEDlUtxp3zVP8bzXytlGA9ZePqmthupuqpx1zV/DorFrEZQfi2PKu2RED
x9z+y65TXi5F7wFTTtkdNr7WKrgLU7AvSbjYaQQ8VuR7Wltkp+CkCe/em6MszWt1
OT8M8VF7DvyjLAoYnDPYYxQL7lAtL9MKI7p7dV8d0jQVQ6tqfsQdscU3scazxYVN
gwNC37E5IZliINjF3vlBQOCOxB68I62YMkF2+v1EBmSdFZ9JbnLtwDkX6u90yOgm
4/CA++S8Vumrns3zwft5VjznVS/9CovU2NUPMiadJ32lyRDf9Rk8tARnWutXBA+1
KAiEn7yov11AaQQ/s9dYMK5ThPYxY5NQs4oN6vM1gR2xArMP6zJnGSm8YcKqKf1z
4ZDL5Ibe2cgb3J7nsTbmjnWefQKELLVo0j3sOkIDe2gsSLdGESW30RtEGxoD+Q7B
SNHI5e2G5puD6f0l198iCIEty87c+n7I/lts/GgfX+9jOS/tQriYofLTtWn9Wgri
b1UPcKxBonGdbXumOLpn6tVwarllvZebHV5gNieev60j/cPtvB9Grxx/0OrJFSLH
WnrMBcuRZ3vU5KRa8kKNb7qDmYFKpMonmC2CTAyDM5ZS8X1Xv8PkGKnQewjF7knT
77UxyF1XXfQZ5oy8dn4IdkY0qbca0AS+yoblXRR/FCGxwVM7b2tUCsLDTr50tPcP
NqWmOYLn+JFizv/MDwVfgfDQHpIEchzAGxqkM8CAc9KA/Eak21JyonA2rFoS7XDy
C/53hgODmWynMwLJ3ky2U910JdI9C9QGrQDp78S+N+WwBDlRl9ChmdmNralGUM8j
MTmqazhFblqoe42GFl7j/y81QwRtaoqKXDO2dcwBIBS+pjksq9R49pU/+Tv/JnAa
qk3LdHx5Oy61GQYHmX51BTmSzveVrbAGZomtRiy3Kypxis61bmWHoKjHVluUHLtt
1KCAhoKiMaKQ8ZLegDgnKo/XWbK6noLnt1OxveXEf2VOehUQbwEA8m/P7kPtJr/3
KK8T/E3M8iBAW355kYe9hb8UXZ3eXZbrMGnrb1hfNUk1xhoFvHqcmTu2SOLUQkp1
8NPdPyUSe/AkhjY6H2wTJjQn+RvOpoO5a13wyvWdpxJSxF3UUZAbsP6ZGN37mZ6G
GvDc56e6k627BZv97x07JKugJsLLGIThadlUinnwmNGKhbeqkTPgtmaQ1bYU4ryu
K2FWGVyxM+igba9rXn6ScqVh6i+0LhI/cS5fSUQ80tpeZcAst9a4diH78bvr0osY
CZcWKTYDnaj13Vg3LnDwMZwScMffHsWuUub//HYXrE1A5iBnxDIM2u83Tkdn5lFg
zQJ8Hrg4ng9z5GENddAfTosCORyl46FqZJ5xeMSvIvDC78hQcfKxgaGV2CsVUzf7
3ZRz2MWBAQ+WG7O+w3aFTqEfSGjz5GkRzCRRR5uDSbypzCVRIdict6U6wFvwXkyo
fkKAIHX91fkenAhN06XcXkujs13iAxcaJdrIg6Lk+pnDCc4YsCZs/lIbTf5yQTrE
U5SWv30rr15QjBrtzeRc2MWJFXA9H6fkABgIbPiw4jcBagU0ROqe/AC/wVX4+Ggr
HuIU2CJO9q0qNQCNwA5+vAcO65y6FL7s/3gk2Cb4MYM2HJHeAH7fWFqWjbkag+pz
uepFASqAkwm7tQ7c652OY2ozkT7N2gaob3nSutFUVsBkP+/pnNyvOatZfnXBc+Jy
BAXq/2wz8GCFWZDLaZYU/y9d+liIUc9xlkahauhMA2vIeTGP8BXas9wRybgQ4hw8
A2eJsDcHxnYOUHnA8WNMHk6CIHtNbCuRw1NpraAJa4lcLBEQ4PWqKmeQyejz6mnd
NkTiEU8qLxbqDw2v9sb+WftRAxGL3+YLXH+QA5y/xf8=
`pragma protect end_protected
