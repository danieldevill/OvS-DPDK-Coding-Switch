// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bfQIFQbYoZjgFRqi8CTsbryKS0a6SXYeF6keVKlqul5KX6OVztkMzYRVFCBCu2K1
s4eM9JOAX1HxjH8rQVbeRd65MB3xtq4cslj8U7r+c9x6v5GylIOLPf/5X25Y+JtG
TgOdnvMvdbNHRx8eY+j1iAM6vX2Fu4Bym+u7id+lYzw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12176)
MXtkdi7RS7+8vJrzMrf4G5seCTAYKwHb0wOt3ER3IorLLIas8eY4VdCa3w1ECxlC
8MIFwSTqqEvbuhtSusUYn6dONXvoleYLQLlhrb0Y4pCsF9q53x6MJCrKrDHX8R7D
fsfiDSW4EWVXybnxYSBcCW+bFb5zbCLFmaQYy89uzGBh1/o8crbrX9FR9w9vRn9e
L1B2ndoL+QrMftv7jahqo3I8TrLn41YJkkeKTafJ9SrVockgi8ooUA/1pCfwDgFw
tW6yLPg+SVMSLZdLpmdu9X726p1GMCB/soO7/dlkJXl2igwuk7ZG2/2SZo1AwcOO
l6mx04381JTU7WBjaQBCbI8sYefppXjip8FPc2CFWbchk8cWwgRLWUHqVNSngqBb
EetWWbtEtxgkwUn/Xxn0cJvuBrLPE+X6pnbBmBOSUwo9jp76G04jiQeuyAP8pnNz
QR0MpARP7Rpib28iwU6r3NmUkXw48n5LUugflYW34sYK3Ke1kUsKGbr8xqQT6R06
ypvGvcwFliHLbF/Mixy8zv45p3gQyBvx6m8hmdUTugM6NJbP70IwPZ+8A7+QecRO
skbfobLyXPrYr8UjSkB3dMy9uMHfb8xQiMq+ACpx4cm6howcuggZSC3+YRerAcIP
t8IY50oLCvlyZM6E+N9DInMMYLpR7h1gxXSfXTz2hsBu8HXQ9Q90vqqRU20YtLXR
Q1rswmNzDysxkT8iCd36b27f/y1NUEONIoqpfhJOvE4RLatubxY9v/QbNryY2ieD
b3gCEHFdc4pk6TeTWMhGwUwv3/MWbYcaCiTCG76BUR9KGwoisoHA8oFJH1Wu1DYh
rUZYo28oAOdvQFYIn4Nm8vkU7EuOggC75JN5OJifwNBBqSZp3pjnjinc6hvftoG5
x4QHq7DOJ7pS+YZi+3xKhJfys3a2QFf+exEVVkz0Gq5KSgPgOUSLsrn6UTppu/fo
/p/YJr4Q9FUw6CIdUCIayVSr6LaEzuZJxpNZiIQdDB3eOWemJJrrVmoZoyuypXeI
BgMVuQSCXeSHncum06WyuaVZSLyuhWnY6JV3669UlcYkmHE6r3V+zg2F9lJ73JPx
MMIiaEMnSKeoOshBHam1PzBSSo3qKWUhsf4zsAvXUmjqOzncGDqNNvwtPFHxEFDE
vWHOtNY1dwGuACSWpo9Ki27z4mqMW3n+DXrWnluGVKQzqmSkXITCuDKIWXS+4XDl
bSqJ5TRphUC7ibKOQOo4uuTVDyoX3ghsTXv8j8S8ui9uqvZ0iE42xtWf+eyVlkLA
Uni/vj36d71N0jr6x5Fyd/KnDaFFABvLsm+nY4ij25ucC0cs2VX8h2qEBFOaxpHn
P4qeI3I/xv9icMGc3gom4q1jj+UgMSBXMXY67TpG/QbrYs72FmTXqNHaw6qY9V6S
UUj3JhYNBKnczT+wvnsiYaLxjeTpthDdmMzbZTKV20p8W8IqGGhNVZHkVHr7gZrt
NdWQ+EEwOQ5PsDAxOTJjisoFX5sIkm+k+H/xbFiEzSwmqzDKnZ1ZnfVHH9mGlBaX
fWdo4KmBGJJlIlPokJsg89aZPbp5ty+dPth7JxSyI8Hl5X2G3LvINO1Q3eQX2A+3
lR+pXlCKvXzaIYe6XMLP4lIu4SwNGv+rLU3u8Vnign1wh4QGVyDZB84AynNKR7Iq
RjjHZ3AndONVmNR37U0Cz2njTDBR0YuDYUfyS9YgLVKaegF0A5SxDldhyf0UW4Oy
ZMH/iumnul40+uSjPDvgD1BM9J/gxVUGAt/WPSbFI29zbFutbzE9+iDralWkn1x6
FEwEhSCFWXXjAkDs0TS5oHxVOCElwUzTq83c7LgdfKzMbkiuYHL3XtUd/A0836l6
ROrEVvgSUTxZway0XyWUBvSd1hjTc1reEZ3xkwL3Gb0m03vYgey1paa8ZRKHchXf
ti7DVkF/sfY7vpYrzcQdGTyLaY9BsPXbXx6Rj5DdHL5ej8/4tsXG/e4tddViGYC7
5IXSwfyYcops3gPI2pTpsr/Z+jyxCvzBx6YCPjroP11qJlgIESC9yFo0Rz8d8+Ft
kPAuhPCcZeEBNi012uzWOrFvUvjjQR1HC2kh5QZrU83Ra81y268XRM69llp4Jg1r
jFUyZJ1XSfelnTFL2aW77NUijX4idmn0N+6qxszqCEsGEJ+rXuugNbQU1q6Vr1Uj
sXRFeZB11iPOzpDIBbdt4EJf3OHUNmF4gG2eJXBsQmpC1Cy1UPnOCGW+vyIP4zrm
2L3rQNrI5vZYFO7CdJIWfnN+Yes3YP7Zv+H8s4D9Vw7fmQA3T2KqBA8bnnEpjjhJ
DUDfGOcKXdyeerm09/9V9ZO4jqcWr3PRVdYN7aLDSOseWd9AWKdHXDB6n0y65gGz
ZGU83MWwD/0adn0rZC4NNCP79IiyRee70CjJqaka1o9VJN8ek7rqXvp3AI5FR8UD
B5mPr/0Yh3e/apWWWNNKCErMC5JSAwqPVOX9xy5USHvars6elnja/jbBngfWM+LH
IOhKzcx/JacndpyKhP41SLpnxB3NvSi69Pf6/H9Gl86SRKp/TLr2c2WdHxNpQwAU
wvARVjse8KQB6CKDE8B3/HOo3qnt/a0O9mdN6j7A0JMKxAIrpbhFvEII/6xxWiKa
NqGp4/QWW0OjBVTpawpnpsbiDBzqLvnvXR+PQOMqbetEDw8ZEwsBSxuRPddsiLbu
sogyUkHp8jXb3UsdMdYoCgY9wItA000Xvo1va/BnFpLICxnwj1TjEeahNAMe2HNo
6WcSJd1nwEYJQ4eAtEddDRupWLrdlScX9Cp3e9O9ryVy4srBKBMYt+27Ry86Hc4S
7qNEXpmhsNNSkRx1L+9IIiLfBBirp1x5QP/mBQiCaim7YZr0g95f5RH80afC9w5i
jxpiDj4ZA8dfFf59v6vnnenNEWzwMC6G4ahGwRR0T4+McrF/xy6RDiqgHS6x252A
/O5UyGB3L8RrewWAHAGNc56n2Za0VKXw1Zb5g9avAUYNsV1cSEgidKtHiKtjmXg5
HUnE0Mpqkgtzh1KwHLY0yo+oIkIcS/CLDZUYFsAqgP+T0Wv10nOyJkoKCOrLC9SZ
o2kKq5RGCcBrmhWcd6nXgNGJr1DwtUWUqT2wMOdOZaFsijLmb/jr9NjW2XzV81YG
n3KRUtTIa4GSvGByZ3VjP0oIa2Eg9tCVtSH47tMLK0nBKYZBPb0s8alEYyXs6wTW
umP/OIgfNYgjqMs1zzpxRf9WY4AyRJxjUUV6jP4F7apcNghMxBp8vu428gow0HEE
iskGYApXk2P6Rl+mxsgHqurq8zC2242nhPHCXDWnFRHHi/wtV789OpiGzKiUKNp0
UuBY1s00/wHdKvgYh77aFl5HiKxrg5cvuvHw66MfhtBluAkJMDyGRfMVdkdZMnxj
4voujfwZWUmz3wOelRtX/pqHkOQMbUCzFBTaWU6VtDoYhdmFd+Qc3M4nMGuafRdq
nBGEGQ8kpnmgGs4NEVdP8Uo7yWYJPyzcsxRzJOLv0gjlp2O0VIxWJvwkjuQBtv9X
Adb+M7zHjOy8nY3D3s7eU5RzhFin6dIcE8ZTx7XjDICo/dluhBDAXBEhlRZRuSAG
xp6xWS4BU+MkYkLEf9lP+6dJhkj7xy5a5HGPKtZqJj/zMU8u5EPyJp1T3eg3KLpB
H8EUS9dPpXtfMeSOJ/Zdjph/Y5yisuX58Dc5PTLklX00kqEgJVJ6Ufn+T+QwmHJd
bTKyX9SvS8wxM23csK/+Y70AczrVQc9y+hqgjWPIoWbB0qrCB59Dfa8nEde9pCBV
v99tzseimXrvoWvCmLAV4AFd+VEzXBoEnUiOciXGUKhWpjjQWdYiiOnmcHy6wtTf
1Beggb4abTaRO3ZHO0NyfYU4GHr9vWL3U7Lwite/PxhVsF/p9dH0DuqecxfMrAga
DoNnrGiaOCQASpbtt8uiHiS97fnR9VBI4iJO0uIH9GL7lNpKYWpxMl5Fuub8RfHx
BU/JhNfACwmoZQWYmbM0LdRaE70pGgVaozPz3D6vJ0qcEpv7Ky9XLTlzTEFTZ2YT
pNLehNHqyVOO9unT6FUpFvrElK7kHQmKqqJj8SkqEyJ8DOCeeIY8o8+GN/4pxVu+
AX/h/XY+7J+NLcz2VNSLXK3Va50jgp4ZAgabqbSAD6Vsv2G4oWJtgSjGPFslIJSC
4hNl5zbEp7Xa/IxsaHn7L6gd8TUnYlzuMblDTWMIZSb8kg4WIW/9/uvnDWc2PphN
Rq/UL+u1p6qjsaGnI4GRyvF6gVEdOezyM7aCxcomF1AE5thprmkRddstLicpuJh0
E8vBOQ9D5SjOVh55cV+sl6w8wJfOdVBsWNoXGkW1O51hFvf5B3dvPSem4/3+cnDP
SdFvt5tMnOQ69WeKrdlrBTZzdPVp/xUjWNysZ7PEyj5GCDIy81LQv0hDEcgO52yR
d7/p9PHaFNwOYwBsEmR9+xJw5kMhoCDvDW3uiE7tNmMJ+AWKg0at2ooj5q7n3nmt
ytXNLMBTsowPDHFXMXkYRsD1kmsjgPfm2jBdAvYHlBrtZ7hpvXCZqBqHU/j1O25F
qfcy4KHBI/3UrXapdoR7VJPby2j3CTDf/cjATgzb3fkwMOjW/nq0QNIB3HpQkPrc
9uyzfp5wEQpeVqz1P472IUD78N31t3XMzaL1OEgDR4arqoaAqvVYlcOCUGM06U25
cn8BD92uPEKDmajdtQF70wwx/03FBKrjdc51N+l9HDmVWgV9oAWvr1GLRT38Vsrc
QGMbw60Xq4sKNUMj1ZJ/N9mp3CVRxEms4M0i0gSTcCfxn7lcHeDvJAgx0k6c273J
Hg/FpASDjB88R8dkeCsjwPLT5CtTNS6P9gz+pqkafK5cw0Aoo43tJlBr+QgyuKJt
w9eSUEL5lUoHYbKSN+OhqV9xZ3ESrhqTOIWLvP/4au6sf59xo35Fi4lfaNt3Ywi/
AjDiJbjudQLlAtjv3NGMg1eNIi/UcB/z+2H+VLyeoQEw5/TbKUN7WWdTzxpN1j8s
5Dq7ilNduBD3M0OOaBixiums7IF8bXFPiUU3FiEwvwB4FvcJs5W1RhlxhimfrDlx
0DXCLmOW1+xXG9CIZZ4zil0wv5qb0ss25QR5KAwCOaGmkVub5hmDXRbGujdrphzo
PVm5PMEkLOnhVb6Rhmps3c/+MVs0IcGy7wtqK4VdA3JNyVO0aWQUr65dCwZ7Oti3
nmYCnsOowomOHi9Gc80rNHTysLwXtndPnE5Y1YWhgB/tkgJidgrnJO3EE6SxxwaQ
rLKpkxitzWv0W0qc+U+yv9enOsJjWQ4GWmhtFIBdwxE4pb9qdsA6LPq4xQxBEBNL
TkrLnA4IN9jmJVkY126jBrgOYQsJ2QPVrZncpwD19+N1x1zV1x17xy5upd6SYDpJ
/0SRxp5Dz1zZsUcIqoM+YL3PxlmmRLjDwNyRBgNsufAdXZKLxp6PUjqNWLNdGM2O
HtL7GVk446qUOwCbVH7pKImFvabScepy8njRp37e79zITeAqjTY75jsLlvFK2sJD
0a23VYabB+ykDrYIXCTbduQTS+DixS6q/1eHucM2Os0E6dA4UkVWXzVqkj+6wUlh
mfDvVTswry371zXi84WGN3NygWTEAApzs52wpT4P2mq3Qdxp/F5z8b+Ig1ylmFl0
mGxoIf4Wcbq7hyu4rQzjMl4om8Gt3mZcnpSuYqXF/4YTxKkmFVZVpo4cEUfdjoMI
jpzF/Xrx43eFclXfHXrt0Y3ZbB34MgwTTDKCeFXr5CPQCegmUsbgvnzjRDp+wzjQ
pNIqVE9lo1yoWnfPgZ0sy/hQVnX7slwGwefssToJs9yXsEQAdLjdmzfyrIrxoN0o
HIJOAWMLXhzDtv0h6M2X0LJgAYes94+e7F9dvVDrPhmk8C1UOorGnvxwQCBOt5lm
NPw7SN64TkkYfpavi4iZaG9bf0EeOWY91l0mlv5FN8tc6f31Iw7XdDxTReulU+Hc
WdDv8+LWYsT2jtrUxjibZlcmZITZ7HL6ji9Wg/1IG1ZAiFXgT/QLj2lVwiSP8c5l
7qGMuZ03fKwWiniMG8foujd2Ycz91L3eLznvGYWgQfycODVGr1Umqm9Od13SregG
fLEHjWRbaLCqzjunmRcEJ2J7PTD/iP6W+Yo7aGmlPI6g3t+JUMEc7gziZUNQbZG3
IzpqMsjN8qZja4GQyqOKCwml9ez0lMZZwh6Qe4YnrnWFC6GwOCJjMgJ31/tvQcwD
V82gDT/KMj+4WIgjnTWMmVUbPSa1/ln6rHdQ0PDzcLgnShi75GXpN4DIjar13t30
y24YqDBzPiIiLHhRoVvjrLZUcfrP6+RV13stYsRGVQZWYyetLreNL8AYOliVgwUq
d9P++QZ9NbN4/yUJnkzgaWwmHO8UagtqqBKx7NkQaLuYYH17mQOFdc7eztyXgNwy
2aHp3z/Pocuw/moYxUNtLCg9X7dGRF81kg5iJdPqI42/dSB9CFp4fi+1au+qGteT
q5X2ib9PklzwGueGoHRIRsjMRnE4x584JGeUUtoN9wCL4kBUIrvxtk9FAdqAhZ3g
klXbD0vH5OuhirqwH9GWtdEBU7gXkvWHifISj8vEUyiFneTMHLLWwYh22QHJZHwY
Gsgr2s2NpNQuNdEuxJ9aKSTBFDF8h7xahE/I/pmfgSPFup1wH7LvHRkPw1PF2EJm
norojDSySTgXZ7MwAfjEQJ+zjEcQgAcKw7AVQLR0pYeGt5pH0EmCZnfJ+MushVit
mGPbbYUVoQFrzm0MTiwD4oy68tL6fAeByVTTaEwgVd5njTprQKK8vyHGTmsc4knf
QF9OhJDoV4zbEv53GXnXlD9k0sDF/QnlHC+MxxEwfczUURRh0sDEmBhBNIfVeq7A
v1w32Nsnl3TY/fhNM8UcbKijkK1Ly3YwZeTmWViYNvC7QmHxDlUrXlhlo0fNpFEM
Nu/x0SCkZHzkpJt4HPzPRAU9Cz6maHCysvf65hq3xEy9hvsph5BYoWMmLoSRqdeh
T48B+IAwm/G5qrJNdVBqO0W1s3+e2ybjpowJzbXqgMAjg+P82s44tn5eZeCnSu5d
MxysPgFmMDVkluQzzfkX+WHu1hgmnu4UPBf0nbnst/3x+R0jY9RzCdbGxfZTJgVh
Q6j3FfUMRR31UEEjsAFyF0D/N0VaafULiyb2Y0eB4y9zH50SlB5Dy9t2XU81sUT5
FMiYCay0nP1Yq+3LAWpJnVy6AEF8oZUmU0YMCkscvmWYnDUGcIfSJuFkDz6wHziw
aLiB6ecrEjpYdrbtBUWjnG3M6kYnrNYhYL1iRHiYIIJDqvQp2xs5La0cyQt7fjSk
yu28f1rKlsd7915nPvTGtT1cKN6BecxM9l2mP+HGlhpUXxJojdUow4gp8b1CEOs3
HZD1ky5on/ItYCDl10KGhHjbV7h9ztlo+XjHMdAVA/JQxN48g0kDLslv0+BSVT2J
bTFR6qFc1etOwbJQroPiSyHIv2BOqPjtCtZC7eCd6mjFuBjUZQs8R8+Cfpn+ag2i
CJnEZrmURRKlOMFIdy4b6h+uoP7yS6bqWBNRcihqqtTml97nfqXa7QJ9wxOlrwU1
zRXCnYsO/8Un+s29boujj2R7pEBaXbQ4kjGCd2HoR4CLxCqahXkj7B5RuteFe6S7
8sVontgJsFJhiW0P18YAFFZmipGQBYjtzDKHewbFDPaXhp8Z94s2ub/zPnq5KXLr
f+7xqQuHv61Kl5tu+71rhUCc312TW/NCyFRFnco8jsyj8ruZaafaUOZxcMSNw66B
CFDtOCKeam1cRunRCJYIHnK9HC8OCcwr9mslks0ZFAfNh45in+LVWK6g61HBWJfd
ZiVx/2xrwTaOA5tO6fn4fPs/bIAcmIWbVFqIqERKGyjtV0rCTjTrcabU0bJgOwrI
wzpY2sIg8mcMHxO2nvUzAFTt3LyfvWrnDOnHt3Ldw0kEzhfGSOXC++yWs2rLhohk
ZfaYqqYf11sre9KTQ9QiZh51Wtfnnwgn782D5OVHaamLJCF8AOTH0/mBRcG+jtU8
QMTNL/4XsoGvsaG34XCTn1S+YgM4wQjZOcoG+NuSzMK6oZynw2VPw6i+cVjhHHR8
YBkLUnjbZxwhyD0e2pmockdGpEtg3FWPF0HtSAamgeo47JVqyHxUIye7HbQT2Dt4
/kOsai0O+hBXY1SzjLjuSDdy3u9wXB5RKDHgAS5BIQXmJSbR4EAHiol4HS+QdBBZ
kcxXrPkvQKAP6ooHD75/s0OUMJcvOAk2AyNOv28UhkoAVdYl9c6fT0UVdBrs1cEd
01eZQDZT3345/A66hMi/NI5fY4tu+dNmdPXfeSpB9fkmyoxJ3rxncPdJ6CKdthJF
aZZMKPI5/vNOGLMAG+q04NggeCrz8P1HpjvZKRwdmRY7AXGb6HDcppWJJnJPQxeh
UIMm6yOXbZSLDEkE7KmSbfufMTNRusECdNeywd4ZHcXtGxsLPcvgfsR/I5lKFxUL
U3TXfjYNwdocTD/slOsXetCBkm5m+0MjLq37d5UjM57ZIgLDUBuxUZ73LbiIAPTi
qJejPLbHR7ehJsIa/cw3sIy3v7P9jUMNF2vW5uNB5JEJ68K/Mt2hwrh5y/KAdBT8
Ncd+UGQUnSVgoZcvv1Gv2+q3nuvj7nuJZPnoQ+Xr2Oy0cqqw6oNK07c106hSc2HK
3HbpQ+GWJvKZKrZr8/ws76AUIgZi/QQuMjB3seWhenMA7CW1tSgzmmPKjLScBDg+
yPN+S6RCITmXw72208zD/ly8N/1sSYRqGGP7govjop1B9825DOUa7PDfQNOGk+ob
RvYBP4um/6v2mVGZGs6XxhMqntr8f9m9gs+I/QJpSiTXB/N0D9nyIjZrzLRn0tnt
BSqLpbydDJ3LI58o2LNPxzwMZCiLUMFebDesNhUKX+/UrWwswSis5fX2AEwK1xUq
ScFVnTHWrRqYqm1ark2JABnwsBSdgyY6bHVnCdU4lGkh6OsCbX/PNTXu+KCds+Uq
lPfTO+BUmit9A/6ijOSF83TZFe6L8h84otmQmIZ58fI//J32qtke6IOsQ5YAszIk
7qlW/ptvIAFgvnn1+S/2VstfaWlIlBRbHlWqfqNVXBKa8XDnZuCAlGpOwF27H0Iq
iRTWMopYkfGjpMUNpTWKGsPkbSUj9ZMoSUza04ubfBYs3fwahUg7T9Sd6xSdZxT5
tnzbfKMSDim9G9IyVG3DrGEXJcBSbwNGZb1ooWVaBk0eVXmE7fjpykNx/8XowaDh
U5C4cev2bTVTg0DMkSNLdQwyWPt6lxlT6IMlvfaS3YrF4/A/xBopGnCyG+xxYko2
NKsV3NYx5N3OhDTtdTKNwmX55V68R5bFRQYDRWlWU7jwZFiAYRMGhu8a4l4WeBsp
W7zNShfkztJv3+9TeykJvdMIll5tALjq6bqTlu8UlBwJdm1e+2rNaUXYC+J51p/j
p3yN7sj8zPV2XmO3aznB8QSrt+OE4IQsXn6ltkDM1kjm2/J9bDqDbe8xUbSuJsgI
Qk007OTklkww8t1eaUQC5Kc3RWW6UOKqV3YxolC6dTlO1iGpoO3VzOnbTN/b4err
uKZNPO583D6tu8UfNKsI3k8Z65/2SyoaOvAly+uNAIkPoJlyr8aRcfZ9hKVUSwNI
fx6id2+ASr09lWeddrIafgwEg3Yl1iSvCmgR39465Wld4hoHguDuFzL0kWp1mikY
Kk7hUP/QLG8/q69LDKE4CLWEno9ubPh2/eRJFb2YlJ1xp3DPSvk1kxqBjtagQ8kR
BVn+gnGeJjttjNXgbJ+clS87fSq70n+otFcWeZi6TKVW2PZ4eI8c2q2CTN2f2Tso
atbT0HZ9vt3rNcgMp9bTHfzD6enecKOd6hctjaaiazHWK42SczNaaHacRQrNFp/b
UoMhij0KmH35nOJiqaaD7pknfHHcSjZHm/nBKDM+1NQrSWCZu/jrtPh5vfkr1Bwq
6kkLkemJYTXIDfzsNr1omJ3kVEULx6mWJPoV2d/GfkgdzA3A7dF8huF47FClVBN0
GN23v7fRFo4n4q2hptWGkqelOum9AVyzK7R7rfZly+caGW0AXoiNFRUkveDvYJgr
/UFx91c35fMLNdgLCati+idg77qgw8opZxbj3Uie0ku+MNeKwLe8JyKK0T9lJpkA
WhttmXxeTfDLpgIqnUS0/bzhzZc6yrCMMVyLqlWjjUdLJivDAAuJSlxrqkj+989s
RNFdWg/VYz5yBOmDx6zaXOO0AitNHZOinW0gzeFeubMcY+LaQFZXtdc+x1h91Qmj
lR+jVvee5zhoHcrnI2luaVM2uZUb08VQE4pj73tu6bVSs6uo7sxkaDujcqw+TZ39
WZPyuBFVSDEaNqz/+xrmoryRmxr8PSUbJzN0pYSWqaYHkJCm+tW9pihzuqooNNRh
yL/LZ9VB4NPqz+3T9bP5HyaDi+F98LzRgs3TrUXj+WZyGgYKe4/oQTVhPLT0pqqW
RCJa2NAI9hiVSkVBC4nl20NXFefDLmrOZQjaN/q/obt59fXqPqsy0tavEO9xwl4p
DQ3cO4N+vdF0KwzVtqRfcTcM3vWPnrBxlouxuxkFLLjCxw0narEBJDdQR/PCx7fm
56POqAB5jCe0VTRLJphZmU2pPpRiooGqvan27OyImQjRBa4ghVRy6gN757aB65yd
kKkid3g/0NrAjZTjjdgeeJzWnInx8nqzyPR+Ha26B3svEn+CUMFMDcDIqdFs7nt0
zQWZ+gMAVlLb3fnKp2TOV8MIrYdMbDaee5XTyi+J7x7/RfM7tH8P/XD11raOy12O
bOgvO09L378scNDd2pMk2HUXMAi8C6LEl1nkaVxGD3FplLKNDYc5Ze2fbiRw1NLh
BdyQIVsKTyxfW9mkaedF8Z8bcgOs/ac6L2NvHO5bz8oEr53gut3bVIibYyotWuda
AOuHC3yiQreovmF4djI0Qaex82ZaPXfB7hWbt1Zgr4kjWRj7ZT6bJCIFg+ltDimd
n9QsMsjKGWGQuF2RahG9W7KFyW9sihPYYMDtlWyqkxYzgNddAVArcwhRrcQnmK9G
dVAs522ns9A6nfyl69dS4dMH0oJ5+cKawDf2zvwpcYWxsdKA9pHOvtnIug+IgSD8
646yLu918/cCwnIjvZBB12CnnFWGHjTJFUlZVKOZIYllgoebp2fbIskIN7V8pHn4
3dlUow8rOT6wJ594iKEs2DX85I6RDiraJRTbb2EN+WljeRZhHLy7IxvYFPXE7lE1
1Qlow6Fe3V5KPzkPABU0aM93qRfzeuObR+gKesdAnYlTN97pv6YuuENzS8UxEX+v
HQRgbJ0asbqH3hMho+iJ/Iy/RaAqGgjhH2q5F+KkycKfVvpx9raHfXBXK4bibV9H
HDOUEV1KvOlQSQNcRwfdJbwGyYIckX+SmF6RnyMjjY6nXzg2Lpm0IHfOgvbONieq
yR6zrwXvdgJWN4Qfvu2kKfaRbv1mhPcuzaT9bB1QFKB2T6M9gM2RziqdpXP7fUzG
nRpb8wZtNu0yTOa3DCpAx7YK8oZApgJ8WF5ipBpdk0Day6ZpOwkOSyBG2vpj6MJl
YMrtvoTJFx86O/hrcUbnv75tgIs06uc3ijovFwy53u5jQICPzfAbVD+XcCyOLC9/
V8n0geUCMWAjmpa984n2MMhMc7mns0A0Jp4erBHjQFMKViHkVgSj90Ab/LC2qwcg
t2xV1vkVE9sjOC+s8nu4jX1gb9YyCmMWesK/OqJBvivEZJN5hu6Vz4qPG2BgNoIg
AbqlHUwppQ3TSAe2cLWMvEz4d0wuB4agV4g+L2rUyrUpgibPBSApJ3UJtu9AAPCs
AUhlzFjn4cd9C+GY0ZWi/94t0zQqkmaYrkRb2rWRd/wfhyl1qlRTZkHpcO4K/S71
UeTv3ANlWqeuWaoZ6fiIAs8FbQ3X1pFeVl3f2zzjgty8JkHGIZfzFS3seV5sIme/
iNhiXSesfr0EWgXVaKHq/O+xsG2SZStl0kGCIYjoCdF2ZkC5lqwrH/faBSnYZ6Ke
rSb/mx1dZnkESkDK1LpK4GQ3FXWMuS1G+tdQJexBH+g+5pHRKSkFIWBtu5kYMwTJ
7yHUYliT1VSKLLKRQiImspOs5TQOE7GZnV0yyus/J25sO9GqaIQ5S/rmL7AzDLzH
7r6t12WYRSv1ac1Bufge8Rp+eWU6II2zn8lOMzimVvYj/OpW6gkfR4AUD2U4Nw1B
RqT7fGauTlPqHXSTW46HN32SVgiw2YTKkyonnadCd7s9gAl6/2O6SBPxFBu5l0QP
4FtxMg7w1tf1cH3+hgqNVOAMR1LPW3MwwR58YPZTSvmoKFC3u4wkBYvfacPjx5wM
O+fKHRR247ZPbzc1JRhbP1aSi1V5vLP3AO5M9k/cpFlXlDjDv8hsXPj/rpY6lccx
mDI6FcZk0xRRVzGHnpvfalN5fPyj9BDiVAoeYVIKQcxCXHxoh8p48Gm0AspCRqxM
/P8chP6OQ6UgrGRxsyDQu+6lLLADBAX3tQvyHWq4goDQLK2nF9l/YbInuSHKVc5Z
UP42mL1O9o1fYas47w+IE1d/as0mxH0YBcMcpT+dp96HcGUIv6VmyRVsU43wgIc/
FEU6T+4Ac1ROw0rtMrPGQspKibqJoSy9faZByWKg7rBle865kbxqDkj2wEI53yMH
LZO1DO8cf5cnoLZfZ/uZ6j8QgdYYvTxDySRh9Mg9sjDCtBy+VgmLKFXpdrwnRejz
B1iQTFFABVBkvP45/eaotRhTkSWvG7nAUOJSpnXMCHD8JQ4N2Y09kizKobw11mPy
x9+8FsfdTQ05a56uZbSKQcJNN8BFR+i77Y0b9+Lf02O6C5u9w5yOjZDhbR9RRVAl
VUlgQs+x69QCmwfyeRpI9IUvRKEXg8aCuOlZqu8OCgf9dSF2gMG5DvhdqPvw9QJO
P9Ra9qKmkPi0yPo9Kx0zcrlLHVjrCOkBfNGQ4RKBs9i3JTcpupBbkvcbEdIP5tv5
VH9SqSlYcAoLLQCdhYmGeVMhLyhwPxxvv6kg6LrEBv6HTT2g+X4dVPo1r1lCHYaH
iqh2Np1smKYVV9C+laeUPD6kx32fBUV0rq8XluchhzbxPZstPzdnZ4MVBaYy1QBT
+3NCJhBpXRepcMI8/tDaGGzeA/zEbpYZFp51cfN/tyTE0C14TU0NgkCxoxzBWSxo
4w1leMbJgBmoinMjn3Kyh1bodQ1/y3tM6Py+qvWnqnhpmCiOjxiWe9VCDyfgEA8m
gmq4t/t+w2lSYC/SraUlF6YXIgMR/sk8XsOh0jrgUgeSl/xhHTZ5jVeqSzCOOnvz
at4Kiely1uQ1MOA/Xjf/mnrPznAejZBqh8gpJ9jQ5rGL/Bs6YtVuWAWxQ0uSHc9d
W5M08FjH9MwtBaj/lIUFTE4TPTCzh2Lk2Uuk73AJF0RCIn3g59KXCQ9q1d6YbOw6
3VzxfCmC3VQCrJggTyM/oeg1+hzKUehFKSB7DJMSLph4IzKzEklhsrDK7MYRvmdp
lNJyq8Y2qiyP9FjGd3wBeCyUTdK3vttB51TSlL9JMXuPFZm5ggPAQ2og5qsitN5f
1MKIsbDWhhWgBuC+cqhsRTIjlGeEbx+uggtmTIv+V/HcCN2C7EWCNjNotPXjvlbe
c6WV49aQUkONRtR5xRGwoWaXwL7dHOudivq2LaFeY3QGzpy+ckh4Ff3v25ptDgZk
0UJHnuSfZVLXNZXztgNzIBdRuUllzD+ZfUX0DOgu20VdPJs5fO9VBFrk6T84oU6s
L6xOpP98VHSEn466cBlIdHyVRlKuvsxQ+IQANjnELM1xyYw0HAHXHNXEjXty5YAw
CFsd6eTAm+6tCxzIbItdbubIT2584NJkPkRtIeRG8vQZNMMyMer8ePtg4nvkm6XP
k3sMi51I4emDlBJkz/zQlrG0WFlEMtRfLbUz77i02UKedZshHmfq3hU9c3+1F5t5
p/O5LpH6fhC9/FJqksGAV8ArJFTGbWnqUV+jBZkxH77saFVerr6W87Qs6utlTFvY
rIpvDO6jj5TWQR3khwtKevILaP1IkRk/7bQdhMEaeH+p0dn0APLq397/2Uuyvoyk
FwLxq6Sgr2ksWMEkPbmZtjdhlTsUtqbMl0f42uQDAeLKAjydMNdnN9jBiKK9IX1w
NnoNh61Noihbdz4GTj4vLfC8exEM/78wL5fNR8FuAyk8flGwdSPjRmdKGj01y40D
LMmjrcZFcRdJpdBx0wDweXad5HcUygHycWuUMe1mLPNkaNeevxNxcqp3wnqBQfKI
qu64N+JR0NUg3nD2OespKnrMAh1cj8DgshjnwQyCfOleaNwR1gXzIyAE9++E1WHM
xvuRcNKGUC6kk6kUP5dSKFXs9VxFOM9xChhu+Q1EalNZgnBMdCcrrI3V/2OqUN8e
Tq4OhVdoSBXA1zNXeo1gzdbp/McDgErDMK7BDVcpn+V5kHM3VDj7O8ZGO6rgHc8n
EPM/LEaEV3f6KULdHKAhHeBWZxamFW6xUQJYtCFysWw6nMn6YANtQs5PGpbKVPI1
kFrLepL9BzofFK9HODKJSU9Prry9bRpIO1G54lvKWGDEytXs2x+FnxJ3cvqgjytP
mACAO+x+FASt7oP4tur6agfm6sv/EIwXGc/snXbNAnEcQh1n5z1A/1/VB5sy2Vkc
oPcqQA5qOfur6Xsznht62K4yLvkuViZXq9f2Nr0dCOupqSmaF9O42gi3x+wM1Yzk
WUX+4KZO7JwHe4ngyDtZRGlh/wtG7n2Winunk/8CBj+OgrHiMmMYA5Nz9VYW4qMe
/yAfLreYlaVlibglhxgI0n7lXC6cjtGDWvmykFgoxCeovhkh87kWK8X8udAMoG8W
rKiq96YQ/WDjDqcZcL9P3Skucck2DuJWQF5Aet5o0NzJo2p0Jh8I58BjDeHk6Jha
5G7OW7tsOwc0tsYZM+3TA3bJa7I5GfzTFJovaf4DMabp1TWTM0eqwlAG+2sGP4pi
NCDN0TPKT5jhLfl2DAYtYeMJmvvSGi/Wyqnw3GTXXYvN7AHR7Qans7CJl0t+rwxO
4pEVxR5Per91Ma2w7jc39QeO9TL95agq3TZZ10q8luVFUzyd5Nc83SZyvtW6CMLJ
HP79ZcmS1DJciNs4hrsGIq+xOFM9JvLOn1WoDryn2/v0Y95LS8CA1lFQSVGS7jmn
RRwST3CA9atZwbBeE+qkmyt7BcvZk6BPvQJG0U+ENuFEuznY/GWNNGoqBAOAlAk/
uwpZCkQw+KXP1cLR0DmTAP2vqhNvYX2BKF2FrzeKf6drbGHA1TuA6PWi7/0z6VMs
th3jS9H9the2bDrHHkGafq7OL7K/H7M5elVoSkXBhpMMSq+phVa+CMNiJ8pQocEE
/d6wbobKzWeezerfnPJCwJIlzHiHWCUuTdJSArtrjCD1oj98tG9m7Uaj1CLXYB7B
xhhitpwukVR6kTtmWqvum6te4ncnMafq/fU0AA5ZbQnHnuEdi8gonyyIxcaoStdS
U0NhaYYfGGtvoyW4IXUvYlI4kW/zfdCbiXYTLfZ5IZ95FD3CWcWs+TAIiYbWbUJb
RBtWtjMtJvfXPGMIMHBvJ/5Y7XdPrJaf+m60Vfkzvk3GO9sVuRYQCJ+GVmmSx272
+XbNerLNJ7gRrfh1uq5NhXPLwQteGALBFtSBw0M3BwSiylknzbQl7b3IkwLYVOdg
ffzEghtFH7L+/v/TUi1R9II/nRu8N3OeYKJYvkcG/f0EbKvPbSE+Puf0KEz5Gj8x
P7356EZ4pRp/73t4f9NNGhT2snNz5+P/Bw6Wbmf0R/EiqRvwF2DmsHRDkoT0sysn
y/XICjJ9BbSu5llHfssQdF09oPVcPDwYqfKEo7/KPF19oAZitRSc7aD0C1fml5tv
N1BwLWNE9CFGzle1itAx7dOiRCozaFwmxDo4hmmwF1ykPtDhT2faQQ4oy4vrv0+H
6+G+kDgWQ+BV0FF+S86Rv0DnxBEfcrf9f2Z7pEJ/0IF07mCake3iUY01/LT/67z7
Y/gQccJ16llE5OF6bhPtA6kTvRTB1CDbMLUTAXEugDsfxaF31yhRnP0kael5ucqx
mjP10pVuuOkYfLojEQhjyPSctRFDm8dfi9jVReUjvdcm89+aWGwjbI/3usLQVubb
Gp+WGzWKlx9WusxZhhZ48DbJRovED8IwQHFkyb0ktEQlDin5VDKxxS+M52KWvrlL
mEUneraa8M8BMyGfeGTYWQcoeCjau2bR8JGRYhmZPCWFXfU4YBDCd4r/i4athJMm
l8GAaYnl4/9nL0qQ1yLN0Goxdwh+j7nd7DC+VmfM6lg=
`pragma protect end_protected
