// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:34:50 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A5tNxBwAAT30ggfdZHXQ8T4nNZTgqo8NbxZTbEl/oJqYQz+jkTWklnwie/CJC57p
r6cnW1JNqCvRXaA3B4fFbxWf1nCCIiSk7R/2pXor2Q6ci4vsp3pU4aWm/9wNUpWD
0kk2qYCxg/rSufpcuPnnoccCNY2KPJ5io9siKLYhGbs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 72112)
odTueopi4cQFB6PIKQjVlfXKDqV2ixqLpn5ItcphkqYaw1Bw0qT7MwSyTEhVZZvS
lfmbRzrgUbjD7wUROIKvMD+z5nbHEVyJcOROYIbUn9OjbnkAPpUAlzH7RBvixFup
1FIVS7WLtlcgYiwJdsi8E2YmL9uo3/jB+ZDKCdq895xxWiCkMQk7vHzaD8n7a0Sb
HYjBcSHluWfxO32Y285lYmA6cE+yh6NLevXVFljU/qc8dukdPpMgbXgGshGwhc0+
zT+mpaTHimcWf3ZEj8q3yxLdNks+uacQh6Yn+5mC3rGwQfcambGD6H5oyir9NDVb
IFxbdQayjp9knJlrORgnPtmHVA6LXlCxTOcqCvjgrDMm0VKJnw6LVSHAX+bufcIb
uAJb9FbKZibnQ13dcumY9JNXJeW4MXOQUCqXOfcMoThgwb+GRJF7I+gZxHJrvvlH
AkQtoANXB8OqZr2kAI1be4kp7ZZweYsnYyoPrT+KwWOrxThZVxEQQr6c0DtuZvsQ
7SIkoIVYys/4iRt/36lCIkthJBDjLDl84Crbb/EvJAhT7L0fTUFnT7aBmQyuI6tZ
VBprzDUKLYpYCHCNxjk745+Q31Q3WfgOCG0qPd9JPVJw3k2G2M//ZPn3VwyF1Rn6
QhAbyxCxkzJ22y62xu6DmeIfWDUY/DV8BZEzP8d0X1nJxZo9eHhX8hu4YQsa46MW
/6RTCeT0ruXKn2ZtS4ewH+J3v16KN1GJDtAJZBAbA1ZigkoJW4QPQTCrkHEpDKtV
mG9CVN50xPoKDry+5ojbYkwk8XegfkUEP7aBVZm5JeevGAQy4PeeAW5mWRFve584
MPb0SSBWnfbPTtGOCRHit3i0beD9oDWCVUInDDUXEW4NAHKfeZdPAB42vCG4sLI/
fH4AM+r8aAt3tXUpU/3zWBQ9/wcIzfCgxLOsC/8LpNsd7UQveY0Ejti2Lm0zUxvN
+Uge4sqqt8OoloYVCoQOnroAGEvmdwgFENgtN8sZSW/M7A0xE5u68Wg6Rm2BIuCC
KGCY+my/q/SaoyucLuakx9hEydShKXrtlMLVSqBGYDPvGBcqfIdTLDTrcLr/cRBq
h0B+OLGs7rXL7+8OBacJUOTl+mYP31Z19zjY7smLPTE4W4MEP/bADmVMjtTmjBMy
UMNrTlGkIzWSNiVU2sf5/1QaAtwm+pl1p1WUBSegLXV9WL1nduBzAlGOTmoFsKuo
4uJ/xJxiFEctbI3gUnNA0RaF1MlAK53d3QBjO9jeQg/H/hyowPUvR2fK/BQoDCP8
WrYN63D6mMzZb4iZwInhvcjc7GtrO2+0xW5k+KBPjfgpbeQcet+v7yc1QRcPg4vd
LoIcgVbcAQJmzH9ELejUtvPKEnc2PrXTBHQHyW//0cXApnIBelHxWMlWOP7w1obp
rTR8BEPX583pjdMxkJ6TGO2N+GsJq0n2oUs2Yh5QcXUCs2vF0Ha9S8xA+8dY6Rzx
KW13r/4EVEscNxqbs4qcSKXnN8CgrEZJcqJX1fLviqaS6xbTjlX+1mrz72jJF6Xw
5m9aiTMcQz7D/f3hyeZo6h/jHpo362TDJhhNfdBW29UWwTHUlZfCPlMGbEPu6v6m
2mdpdMX8qvMK0K80LQl4nlsRlPscAMT5/QnfyRDUN4+Ay37n7hDqP7eWdYfthK90
+wpnI1oMtMzAbqvlcPNtYodHMWLXwuxjub7SqwAdYNS3yMqk633t/zJ+64+qO0lE
HbEOEwZe6n4XV+AD01jVOwTczYAAHafDNK3yDF8T0ad+iXdR/rg3su9nnzbVptnC
qd8cWLfoRvQyyJytTRIkyt5e5WeP1lY1jDnQK/ohLESWeo38lkROxTsYjKTek/w+
Uwv4cL9Mm0j7R30bb46XPFzMD38DIfdN3FD8ulLkro7oqI91LTR3FtrK/xlTQ0A2
1gA+iiUAW20yiY+2OklwZQosKypNHkcOxqonctTSocp+rV+mo11iNs3ZdD/6tfLM
T622wjdTXynK5Mm5VxpYCIEb5tb+1GGx0D0UmV+klkdsIJz27G2iSqe6JoBNQEg4
3YPfKMHslYabdXRZoi7oONgTFG+x3g7/DtuEsT+IOn2oEHGORZKcz1Z+UyX90Dyn
/xwcaedscjMhtf+YIapu75Vp5chC9BBSLrdR4qRt/dTru8IuRDZnOReNmMAJV/L0
4n4HudS3cFWsxclRh9Cyz49EB1EMaQUTKIhhg14zvxEKzjCcVk0rb1hMt4IJ3zS6
PHHrBU7c4dGhBu+2Xzhc6BkgdmUk4MK5mZ/Xm0zMRWMOB9NlssxSdvxYMS7guVRd
J3aw0LFtvVqouxqNLZjjHTS0l8I/TA4o/4TeHb9EiHeiOU4tHX3iJNzODMR8zf55
YmS6hMOzSzT2iID6qegS12/321gWndMhUCsU4WUuf2K4z6IDSb7cLx1PpcZNwpP0
rRx2J5W4cRqvaQCIN4Tak08PjYWUNm4zEEAqQyoVJE/d0d5/HuDR7ely7i/xpmBU
unydxvWWeP7630gaJsDiWCWhbL9lZcv/YjPXFqRkYcoWN0mR07XEK2HAr7rwIZka
MoMVSIRvcPweYGuqDZpmkTsItChfITQ3peQ3zTaRQIXJRJ2wGsiAEJfHFb5v8XE1
nDYGyWSlWd+qIivQxIXy9g0mbVjzXKTGpwstotbEBdNcjv8yQVCbC+0dWheZGXDq
PhAalQhZ0sukSiS+d0fznBIGVVHj6nPHJROUtPTeKLBpov0ZxmxSuDJ+JYPqzQon
5aYtavmPAgyxEs4D4l6L/27m8c4B1kvAMtdA45TnSoPYI2VqYmKcZukLHR22z9Qy
9uW7TpJbQuDdvzrlqHs6y+4BjHZ2CdeHi5hIauistQstIJsUkcJzB4j4E9d8z/f6
Y05KXiWyg1Sv2FkOsn3+3MT4BXQAdrwHydI6SbOlv81cain2zi5TErdlrwVif5uu
/M9echXxdGsqmRfJpun4cLqdlVdSSqMNiFFBzyjS4keGYk3fWtggY7MdIL1MD1+J
hfOOUHOgqUAafVZ+vJfIeuhZGPa+aXmSrCPzkca9bVsXaVwGJE4376zbtzVzTEZo
qkhVsEo94XQuX+mEPJtMHztbKWq7id7lPN5vKAuml+o245og9ZzSNwbJ0wsFw96a
CAz6Yw7MYcNbkk+lqiNA70i3HnUscGlRUii+x1XK5Pl8siZmZxpQ96MHuosH4N7L
/Q2GdhwHuWAmtB2Qxtjt7xWbBEaKuvp25hbXQIV4dtiTEgi++J5AOXPouWVCA/eO
V/cifeLEKKBZmUbP7JIuwjNQ7uhMfK7JiI90bmIX8Q01yOvxE9I6yzqDW9A5XGtS
umAtw7HyRpo508tvEdCYgAoj6W1yKjCOTOHRCLq5/7NcqwZep6HR3FB9QvuUx8tJ
4bvrvkxR+IHQCvB/PXtxUxRDystFk2fP3ok5GeSjgO7K5RBGfYWZtEGeoJPbcp7X
bfUFe3EMcvngZvUJQjVshQEJgvJfuZFlTcVAbKTSnLkZaOXiI+Bizke0YZ0ulvA2
/nizAwe6z4MbGoz2KQCO9tFbxbw4hRK6VO3X7tU3xcParV/epdnHw4Xnxg2XJkW2
jKn445zAboWJjmtVgFwPhnrujB6KBT0Am764pjEG/mAFBXEI8J59vZMkvV1bEFbp
yDUlcOHNcYKoeViwikUW85IHE6qsPIFpIhRkRL53UfD2SB+Duw9hjxGkG7+k1o4D
l28thPhgcYA3XWA57X5eJfxTFEPFFeHsRJ65Sz/y7ssZ4Y+RUWy2QDOTBQuECP5l
asHonBhQGxaLIW+qJ1XY4EhxgrnR/QC/u19YjLuHkXKxjDHYtfgqC4jmWAg9ADXC
NV1r749Coju4MkG+Dm3HeVwKlfZcAEr1qiqunevV1H2hBZvSNBATzBKPxulhKTub
BqLNARs+L2GPFhBVyUMxDs+9ZHig1SSsc54XRbCk63viyW5udeltILYCOKrgxej/
N2NQeeYYctihXZA5k5Us5wnILqQ8E/krrM7vgFUrtdSQXCwR563VRDSKxrjAV+yU
PPQAH0gNxj1wwyUT2S46CsU6YuIs/J4aUuQlgh7gCTMoQzWHJkjE6USEKxueaNZr
MdTATgvNC4goSaElYzOgAfdJQJ8tX5AiyoMHF4j2uTUkjn6cYJCBfA0c2qce2JZL
cVGgZEPMEk9l0V5Wj8p0yEX4gxN4Fd4wbUVrWEmfYmxJ6Shuu/WLPkLEglrYwdod
FsIiSUUeWQ66T/kPuAdlNnD3g16ZC3b0TrCLT+EEpHJlytf3701BVOmLl8dPpky2
mUei07og7kCBamFCkOcVuBODHb7T2go0gIwRKdEtZ/ymhq5muJLKzPxJmjwSzhhY
ZaF92Wv07EzWBZtwZByUXU114Ux6pAVueMjZWa4XiLiqlbo7o/OmDswENM3bkZ9j
ld+P+RQLki930PFVRnoRdJZHC2Aj5QgK7iTioNbNXt5FnoDxFtQ/SWQrRCHT5FRF
jTveQ9H72XodqzyYwp9u2sZI+AnicGtK7milKWRlSaOUXd9Wa3ACZsIAEizOfG1m
M1+Z4zGQfW6ZZvNPOfZ4TGgMhMmsz97g24d4dptS7VW/sNCl0+uzDBMteG1fOIVv
t1KOx17ZIs5yAwFhJm3y75WPkc3jSi+pczh5dIwyERHa7nK4+JWkc80crYGtgRkz
g760pWfBRbb4l/bBBwGkPLzwbfD+a36/Fh/8GkO4ZVREyE7LWrWM/fiV7C4+CNP6
0ERt+a8dhk6Tffo+Hb7bxWpaw0fgt8SMX3r6+L7ykge3ojP/NU/SnCxXAlB+KZRe
/1RUtqwN5N0GTUKQ8LJwCzjdFhn/mu64pFv968rZwHO3f+KZexq6zxYTaIcXgLQr
DDCMUU+NesWpGMWEcrFXW1MMsrrxwlDmmTccUuoxdOhVwmHp0+TH9PkV/SFsw5Ma
faJoGlJQPULzdp84HHCAWJ54xMxtIczF1IRkzHRxNaHCL0Qatf2VrBq/rowyvo1D
spPjch7DDFIddxpGhPWDqw/8yvwzu/iboeX0hCOcTk/1M/Ldjw/YbJ3v3a2ZxTD6
EgJM69nhRcDD81zPVnZ+WmZ0451QJfFXfxHW22iXZu6xlVACtKqWgB2la4errB5b
5KHN30bJ/i30FItRqZZnM6FoEekFgN7Y7d/MyaXi0jZVWqchc2Q+gk7PdsMXe7tM
kvESafxN6Pwm3ABEibadrJEk9Mg/bmdeWZ3n0IlAtaOIqO9FtLO0qLN/LNh1lv+y
xJEYEESnH1qWAkGkGW0+6cKr1nS+GclfBoBS6WF1d0klIMUzZQGzNeaJ9pjrWInf
CfJOTzv9xT5cW3gR6MZpVZbdKPzLuyfZbgzzx9GZNOfgNIMSEdKIyAtASPuLT+uP
C5ohS0FWmJ3DswZzf5m0/V3X3Wy0NAHmnbMIamiY8x258ACwBKhB6T8i9vwU8Z7+
WmpYVq7guGc80P67J57mM4sfKkvLLzb/Kp0alZJG4iBvpNNPk+rLDia11d2NkYoI
kIA7oWODNQoQ1+W6Yoy5uQ6VmPCF/CjJCVf7ajg2zgsrDYUg3UHN+E14zkYoMyBz
tObor9TBnBKQ3q0/jz0dZgZ/u+zU+UXkEJBOTESrWCbX9J5AGLTtiaQ+gfowZvE4
rpKzcd5iNJ5dgE3NNeIldATe/QGGCKAxzJgCf5WjFNW5mRXnnGDYt1Rnns4SGE36
MCNEMX0+J9ajuh//PfyblbyimvtymVt2U2lRqwmgPc4SwBsXLGSfilko9K0Ije4s
C0B+QYIPvOFJjSji1OJagLbvUp23vZZ5tDNawGZXpO4608tD87D9ji7a3hTdVXCv
glIuSojZwB0Wk5G7fWQjyX0qwfTzqEeGLsPIIOSB5CrGH5MevEQ8m/dmfqig/D7H
9RHlLL4HiQdWnZNG6wmYc0RLwJ2wHjWVYM69hO7kCTjGN+4kNkoEvWY7WsCmVDWg
ufd6ms8Kpow6ksUPpavRak2g8ZDTFH7OJ8WSpTwPZv/T35J1RCNhYQ02CvkJB3uv
Ja0UZGssYOBu86VjNoe0Bq9s0ucnT8rTTVVwGrOWXirmoXU2LOYfN+iKWo87mfM9
q11jjtR3o9NnaaAMvm06fjwGCD8PIZT01BLVoDgjKvg7V3t+JOtp8gOZkiImccjO
LqYZeJ9flPIpxzjf0BrCQYvBp6yNXmQd2gfBxEe3FBXRR4bnDxUia3GhqfZOR34G
jfS24e1BfqQ5KAl0B5OuQ1hYY8ccp4s8idA2uRt6m+D1zn4/2u3PRCiNfRITNgOo
1bolHYVAHfXQL90i2+QbPjPuG2Jn5yBcSjGS5xmeZmuqMDFfAtHZqBFLdcuD2TAK
h8uphh1PkgclRWz3H+fDVtsZ+n0exXyEKt4eyhdwFkooCbrif+d3zCakaE09Lxc4
JT33rtbyKgK8KDlAgDzf8af2H2FvPSDP2rLAxvx9xjBjZ1M5Hu+CAosXGQEZ0x7G
Th6Iv+dIlVanVNDnn3/DcbTNjc5u16snCcuCFl/zl0DxH4fLe02DeWjbVeraOpAs
pAX23gAeJJ/Au2cMtCosKtpMZgyx8i2XSTUtL8ezUQvStxjKowvII2Yr4VZ7X6Hg
DO3tMy4OOscDUViTqiM3djTTp5eSeizsa7kx3ATY4Hbxc02zzQABpMflsLX3vuBX
Gg1N8zlfU0f7/aZKW5ciUcS+Ehc38NQ/aaoz9jSely2OsbyRgrkF8XSjLnKTTdMo
9BeAuU0n5CDCllUlgFAq3B9cIXNGPCdjPm2Kf38WqK6HGYaFJAhN3rIM0I/oPTbp
gawhoieHbxT2U2I3Kq9d//xPU+rS5ITKtO2kf17qaznmaSgjpYOwhYOCCLmPOoki
+++D/AWPMKsPlJ2rvgE1sgtzHQ3GXzJMV1c634E54sO+VVrJ+wY82Djwbed/YeRD
zEHJvE3iB/7G+Ecbz4PZC4keZ5r3GPXMuc+444zIpjr2VxlcTsIpwC+F4JYcbqZb
TgGKETqiM7HNAlk02iKbLducVpJ2YL+z+kUMT5qJlG/tJq/H2gKYnqEf3Ha45pNO
suPQnJ0rB0FQwKwGcH/TLGmXFjH+tqUir54pZV6Dq7asOYAnk15TsgyHTgjsvHbt
1cKFox9SRSXfYKZA2y6EE/X5gnC3/7vV6pYBJBHCrA2bmIKH+Ws3HDUQveq4EgYd
ZBj3LWo5y6ccJZCgIJiy71QwQMumpUndiGBXbxqjCVhG08OK5HQ2LBYzFXQBZ0TZ
Yod66edAvmExnEOIoe0thlBvxNXU2/aTNfYAzJ0V+VghZlO5BfGrSj2DRP9z4S+m
Oydc0PL1hrf8aWbRAnkCbkhWiGNQQZvmIvjDfuVH4Uk6SarRojfkrAIg1jkcdyhf
GzBz1LZgOHawUGoJsuHyRlu8xu9yJra3Og/cLhZK/5s96PczMVn2PRuGlqikkgC1
wJWkvletY8rexDNSCU7UPrSkNHAohnfeIHq6e2kefIPjoHDCyANa02omIvKgV9IX
YvgPQIhqamEhTVeqysqGVVche9tik/xSXxVz18iEiXYMLfW3iVUi0IS3Y90oTA2R
9vOPbdyUbir84mVEUZ3cXQimVlJ1MiIBVi6xIElWPc0wmgy4dNaAI3FiariHHkPk
fPgvU1sHzHat2tk3G4NQ7fbW+4EZLSdubAwpMa0ThutwFAcj917Ju1kA/53zc+kS
HOjc8a4BHW+kbgp0Web95WnjnxfehJ1TtsMM4wgy/OwBTfMZdQihWCKmJi9z2lLB
csZuCJy4ca1ggjSfFv0wOyEqcBwTUx4Vu0Hb/gtIPUFiDZpRCo5pPi5uscmiLk8q
nl9kXSkxDGzwCnPR3soFLwneKhW94Eq2l8BFM6RozUpoVDpFK7SWtP7SD7Dy5Cmk
tzZEEEBIeUrRk0BvLyYOWHYKVA2F/vuvmZcbTqSIyJ09W0pwvZmyBdU0W2Rro0MG
ApnDfq0jNR//dX4ZJ4w5rIJjVImNMz9TbEfr5panBYqeDWA1K6iDSgMOprm2fikA
YQJNk8ItmTfup7P/MR7vgstgOXxqzO9J0KjvDfcfFgNPErrsn/vSPFXoM7wIeFz4
VYwOhQ1ggYwZXoy+UCGfa73CwjIJsPRvh/JED/HJfBbRhPf2+U9ecIOK2HHD3CWD
E4dhXhLWQV7+5A4WljTmQQ5/lI+XGd0UNY/9YmwjGUjNreIaA4nAFVH3ny0cdnyQ
IpCkWn5/aymZvx4QhxyyE1Z5AL15+OAB6g0Kete+OjkzSpsv+Bm0b+bgf/BdWs0u
LI/5xry/ic857qEA5UAtMxEwp69u8h/fK+KX6Tyk5FTc2ui+el+UV/Pzg0YCKFOs
IQBO29nXvskRnPtKvLQcU1PEPqbB/tPZ4I3P9ifvYGz48E3u/Ly/6d7fzeDO4dNC
D4aNJae5DVQQ27MNFNIxCxrVnEX8v5qOoIHhAQqQ48lH9fMByWj5JF3ojyXoVQOJ
/46hEv8agFbDBDC2MwOWNcFHAmiryVeWUv/1VQeCFotVoYlS5QPDJez9N299v5uH
s8FQGFCbx5xB0TRozUF1WscdjWv9QhIZDE2u6HEHBh3qENGXR1mkdDwGyRArLGjV
S1rBYeYk7OsKh+WfF32aS3GW8n8KHR2NSqHY8SF4vgKn9zhHBS824r+G3Nf6L+p8
tIU39ymNOeo0/lnetnQtuirBc9ASt9xB9KB7Lo8tV1Npa5suYpWzhxRip4cIaE5Q
e0ShqwcyG93WXUyRvMAnvWvd4U11HT2kPNcRmfXqZ80bzVfB4XnqNlAmliWKlGcc
PDTZK5a/AZehY8H7OYTo5o12HQfIg1L01kQa5D/c5bd+oW5U71aOELYMurbur3+c
im9BAAEUwONT9xlIk90XxroEjwZ28/KP4fe+f7safgUBdA76wkQTHvcOnvDzMRLv
jtIlyS0FTkoG5W7pfMT34x20PTqvDpizcY/qldCu+KaOJtUdBD8/GXFGO936rQ5f
2DVgdaP/58kXaTqPYd+tj+4MrWtSMkam/mwovCOrTCc7Zr3XAVwiI6pl29r/5DyF
I7SfUsEeSdopp0/0mmxY/1hGjCX0wfNOKkTcIOXpPrBRmsDeiu/+yXYDLvfvk1Ep
WfkBFhbBEEZUXyL943D1HFThDNj9Zbd/FJnC5LTY7R8A7qhFhmOqLIBGJu6yP8fx
10ufalH87j0ewe60p+hiob1QmPbOfKGkmsNZUqAQXCx8ZPmkP5kre9+2/5+jeiyg
KAhMwOTUPVDWASAGuSGE8bzwPJ5WUgFlBTIjc5KkrRhhLo56rWEuhWj+0+MVJol6
CaRPcJb6nOH4ji5pOPBwb8Q5fFK4sDSJ7BxBJC3OBqm6sJ5RkCYxEqCTEk+596OY
kNXN3IfB/2yaqgzPK3OUVts6lZzbLrcjkIDXOSEi6B0zMFghvCU0Q6DVT6s3nLnH
DOZAtjd4flsC7HhxC/5iy3DZecAgZKJTNIC30zXU5IBHbTVMToHfFBttDKxUBoeX
F/YCpk/s0pcQYqffUQplrF4Zj3fQxZjmutS1NFQ0w4D10bIyRhJHwyPsvrcSifYT
7Yp0HpdSs0PrCIQzqGFLXjPerkDN3nklpJj1k54n9oO2fp3ci9Buzi9TMXt6PePb
HqSqM982KKqez5B82Rlnqv4aYjP0wBSe0vWb9EzsfTPyjydiMaiTg0KXMQLeX4mh
SQfhTIrvCekdpatSrx3hZOTFD85YlVNO9rMLOP3JH29RHdyT6wlHwWaiIy4SCxej
lI13Qv6EiTzCiTI+HogAtVQc5IbLYC6dFVGHqdFOHKsGcgKK6p6LBo4E4G2o2ejx
KaaXycqYZD7pEQWSi67+K/0cfRFRadluRmKF53ZYGw8GzBLda4UYX5WjAcVSPNpI
Sb34r7HSuYx/ZQWe4gC2SGLLRByMPCpJhMahLe16bZW1eGMpfM4xiceqhzu2J62m
nyp05/6dm1bS49iwOo9cRroJ96MJdZU85t1jmSVaftIVNr0X3bxyAaK2yA+z2FUj
idqRQrHiDsnmVfT3wsP4eukFrLUCqq6Cw12hWETPnldDPDnF7mF50/S04rCazPLu
TJ663ke69A6JtA8j0imxEVKfnkQPU9DIJzsJrlFLWi3m8/0mcY/5dnrAA6RrB7x7
UjjsMza+shmjvtX5jiJ2krT2zjnk3EAt+1LYMA4O/uQO0xLQLwuwnlHCaOIGyrjd
booKV9K5I3AlAxv9e4apq0kWQwqU9hdwU0pqfk24lqYsSCWU/v6oTvrXJLtwlwoi
6Xb3cPnAlWRQ++BjLnqcVK34AtuKdJ1+o9ayau+Z2AZLfqy7w4iMqW69PPOU5nra
CBbqk2ius8PyJkEE3wsl9KkfwaWBqgdwJR879Y/RB9DHtGHxe1UxCOIVm4IZjvxi
p9Vp4l9oxDXio/CozUIpTnmt79oldXptLZIBBf2uFkzvPB3sJMTLsvzuuE34D6B+
Bij0oZLrc6vtazS6mLGiVQZfgONIjCl166Df7T76YNjjFQvOJ1Z/UWCJ0aAAOhVV
ro0HAZw+t+sQNM/bk1gUYqvO2ixhGreUrfuubVgLOru0YXc4tH/1kGevGF/+Kvqv
/wktQmVF/Tok10FaxrgRWuFuUpndpZ95bfGf+P/Bg1ZkMRq+Gja1G/ll6tTwbSCE
gZnZ5Wx8ZKWZSD8d+4AanZ+Kp1/kvNmrYdz8DMNdplN/OmU6wKHhacK2myofuLUj
o9JXdqV9mOJ8YDomPyAG9AGIO1SJv1W3sszVAatPGq4gX+18dA8S/d3ZdCFFErnV
Cc0SMbD5M6TW5nFptObtPufbsjVdGWaFbBGjmKB92l5LHHpUeeDhDtYJVNNDl7q2
Nt6qy5IEqVVgHaXscnFz6q+mLzt1tN1FuCKiyLmmluWp6bxurtZVPUEAJMt4bn8U
tBkASz502TC44NjE4/n1OgFxB5wESvfS1vzMJLX7FFCTuxyKMb68knQNxwKKdaTa
Cs+PuI+Kao6viiiERF8jU0SsO1dd+pKqoQ5bAs8K7+FdGdJtnKsU+1SLArsLzTzW
udUC2mtQXXWi1OQ4RS+S9EsLCXx/vBvp5Bp9MK1uL59kSfVG1McqqoagMsas3nFw
VdR9pPcIS+4VTMP5/nObKTYIW6HNpm9KmQSjtaXcsLRmBy9yUsCD4AIqjtYkFuum
o1B1PsNWGqGX2NeS7TxJdEOOSXugsH24rQ+QZv7gMHxZ66dKFlhz8pB2gl7FL065
hx9mqXVOs7ht69OvkQjvQG1W/Bxa2NrWhRo3wsjscE9QR/nMrkuPhdFHagKBAXUM
UWjK9jUcQj0C64+mYGecK5Whf5ziXaGkIrStQxdJ683TfezpueKrr58fJWZHuOMh
YhdlroZ4N2uA78QaiBBiaaJFgs+xLgphtZNSJb0M8p3/C8xhJvOIaCR3I2UyvT4G
3FYs3X28fS/5qsz5Os2ZVQchEIadjt3MObppgoDGdTihjGeS8Qg8BEi4z/d6SdgD
LZHzwc9aA5Y+cylLTZ5wDxOIOlSKjLIFegiPcYz6DCQcylwImVt7spEquW0RkLCc
9ZTfd+G4FW+Md057z5Ji3ot9cjzHUb3MRrcyXt2OUOTeYXDOWACyKOLp4I0DIHLX
LnVR/WpwaRGiNJ3ffxxLnhNUsczfsPKxxpj/xc10ZO4Knrc2+lNtqpkMj3B0kxRB
g1ZUzuZY06mhHVwf4oqG4PHx9knruJRIVsbbU0gzNMrS3rg4Vy3L7DoIUwUbs6zz
iGbxjrWnS4LYvAr/PZPCHlloW8Gr6I8s4+mZkgGuvbclWgQsHRy16ZULz2xzLsyB
rIcaepuX73fm1O2wfb0hh6/tH8rjecDCro0sr0/A8bD4YGEml4N6KQSWR5bZH8Ws
Y18UkLyEIs1U6RHuPrbIzz5uIkjI9iKVmbBuC0zaJYaf3I60vEFPbI7IGBsI9S3y
2D69pvEUSHz5PiBqSP8VtlGuG+ethBVJm8d5biCD/pgPSw/P0R37xtTw8L87kr5Y
pnCpaXlngx3dZ5QFed6Gz9a6ODZzBELO9GdeChJaM5wF3CtS2PnGl/fK1ZbDlo9L
Eiwca0kJGuce8FHaYZNyKDFEP25xBNph05u55CIFSz1lWi30FZATOPSt33eML6ro
59+wajaZv3liijGO6LrJkWpjBt12c7REFIXQwWa/8Nn93Os22MGyoWap3pphFo8E
h0PhP835k0vFzxnJ0VfeMXqlW/M6Ga+8GTO1+Dlmsg6g3sNdq84/A8WHoU28+Qvo
vyqMjlQrX7xXAz+SN+v2KqGOrmB495EAUuJbYJu0V76+WkyvKQQsimOfWNYrHZPd
r7PMhCL/as29pzn7Ow8DltENNzc8/vOWcbhAuIXsUTBYbkLutMc0pwctXLVNccWf
6vZty98WYlte6AzFjwFSE5DunXJVH/HqNz7fli+WYUHtogzMtcLJrH59S3vIZw3v
IUAjaV/XtReYVHxnNalCdVAIVrIqlLDVICcydTvwNJyB8tvXE9yDtUuiTU5WQ2wM
OGtDbh4+jJlY6SpkQ9SBy1cPjSfscrfcRf6T6udqw+7BqK5Qo2DNYBHDvVhmRMBg
MpdKqqnAJwVN4DxknCO/aO8+ZPm0985UtaxIsYubM5ktphpEPdbu5PJuApzlayc0
Z8NLpwgrzo5aUcwQfaacoIpWsNAKuRBicVuHYKBjBDWpGfyWtl6lWRdYQvD9bIR0
QFkBpBnjaOAmJI8JA+Q0Xjq/qRDiTuLph476BDA43j/xCMdgkrHiaKwB29S7CHpL
U5EpzZTYP+0p2Gc4Tv5EzZn5hCTsoRvt7kITcDiYO/K7gP+6a3jP8Jr7tGEbIC8I
Nm9kpY2jLVf5gyx1jBvMGGErQ4LCIcvvo4qetdwhlPKXTn7j4GPThsrqjT4V6yye
GN8iCiMcv+L9nG0gzXidKT/azIoDspgTiq7x3YytUrqRB3vDkBi+Oc7eXzy8no3B
Zo1P11OXBCRbUgD+WoBS5XftWnBA/fG0Tbd7kaJX8xHxuMaN8uBRbGa4VSjZsLG0
HWfTdwsEacNcr+EY5wm5c1FLvFtSOjNe1dWVEylTH4ZpKDBadp3Xr6LyD+2pg1Af
ccVHJ/vvUOTrEJbyaR5iVB4hU69Pghs/vFgmZ1VES9nHEfwRenC98xTRCCY5dYDJ
PbKm7uIF8v4hvKesWwOkqV9jjQVLB7rM5NJyrDEEQlsVEfwIEmenjw9DR0KoX1Ej
5S8F/0UKLWI2GGSm/B/nWcHCdMGOlqNq2hjEuEtYExtnUWBiLhFFim46UDTZ//+a
DUtDNWKNhBg+xmPkMxZjgaR0Tfps+qRbRZ/CgzSLCMNH72pSgFZOthWGLDEH5yKB
OZ2EuzZe/CyfCb+QhhsTc7EBnaDAmzSgl3bbiV5gMZB3KVIQ9CII5IDTJVuorMu7
2sja4RZZPLkQL3on7/uhZm2zRUTrFChoF2Pvx0/unx2WuSCYQ015rKRH2H6bISz1
W+WWJuHVy2sO40GcaHTy0wPP6CS/mgX29uGCMYIS7jVkizHZYxcpX2VOtz5NEUyg
YRZzOT4svPg1EAlPRD9z2YYRZFTtxBzQIMFEEgKaXovIEY+4m/jN6gpHA/jlAFaZ
pan/K5mOOypMg1fkzoUWsX3Mu7lwMCdM2P2WlGwdkkHxgUGP4sziyBDud74V2IUP
rG7jlQUABZB5uMtOffqGHZtCuHapgnbhBv8V+lL0DZe8KiDHhbV5h2oDXkOlfEl2
LbdPC6sVLRoFu//p9NFtUQ3ZCAW5uD/d8aan0McP4lrXGNI8BufYsp27QdBeWKBr
mwR0n4AUqCIiz2rGWYC4ZNyiP9NElVztYVvXF3M4qE1plhH6TKYmqW5hpXxU2ZrW
KvRU91r7YU5Wt047fgYidRCiYnSG3ZqNJ0BKN3ZMvsUheav2v4TcS1j/yZg5GP7Z
qS/HgD+CEfDR1KwnzlQI9Uphuh+EJWFGkMuFPqGfPtHJIsY07vi2PJwQ2jAD/FdD
l8fbfj2kBnluVpukmjJTAXV2wYK+dNiVyMdFrmioq3ehr6crtKQgwYWIqPYg3s5M
7uOBgYkkXhYOVxJlLBm7x/Gyt78z2TEoYQdIQ9zlOmBPGImGbOMzQYU88RiZYWbT
9EQHyp/gjlaHw9oY26YACxjBz/RwMi15cF33+jhFygGBj3qMvfk4W9fIPWKIo58c
qggAaaOSWTbWx4tmgiY0c+LWgkoFHP5RHQhVNJusOGbEqltxN9OBTg0CrffAK9cB
Bxs3m5ZeaDB3Smj6/UKB/h+2sksJV3X7H80Knuxhu+cUYkG8w3h5t6vH+QtopIBJ
UfditSXukiMF/l2xdOBmj73oCn5hY1ERKaWIuk6uCBYMN9LhcWRx8Jgu9bIIEAnW
/hmrvIVQooma7uErtyhD4bqXA7MEZDqOk55XnVHjsz2I5HF+dCdwUSet4sYKJPJO
lpEMbVJlQnAYS32ciRVxq8k8gjHf0xX+98XX2wQV4kKJOZz3FYckO8fZfvE5ZpKd
9LHululniMJI6KkfxEWKVWNGT5366Vfvyr6VP/PcFxcK8M8Jkzo8SxcvkosYUs9q
8sQf0b9O8ESqLLV5Gfp8OgSESrc1mTT93qKhJTZ/GcxE1Z8xpvllfkI/atYjRyz7
KAEtXW15MnRGdXQ7kZztEhmXKfGmHilaucEp6oOs6yy16dCNpDXBe9CqdEQyIbgC
lDHa6vtdsc/WqdSjbLASOvJZkqEeXtT6u3YttCoL+ly7tBFTXdM+H83ZHiW3Cppu
//GT/7NwYOj2t99+1hlOFkBI9SBVYGX83/lDQ/g1CHGghA6q7W5XK/y4+opjz6cV
oqokrY8j4nNIyfXfEIR8qhYnU53qHGdpzRe/ogMGCHV3Xdp0oxUXmpysqcJXySyH
NqekoV/lD3QYsHrM2UGey8X/VKC8usN9Jr7wCGPVMmex/M5ctzuGW7bDZvb+OlFI
A2JWAbblWdhS2eALofvHPyUBP6rrFf6nUNtmOibYouGRc729P0CSG1jZpUeZsLu1
+pkeIba37LirOyUYyEJW/RxGcZ7KfAmusIqrnGgtM90toxcHddIlW3QF4UR4J16L
EZwWvixhSUL7FQx1cIHw/bhXwD2Hh0EaY+LL/gQTWN90ikcmM0B93znvIGZPee1a
kIpGGqpSFytBM/sTqSkKoMAayVI1QyYukrVuX+VhdMufck+Tjuzzr1nwWIu6D5AS
9DwG1X6ho4LzTaynkGohH117AuPmBowpF/p++8Si8luVO1QAuvsjMlHce5v9pFVA
9GhKI0eXFK2nhL7z2aR4pLAWeVlWI///sN01CGrNuGRzoLB3wpUpf4RlzlFGGn/1
slRf1ZgA5QxaiuXb1TdfkEn2fjP/ZEyv/w5S7xdcf1W8zhoWbI4DzU+RHykFlR3t
/7fANVp6XTdBfJwQV/6B4AqT+XvFDgrA1ErCnvGXirHwz0ikep/1SuTZK6K1Fzzd
P8xvYXVpVijrFpecdHxvaUO2rP2MwUZm/O8a1KykPS00lsEI82c8jufURfXrC1XB
Qr7wG71hiDY2bs2lcEy5zQAvVea+xOSXeLUX03yYQPHi2/QNzJMzP1MbfNzHutyt
nM7CLKNDrxP+GSr7AHkhsAllc7lErP64L0G8YZj2KBkDunTPrBXAF0nX3QKbtHxW
yI7w+XMiGI8WA5wAN3Oa6jSShw+9bMGaUIvjFmSTHUlZkvedrU1wPr0Xqz0xda3P
/q2gNhZgHDOPXFjzBYYPePhLv/bUnN8S+A3O0tIXLW+jlWWOgm6B1afGrUnSCvh4
5llSVY/U8qYOmMmg4j+0RrRezjR7cO4T3RUmKLVXboJlyVjA3hLkQ7mAh+XnmaIN
Q4l2nX327L4qWe6fVEShamHz1BF8vb7Ekxc3Uf6Mo6OGecaJlPlv0XnOy7A6kE24
MT4+HZ/xyMiAicbtZFwWMW/whM3WHCRMeifD6E+lFQ/iCr4OB+BQ48bAxA2fRfiG
9yRtGmjm+F9L2k+oIe/jb5FcHnr0WvdlqFxZXYT+LsSycqGSxTV6bYvMWoeRqI1Z
Z+Mikg63fRTDNSmG4RwIs1YM7+x9PA8Pm+u3h3Ho2SxVaTEm8MrtjLlcEGp/o6bT
cOHEVoil7yPKeusMfCXVxgGwtIibphd8N2xpczh49W2xMLO4+dGIP7gMH9uRKAZO
SW3QDz7tH2ejRsCojZVPLk1JLQQZ+EnImpKJXLxLNJfGvWL/LtW1/IuGFgYGwl6E
Ma50xFv7+P30ziOXEvk/YpckUEZNpwjaZWgDqUFPTCBk7/fRz2xo6PyVGL7LHHpn
MF2DIl+X7EcjC22nsW9yQcDKLeyN/8wgtVsr6G2O1TZYyEqilhXoN0b79NM6UhxL
YBFz8E0pN3DfyfzLlTCg7D/quI8yEOmZiuh/OkKAJrVTPR0d/oiDQSZUL67eQEBD
yvyM0vJe4u+mAnCmrHornckfTuANRfUTa2UUhm/TNTTDJyQB6GNzO0Y5HTT34wl8
oyeJqf120LHd9hH/YnrgxupjlkF4lluWC219CXw5YbaNj6m81Ne/8Sqp5H4bIByJ
XPJpBnsJ7NnPnofqdgOhAwWc3dOKbpEU0iyh7+fwaO1l7VRssaqUjtv3yDI3HdU5
qVG/85Ph71e1zWw6WA0rZfsQhHN3Qj16aGZdPByjnhqmfI9KH9+6w7/bhOu/pIL1
ITuNpOSz519Yq+nBJoPs+P5EaG9G6i3B7+C5InHRY/aXTqHIFf9IeNZw38KW8ZES
nB+RkXCXyb529xMgIQwZdAbEGx2+khYrHhDMtHLLfQ6XFn+RC+2+WaXdDEPDI2CA
DwRyUEQLELnerN4PTW1hy2R0uAUsr3VMDZP5LIQoHOhcIzk/3FHTH5uCsM4c8s8p
aUepjExq88lCkqXm6/B/mz5scQ+cevXN9fT/lM4KZBiSwckhtv4lMUarRbJULQSf
6ydepIfOk9kGHaf8+eVsjLVeLbZyCCuYvvChLlcXlnCi8curv0N20xk2ddrAhXZP
nKLwt6wmrMKs7EvNCxvdKrpFjC9saOMKHJKE+M9M0sWVtjxWLl8bw0N0t0HnP+Bi
equsW0+3qUXgkJT7sIfEE0nFxCuNVdMjipajhrDG+yARYp9Ln/5CF+BQGVJkZI+P
CiZEwHthw8UtRhTtGlHN3C6MMs2uRJ+sONO6IUyDSlNylK78bkEhkPOlLcsXYPrU
szSL5XTANif+Gq3YEmmaEu4FbVmG5W2kbZ7n8Bc5H9VvNs2HeiCh1n8SSIvv4kLb
Y5cDKpNZNQzu0KXDmbrmWqq2+2OgPJyqG2s3XG4ahALUoX/nf2JBU98hiGQSZsfg
lix/1fixXqA21+7LFGy8D6Du8/UkG1f7S/2PZ70BFNjhFT8UcugSHcWTLj5S2EHd
WPGXoydo9B+IoQcUx0EPd7RlJyE3liys8LVXi/hmg7vxO1rhSobLW7OSxY47eOOp
RKnrp7oxwplGfBu3/dV6knifj1ljDs9Z6EKNCs7L0kNLXgs91d58Pi8oIoZHZPKs
BnvgEpCsRWqWr+GmFNd79N3tgl5YprEl8wj8iwnzcHRuOCY2eQUpk+ww0xp5r7Pk
BSvPkFWwZGnpb7tmYEra9J2wdM1Pyc5zVni4zb/VD6cU8nQo5lhvznAYXk6FlXpC
TQQ9PdA1mgE95JCsBlKTHjvmC1ZyC9355SDybcdvX5iRY1LMgYe11QAootaQtSyP
8+wMgbleENiedAUyzs/XJM9MvBVWBTlNn9OEHeWNKpCrKTcBVCzl3lz6rh3SKpgX
iHfKhTT8QX32fQsckCkf8+itUYK4pK0PBiPH156UZ3+HWpIe+fAXCKQSlzUN1QF/
Cyx4MjThgTMeTyl/W1VH7x7tvJa/PRBdH8qrUmvRI1r0gfqEuGOkU7i8PqWxQOk2
C0YM/vjpY2O5+AAnlCi0AaD3MO90qBBth2RzJKli5ecmq8HypwiZS7Us4igEgNlU
ER/dbcRO0GAQhhs5Ko6mU5qHplClGzv33vpOBWjqt19y1wdikOavrHLYxiqqiNn6
u2z8GChuMfm7sJQarixtRFPKJr6ZnWT7iLSOSIoB2hN1DJUKf5W9zAlu79FC9IcC
3Wn4IUkbrofOvsMebYwiaTQJW2RLW37BulWAwSEjJVya1SUzGQP6VsJslKnldv0E
sosj8/5zstPRwtd2oDT/NWsJtGWxpMBO9dBV+MJfsVt/P+BYeNZDmnuUQYPAf6YY
9yUBocje5WcQxOewQ0CIqHj9T4PaR4JY7SFnI+A6n/QKjtnnOy4Rg1BJPAPQtohf
plrhE2ofYKlaafEwyIKUYo/bVhSooNKPdqkhHi8k40ZzU3cOH0ThS9DDygecvYS2
2ysqs996hlJXyl5YxjLsBwFdUMJhnH101WrdG508ML5VRz0PulPyC7bM/ZwoZBXp
B9SwlI4s1JKBilrRK0LXdOWw2c0qRwO7yW6o2EBSV3wdbqSsmKARBmEEiBKX3Ctd
UA0P014SC1E3TidcMP+VuGPVLjs5wfDCPkijtez3NpFV2cvcHD6QYpiamhWsdTEX
aIwek2g6Lftfd9uCUk+r3iFZROouXa62+vLC6p3MzsjbF2MCp+MW7fAtUcipmOKO
4KDyxQUGJ/B/Cv4SeHuUXm7SBPDK9N4+Q5sQSNGj44788kDRsrQzzCM+Pcg7d0pW
JQsEjTQTes9Qww2XMaduc7zTGKn6TyImouitUZeT6RSJK3qv+WQGETKV/GCoFpcw
NoQNF91XO38vQ+n2wNmqfrmsU4p92obfZMDbcvvXFHIuy+HJ+wfVk5f+7KpMn8OW
RoBc8jxT67GcSbBWB7Mn9A2McfWSciHYfx5v+qhOdXH8objZoyw95RHm8nm0eIOe
meLyYBeYr4SAcjPWWZhvA0oz1lfjNqQTV9zk6d4gJwYpWaPBzHO0AwIT3EhlNoQb
qKK6F/P9qTq/RlaE6xNlgncdfzVrohWnAr8+sTTsDTxEh1b5Dn4dPDSGrKLqVVbV
4zJNIqQWuJw1ynrQOCKWMfu+G1Bv0KDNtWjLXxSmTqKasr39O55cfIE3iQzoTpkP
JR4GB2R27WmhIQXICBnPk4U9X1JpYJcZABrT7W4HZDVO5UsDrQzvD59mpuiEZY8t
XhUi+H83FsyNtmQOx7SzZ0pfCyesOk9rZNaBoKPyVny1hQAsqRD7c8EBU9L4BW94
W62+0eMYSpwGconpm5KIY+8C+c5j/XCV6sT5hP3ZiVBdkhvNpSr9Q2okK0scRBlt
/4guS84SsvXLPh2k1OWVYRoS9MMX0BD9F0ZEhkfhmVHMkQMswh976bwlGG/CWb1n
RN5/5XbJoqcqDLXKQ6g3DjVmpw/57xlGXCqmdpKC53rqVdV38/4mZGnb03qtXAHw
3qYz507PIEZq5Yj6n5cRiOlCN3uwg6JgKhUVSte7Wbfl0RdJVle5dq+dT3utVd5L
XNcTGn9XaU+irjsietur0rKvqizNe+LOfjKg1Qxjs3f1QcjvV/p80Yv1E8oA58Rn
f9x1OOvWH3NywfOYtB+fUMBUal7v0KinUa5K0xOdYWo4KCe+FiKREuwPCL8JSR1z
J9eqm7VQqhPKvBL0rrk9vdFpJLACf2hoBfr6GeMbN9V7KCd5jvmqwjNYYxMochZE
vv9bTFH5UQkxLYBqELWcgjiqxl1FXLZQnrKoP31411LmnNrivwOsCZ6y7+OiByMW
9SLuIqjhemXEQvaSxtqUuEUzV9hdcIo4Bf9T9TaqWXTeWAKGufKNxoVElGO5cfwE
X6snYO5Ly1cIWVkWrh2kM0AkHuE1N3AQZyfvzJ+CE308kWwx1ta6NlnmhGJpZbY1
4Qk7e/8iptNwQfPV1yMw1UCRkpKDDRA3NaMw/VkB6aAiewNVMtkuTQm2bROSp7jW
wDSSfX87W1viR3w0lHa91XDgMbcWvhZMmBY/Vj+wTRATx+QFJdTA/lCSPwgT2sXG
x/pl+AAeVfDDI2YYSW4k4zBOktSBAUhZDQfvFu+IDYoyR10nw6vI00nJpg9FSuDs
41BPhQbCTlUu3T9qYxX3jqbPkLsdMIrzixlPe7xpgUkdlcXXVNaVz6bOfHTHxgPh
ACYsBgRBZS2T3zK0JoDue/i+0xoTr21cUwFtiAP0QXEDcDCXMTTSwutI6HTd4oH0
NcrQdt1lp62ac+fJFh0zvtQ/EVu2s/KyLPWLqYFmFRhWFbj3sqP4XPFVSejfn6V3
nzSLSUKEMcyw/RZwFZY6HpT55NHrKK4PaiEs7izm9Fs4isUi/IcGisl3NhGmczJx
oeJ6/inpQN2AZ26smFT7m07RiosnldQpXq1ZAVXu3MYOOxrfpJEDjOiIqUMJQTPq
QlEEtj4hgsvisco2b/GrBjw65ZUy+Q36xyrsFwXqxBodK5ti8tH7uVPO4xT8XwPF
5TSRHMppML3A9hyi++J/WqZwGWcpVpc1lOZnQv+LH7EFB8yuUUul73sC8+zyX3H5
cznW3jy2jaoH+hDEh57iPaxLUe+VD4q8w2SDfeXTBqrJpt+gMR61amvhQQJ6gy0M
E5PFbfbXl1O1thyrLXt1P6JT3EfznDilK1sQl9h9eGi4LZGILk/zE8gVo+lDc/e/
Lbfltrq4AlpQLxcbGJZe1AqJrZ9RLjalxpIMvdE9Jhi3RE3it5Uu7Kaxh6KVGtJu
U+9ygG2FCGntvtgZZ2OhlM8F36N8KeKwz40SkXYXvVVGNjZvrn6nQo5jI5BQUryD
WsvYE16PamBJ+MYvxzXH9ez9Kbg3dHspLEXPtllrkDdGKy+6fiCcRyqIFDGjdYZv
kECqNOlBGCZSveIqJJNi9wXm4QW6qoSDjkTSnEdzJ0g9M1Z649bwl1Pykp7Cl12j
3gdSBLH9kcgvvDHd5klcQiSuPQ9EYzn4EDmndJIQtL8GaxCIIRxHTdAb1I0+U/nK
MvQ49mvg9A6wtlwkO9rlRq9R0qQjP9qSxbDN0fdmYLVdUkOGuWRZwqVZsUtSuI7Y
kVNA7/VnH3EIqzkz/QQ/Ie4KII91VZ7CbAWeR5tZ8sfx0tswdPzouAp5eNXdO1ez
skRRli2rqqRCiKPOwVxYTZOpvq3ycgdryuYOWK/OLpAzveo4kQemktYD/q4SIPzx
Q26VFadD+zQpvn6z+xQsFRBUrbiVzV1TjiH9ZIZD5IbPnv1BkQCub+RtW4N8ZU21
Tn+hQmasI36dMMpi9SLPstHsucS0r2HvR+aZZ16SNFcdrIaSG8NLsm5ZL8aBQjKk
vUyW+drZy7IH9HBmrP0Y6mX4w5sMid6Gc0WcGJSIO1apUGBUE014yY2tjUvZDPC1
2ZiKFQGolj7/5S4hggPjFQnPuR2SiYgFCVSfT06tvD91elEAq/sMB95WHkdd/6uK
+5DzfCgM8tr+dSiMtXSqxqzPTsZVr+SUqvOq0WnZCTsFjzu/ZO3FxgFwuouyIrTp
DC4kHeox6txJF2jXqv22w0sxgh+rmmMlAbfiFERsFRyrzrAZ4htTKQIfZVYJxC6/
4oCvj4wgPLPJK6ohn02zCt4gyycxmfTLU25AKzc6SzetTucUKVpa65rOriUSCu2F
AKAJ+vzTYgqNHwcvwhnpKY+YPx4ysRWoIVqGhilB4y0DOJGkuJiQa+sevQyJp6Bj
y3n48KgspSURG5UhrES4n+4gLJFxHQeOPlv5me7JJm3aJwjnMSwuWT/LCm3ooXJn
/v8xwQkTI96MDmcHJ2am2Q1ge2UqeAmVH3V12xDhx7uQ2a/aT+MTb2NPa5GvLx1h
iz/Koa+N+22pE2jZwxi+TtLj4vcZXkE6XFPn2uz26EGDKMwaQMzUharuCcxW4THc
QNpxFFRTBXAuHMI5w9Xqk5Tt7nbBqT8oMtJeHDnrGFC6ZbPrawMTRb7eYMfOjRNd
pumgVl5xCqubhBZppqtWfveIyMVnYN+JlG9EC8otq5dZRHe0utC42M92XdTl/Id/
UT/eRBlbkmTngjNN1F3jZ/aahoMGi8yE+/dAhak5kFBIVUpr/JFPxzMt03IzYl3k
2kFiJ6XPaLpcbTfDMaQbY0PKd89k59GL6dD9v2Qlp+JeVwaHxuONB/WGm5yAIt+6
PPNPu8468PicpokQG3iobq02NOL5MFrC7X8hr034Qxkk9By4+JM2XmF6IDno4amt
A70V753IITQHVti/XEdlKxB3ez5KqE2/Q453uX1X1uegli+J4RbJJDVuJo9McREa
WN2nBXqbUemzBDfWWz53WLXFVw/VvrY+rKlNKJigAgcy7cyjKcQyTB+QQ86DmVy6
9D8imdyZ3SOj3oFcl9qlY0fqTjp5FuOx3OGRvI+NyIa/Z5FGE+wXgRQV/dMKvn39
pXijzKROCAPaX5wt2LG4Yns/l6bAPXyk099JzQZ68RP7TYtMnPMCPB697Pgfl/ws
z+gEQl3YDx5X83twNImC3AROBEZWbICsLqUgaBG8kncUaz9tFx3uZBEbd8FSXflu
Rm+I81+DpYibu1xlhuPA1Dw939toqxFWIUv+CAi4K4HHxCLbWMblOVrXdY6wzzeW
mTrzv9f/S4dXQAowz0GIIUXoGXwGGjjRgD6KcTUUIC/ZgbaTKFW0+u5fQZgsnWnq
MnXgDp4i/ahHrjzH6BdEsvzVygVPJjwN5n6QkEwuG5615G1KLz9e/3hxSKvHlyiv
+B4QTz+uu9a96xR5xHJAFQQB9A2T/lLKbqcLHFN2BkLD9p6phC9h6Qqxsb7eqZhp
QgpYpP4jUmnm8ssgMnE/n2TXodtYRbcXtdMjSrherWFphe2+Ha822h/Mch/e/X56
gOc5tzMY9IunCJVwyQkCHKB8ZZ6gZF/da9gJOwiQ/Mnxu/5AaqTedx8W3RJojE1L
cTjN8KrUc3UnxjhaeyYdmGF+9yjbfQ0zBw/oxol+mub76+GXtS6lJlyXcj90CGe0
BwLbDj170ECwra27AQxDUf0Zqc++XR36Qh5CLLYVCzh7Ya9F8p7BMF54JvA/kp9t
8pQuSqrEANOLndVDMmiW9iGUNSPv8/8K53OPIPuqCvduBcAYf5gI/kcSgpi2L+pp
VOz/ofvnVdSujZIYM0f3469l1MycbXLRMCU4CB1LeUUpjipSMrJA6LUwiUiMmhA3
JI3sDJmGX+1JEF+ZePsUFVBbXHx0x6qRNtGuD+K6TuCusIMBq29gYPeceflP85fc
Vh+AzNeTS8vpKWVk59PNlG4NyYmDNTtKsO2fJNkfgfPKOEQixJqSeqgJ8r4+kUZs
7i+rqJpbJoy5f+orjCSSdxkpPiJ/GHQicDjrDTTPDcGhfSfcBiJxxw/uf1cF1SBG
Uzk7l9o8S3hlnNM4EKxEuiptEzyBteVy0TvidIxxxEWqRYJ/r8AFohOH60Z9J3wm
SxsPtGfNiEwhh8AhGwAlGr3AU39Q6P9wxiRgFGXcjqLFV8GJ3CtI62omMeigndH3
iDQyEVSZZSevCWlwMZLLbfypCOCDdBC8TVEjsn17p4bRrPQ53aN3fbl8Q0BsqhPJ
7FwvzusKonOcYWS/GIHLpyebi40agiVdCbaL4y6BNv3GPIfJWxaC0yviMhwcplDL
kgUApy/aBWW7vjVMYLo7GlzgTQt2zK2ZWBS7s67kEy6SU4dkcU4AJSWUuvM2TT7J
0bJn760KAzSfbK1zGDg/bOgcTTFKnHwpszIFle5JN9OGdaU22PfiKJcNhtclV/lD
KpAVd67zy3fqEL1sfMep0fV7ni/Fz4J/yQFCFv98skrpYT/ftVepEatfV987PFOW
P02ziBRuIxSnVKmWdGg8NGWO2njQ+o9uScymzvrOAIuBBFRSW76iiiONE3ZGAewH
W1c0XwN4mAGmwo7aXaAfDXNpAmZTeE3PSarJmp24LAEk/fEYZdHDvJTtbEmVvUPh
DZJmj375RKLH9gxCZNT1U/kPsxMYyNTlvCoMNon8QCWeZWCMxwn+XEcbUpecgsqL
IRaQYaATz7VdKtuWzs/SI22U5sBPKUdUFeORDJEN+qUtuH8JB/l9Xx8r4QS21/89
yaZih/8kkvy4bWhUb5fRcu8W5OGbpjOguqGA+QNBz17CZ7ZuQziSrG78dMRRItxH
mntWmZrQOE111KQenRVP38WrYzdKKOpl+yuHGEr9uRjgBph8y0YbxvdpWnzsfOC/
8kMAiHEx82t/s5cbu2cf9r7ENdUgOcBL/J82E12mseAMyvVzOt9sLziNAtzFq51i
JuGIu0vDZOUcIDlOAL2CC69XVUCFJD+octiNi+8PkBGcNFAsMVQGuPxGT+2V+qnT
5+FGShKWUfVFkEpKtKRgOCQEoEkf92W0QX7pjXBEiD9Ht3SnjaonXmds2uMkOWP0
3qL8Cx8Sr6AbuKPH8Sd+mE/5vn9ww2K13+7p4o9d5Vn1jjiRTMPhTghn/DaUsyJA
+08Fqhoq5MdSQ9+Ut0QZMD84aOxkyxdoIpnDpUttztBmLvxhatj2u6Oc5kqr35WB
39GLlgV7JrhdSdQpZ0yx2wT1Bpqx4N9hKs2eygKLm19HUre6voKT7bHpZgxfMygj
sGzd7naZH+fK8OuGMvYYm6AgOjBXuHdeR7RkLYdrTY6O8iVhWmt7AaC+n1TNFAoA
QH9iVHXnGRirocB66He1PqBH0pgCAGgswbHDZ9SBLNPPaRG7To/XvdkmLEZbDs1m
aoVP+oP80q0GIgAwHY6MJe3Ll94iYEHxEzG3i/zbn+ooVt6mO1e4C8LgEOjo4nFK
DHz48HxPiH/hmG8JdGn3CIHxxXJKG7D4bhyGTRcBME9nx3FS7sf2HFKtKUv5k8ER
CWyOrNlgUjn7/VDd4LtFxPg2NTzetlnJiFSJVPmbz8+t4j3wGveZT/5Sj682U1ZC
n1oinIpNe/0Z7bUBJu5hxk3NJi73J0khQqCvl5QBEYUOxXTIWMNboXMPcP+6EiAQ
3ozniC9kbFryamTixjiSP9NIWngHuTu0lnpE9eSmojSbW1KSa04k6t09q2ZC8s27
7UX59yhnVaGKE12zM2aJP2IAEkcY3+cJPPj5CP3UZj+t7NlQXitdt0k1PgR23hyQ
jeeGHmimZi5PqXIgQ7CYAsp9wz/DeJFXD8jkCP1cZH68MjR+9qJAM1c8smnocSys
v9FKymGY6d8ZbZ2aAapusYLd6e1GakiaZelYF4ruTJmy6lEIIlFt0UcQCM1fBsZS
fVID83LXFj7f+GBhqz8sydEznxDA+6uc6KelXLFY/fNTiSI7mQItAluEZkDBoCRB
g/0aLjpx0bk3s580YIl3T82IOe+hiBDOXURWdEgnJZ3rNcJ7EY0zHjYSsC63Q6AI
SfpBBp1OxS09cGtQLaJOk4eztxUK+oP+dFTQ7mgk5M2BcS/OKyH0SbjhLYb++6b8
7U/+NRu7dQ0eBnfv0QX8eTVhHqIMGo2SP/2wkqt7Qm3Dp8w/6ePNUBJKYWgmY7Z8
ALdQisvMTmVG7OvgTNhTxy6xaz2ADtZerPGDRbL12Kt/rfRohzAHSzXga7U+EzEJ
sjiPnpVXY03o11aTCsiD9rxyIAkHCr7XburI9xRr2Wowh8N2WpKZ10n9anz7O4vz
M1oryGbibIIk0vZJdg+m6t5e+PL7EYx8kiHXPLd8v30pzW/xk1o2pH4Q40FbPPL5
7ZR0aWiUEQ7zZTpAHLSjSXnXCNQ6kOsJBEu9Z2ad5an9ccx+kue27c7ALwDRV0Gx
6BotoFYTR5zML3TVKlfn00QsrChRizUqu4yVp7+9gP6GPXCoZlnSjq65Xm9RGrIJ
7t9HFLykSrVHZzFeBRpwBchAD3M7EzKMZJULRM+NuQiIrOs/lVjeiaueIF9rFGuA
jDh4PIQV42urwLSSMq/v9a5Dhd15CZgGv/hKZt+Lu6yD02/pCZqNTI8wWFjKBtdv
XGATDnfTs3BcgmR/1+wyiLOhUUGxt5x5iS1/+yuNruIVLUChfOnBZdywZV5utdyq
kM/riCsUteNt5hkt/Zb0gA2l/XKrrbalZF2o6LqTq4WeJUgW1I9hb/TOk5vE5fvR
vGmsdlRPblD2xVGwwuq74d7AajAzpv+N9u8aKPWgxoHKMl2ccSxU5TsPcxIOsY+0
X4sf+iFFY6fA6OmKr4i+rVePQFl70up7Ug79Zah4f2mRgPwk5qXWddJYen3S8ScX
5ewIMiB6UaHCHNin0c+VFGUtIHAqJOtuSUoh9PQ3+wyvI6AQbZgG6BoAV9E1TP1m
LMsOAcwDv1+xTx+EgHF+q/NZrnYYz35vGQF0nvFv8tqfmdUHT4u0w+hasxwEl4FM
ON6YS3h7UdBczPu4vxGB5BrG0Np2NCqNyFtAsBs5E89koby8O7Oqp5Psvwi1INPL
u6Vvp9j03oWIHxk2uyYxZqbX25x0q/v1Ol6ryr3J9ol8nBDL/Ui+Qj8Wwm5iU9fQ
lkMupY0zTDaDnUI+pxJM7+Kp08cTcNni86Ws6w2/VZ6op5edyqPboNPYx2Loxxg4
PeFtkC6tqNv64EH2HcTUzg2lAUKQUjhuT79gQ2mvyX5xwkgI5sQYVzQtJpo1se1u
+xAO0bsKtFPqnxC0N6AzjCD4idBmVuWbFYxVEbFzHyoC8zAGMSBNt9eomc2s3Vns
u+vM/OqvxGGjgB6DRYhUD5Zd+V4bDiJowg80Kc5/QDdxgh4Y/Xbfg3tvw5XKxNBv
116ppDFqUUboux3ldNlo1cdTkFFIpO731wKOLho8MdwzXOj+81CFTv9jbW+VX3du
IzfCAmmuX3Zsr4lfRrD08+qWG40yTCxM/iGsdkyAuAfRbDAY7OB1/AOJPrzcQJLp
+Kyp5iTevsn6Sy79N72S/vUJypuTUA8YMPMnfPQZjFib+TdBW13jFliyI5o4PZgt
vjV06IePz8MjdMQnDsustKmKkvGW9hRAsKT5SZNYUfafD+yEKL7CFHDJuDiyTdIo
QvPtJCdIq3rNpHXXwaWuJvPS+Cre3+21hJ/c1rTtdRlcaEMwE56mAqL8JGM/IQdF
Zr7jWvDogmCTGooyrYYj2/2hEGoblApKIDFlr46axKQ3Viny9pt5A0r0FKnWBpjw
MCy8aJQnLowXyXYUwHjhTPIBr+7zogsCaWrV6x1TjoDO4FIWmSASo9WR6clL+3gN
IvZFY2BP3/VH68jGSp9168KmGEYHuYzcExHdw48WVxDHhVM14pJZDd5iyNVX75FE
mxxpRsuIawGf7sLltzF7YWS6LR4fBbbcTAOp78JKqzm6tDLFICAI9sQ0WG25LF3j
0IQHeUW/xCy/ErIezoCHOsZcyaJYq11lEIHG4zDfDTWFfIcxtvLkIfW8XqqWFNu4
mktjIEXdwGFn4wiaZBsVNFyhDZvQsPpCgTHS+O3Z/JLjTzWN2ySr3fw7io8yaUuO
m7qo35TUNHPUuAOEzYOQxYJYA1NXkGPntzzh6OO7bF4ZwfNGR4cp0V9Z5ZzLLwYL
sjchRfU2myzX3uFWC3oB282A1G2z4fLen3lzVLFpu4lRZERJrRxvBA92fUN1wMYz
yLZoQqb2pGXML+08aATxibj4rncv7PIBujcjyIP7jlLs2bZSo4IXfeUBmM5TCbFr
3aiDODlwdoySEaFWfyCxgC1ObeZCvdKqQkrxKsIrgQZ5fH4UL8BnTjp6ePM6uQqw
jb7Ow2MmhneggfzwxtQG3l/YMYt/pNSfqYeXzBY7SIeCi32jRAJUpeenP4hZPR3k
yuDDHdjiHo7vRxQBBY5DtUWnu3L7jVSuDPe4KccvsZFzk1B5hX4b3JicIcas0+8j
lyjLPsVsFWqYX99gDAy9mXaM1Z4iaqUNw/YX+yLPfE6pReNokXfsD0SVKRxWdp0N
5B2qdfWMoMcdrzw5drYKdAwZCyzIcEZd1O1nulss+HEJ7zdd5Pol6/ZHmsqn+/9X
MwwA0pbEV6qwJPIT96MmneakvzsYQQv77HIo3m+OpOjWWMacGqYN/S/fYYO25Dmm
t45AEsQjb/UEmUTSOGx8jCP1Ao57HwU7E/aHphmBfDlvnzj4lsveZZL5V/19OGW2
klKwaf1/neilIZN7c3M5y+Ius6CyVL09Dt0pE6zCwSDz/ecSOT7DYhMtn4fmZRrw
ftMGQ86l6wq0jvm56pNa9NjBOmzrXs8cScBd87x8YpEMLzfp7YXROFnqnyBkfHv0
v3xgIxSrgmU6t169ttRxM/qhWoNjwsBTm+WOypDcMPEfNX8Kteim2bXNFsh1f6Pd
l1CQdEIUyHVgeog+nTI2n0TZzpZN4R/LF8gcI1GsJS98uq9CfqRbi7D4j8r01Xzu
QUWAIQwZC2cHYy7uX80tHaYYzVub0EetH+vEuK976TNoSiW23PNyNceYiqNbykhN
oWkpeZnb6c8TtoOIyeMPTNrYB7up8APhHlfd6KIzjvFQfA9S/BAo8KV4sA3l/yvA
ztu10teXI0gu6wqgGEZtK4xBivF723rZN4aEtWMchWU9VjzzKUlpJPcwG3ibwI6a
ymZSrNB9hNNexCe9ALHAcqRrKXYrFr4xsRsOSapk7FaCh23XRCk8Z1UoBmtRnaeE
9S39hWKHOBmBzUxKvWDB627x8Kk49fyjHnM7nfOSd3DFWc+iJv7Rsou0Nz6VRmpa
/dSCrS2ZnCh9JudIngwIqpCgmHfE+P7chPMcQpdAbqKj0gpYF+c53Ji5hogOOQJE
UUZLrr9p1id14e/MJ+LePWXzBpWJrsOBItUsSNsUkZU6RnC18h7nBPi96mGWgXMd
xcpqNFnNlo0zhYFEUyrkweeFOAnP889Y/VdqO4NLwLScgm51q5nRaW2hccrdzA6b
mOQAtgEDY0TcHkwSH96W+FJBr5VQ372koX3dPt1sIv8u7I/5yY/DVrTZVXOAkuIB
zOOp0Sp7d3NLOH3hczxn0b/iSktPtuvEMuaLD9qIaFSiXz0Pst9SkL6xIExm1FC2
lLO9h5qQpnrPGMZ2mbc4P0xO/OsJNtUuQyuhPOXVA2UJUW9dDnWx7fLyboVuU4Ut
y0AT4MFAO5v0foFFb19dxFOr4ecrFNVwcFqCd6p0RuHE1CM7Sfuw87iT7D9rIZpU
qAZEVf8saIful1/2EG8xhKPJfJHITRVWGQZYHR/KNvt9XL51vIfeutKJ8rzfTGa7
6idgCluxcsrXEr+SFJWFHGcFaoMSb5NetLIiCu9qRrDUVz1LYTBuOwksrdZ2EIGv
FKOr/ESaMIPjEjYwM8MRem29hzQTys0QxhOiYzAYMH55W3KT9z3e7mX0mdDi1Gma
MkHz4Iej+MYkvdgUVt26ndh44pQoynUMCywgzvhQAHKmD1QkZdD+QB0P1uah1y7r
Ne30kh9XMdD4yWI5R3zPNf2dHsP0c1kO3AGLhqQFK94OL8wCf1iry4U02vMS9b1p
V/x3UEsUhMfZlhadxWMfHpBxfS1Isrw/lVQGvGrW73BM6opuNWXIC02ky1Z/Y0vy
v5lDCDnG02qhZuQ8ENBTAVOfJyIvEbcl9gOOt7QIqBJgvDhM+Zp7lVKtn1n1rLmm
sKrpMevyDQPydFbFGvIV3A6af1kNyWFhtGAfPrILT2b91gBnVXEtsqhLBCRykmGo
Qkuro4AFLMw3WTkkuxUhGTzkJ1ZeVXjZqxB/IGLPTbvNLkTWHCLAK4lGFQ56SFyu
v8vGcelpoImn8B1KATqG7wxwYG7/yYehzn1DxIZt2BMgEyoaiD77d1SGEFBVcNZg
EfxmZtrdNrVFJxO+bmw0jFZAiPO2ZLFPGvrQYVVcPV2bGzTcAFVPPCdAvQ2HcdXF
s6aoNb7uKjfjQSDJ91ASoFrokznf6wK/oDJ0usW2tj++v355xYUI+SwKYmMoLo0Y
z5Tc8tj3Tml6zMLrngBdNFivaNgwqSgluYRUpC4eijNi1LP+03Vkiqy2N5WeMG5K
EomCizIUzFsEH3fWYp09zIicRFfnGoHInOfB7Wau+/Xa76kQksxYr1C/ianPqgv+
k010wPJP5PVrKoysuU8xiMeVY8qopCn8n7/9pMVyamCr2j01mFWMfzrzNX3wCNEl
cx6mxHb/NynfLWawsxxZo0dlEf7TjRblRlxzByYsb43eAhIrSPbq5hksFagnP5Em
iC3DlcLt/y9B35DmsWtB47/89vGyfrVfSSy7Dp3oURUpRcqU/VzDoEF1w9EZeSb7
5u893FCbIaUsVtLBGNFEP5ZP81KGI7HLnY10V634xc3p9jTbgdKWXdtRCzf4w+GZ
82qG6Mz44JZk+nS+WDhAvSCjEwhKoDJkFtsXpoTyHvrFl//hfjj/bNO1wBmGlkhF
mDbX24+x4ehDre1vje6hk+x6nFMf4+IyG5mB5nxgGa8zpNbkDJPlotYesWe6+B4P
Z6nISkRwztid3862ESJX70ERiJqJ8a06w8t2bk50VDCLTh+sOhnBJpFdznTmMSpV
eAJDvfC2QnZIHzkGgqlSR4VhaiwdAbEeoDLCMklCeHEWDIGALNUhG2MPySjJDAGl
Ya88oTEYKlWkT2icSM3M3Yl0lcOuL/21Mr22gBVtVu9O7P7dgqNmz+jRQPt8l/m8
CIFrAwokEy2+dST3NNuXa91OcDb06f3lbbPXUlidpc8Mx1ZMQ7/XjAEOtcDslkX6
Gp849/hE+LHvQB37Hg7FbKQlMVfOePq+Fohe+Sc1oDlCBRAzpzemPIzQw/9k3cXY
mkywRveLrkZmi3eNs+m7jhxZksltxH8XuhpYd6WreNRlqwRTRhl0uojLRCs/fX1c
D+ZFDKBO/QOvlRAQ8FDjyti/EeuBQES8kseI6dZmi5nWyqia3MtKmoFywFLKEAXA
VuuP7kd/LMRN9QMWjiUcBl55gZrE/T62X5RkCTGUFnMepHLFY4Q/k/e2gwTX4xuC
I7j7c/YxeSwEyOsGq9PwJa5irgXnTUXMreJKbnFVh8qa82h0ZAjgGqE+APfBH65a
A4r6MCucQg2jBTY5e5ccQrx7jQQfLUq4RI3LSsPnGRiMEGQ3fAOcBfSwFOTiwzVE
N3nM1Ao9FU3lG9oPvlYrteykcKNmGWn1g0420ZY58KLhbzyCiOx0PESsDrScXAdH
dAiWudL2kyW+QTkH+krV6E8bVbx0gG+63mTx2COX1fkehG4XRJBh3+2Uo6Z/sDz+
jHtq8+KJYJbKhflZ49k0jc3pE37TS6gLkxLDtkO9pxw+BkRCIBHS5GRbZjoWvA7T
jCqRv4plolQyjKOWuAG5Zs8YvS8E4vX3UiNRPu8IvvV+OjlQbxkc0lpLC27SgrYT
hyGvNfeE1IA8KhCyZopZoYbplXhdw5o2tC5pMQNluyBk1O+72/Akc2jQLChPEHA5
m+vAHdqnz3qTTrAKwDvEzKrxnG6/0kOYyxg/q7Sv9LAzFEsS6XxwFzerkcavE/bJ
0/ZzYnjEwl6tFqJQUxb4JBtoQgiMzS504fd4qeVWlXBcFj3MSqdy6KBQ6AKBqryr
jHtNde5IdP75QkLZ670Pkj8MZzIZvuy7CIk+RAxgKU98vyzAJa0gHDJLYWyoJhsg
M/wN7Pg98SaSBnh+SKqt/fJGg6JK1GtOJwGN3ZpYcZENnp2lCu7uf7kV3RXavnVe
JPlwhjpz0gEDmsUFR5z6Q7NMD+x/CEKdi6Nak8O/WswTm62/weSgCnNsuTAZW5WS
i2+R1HFn59UBNZJdZSRO7oEEaoreWDIZ5spwcZMFOOlQb4XcnMAoTCtDny+JYSqw
QfKoes2xj7QMy6Ez9xURUD+ugdgSM22X3p8PTlNlF58Y4QDHkzQ9HbfUNA8GzX+i
k10k2fxA5xddH3MJYEPBD3ixA+50eA+iOMHBzc+JQBqjz1rf/TIWBfA6aa8iOr6P
/WIzZj1jH4FwuBrTWehHyrfEzlnadnwf5O5bmx2aQyCR/KMJ6b9jAM9XORcmfKS3
p+vzLoeKutU5U/sGtdgMlzb7zedzI2+1KRr5Q7ZEh+XYszXr9Jr1EBOx8aFjP1m+
lDJATqFbLPNOa2btA9/aF7C9meEnZr+XoICRt1RgBZLfXSC9L59ruu2XENlH04s3
wJtrTJYiV1gfs7TkSk7GIvVn0QvCQYEvg06nWBwoVOHwVsufxIqXIpAR70LEbDne
g7znjGIG3aDB4K7dzP/ob401JNDll1GCd1/vt3CTjCW5TOWVg24wbugxc7M3qCvN
LljNvx1B9NiJ+0ZjaKV+WkdubJpvUcR34xcX8Mzv6BAzZ7xbmZUlfeBTaiKsC+CQ
14zAlNOYPbJOmB+995JuJNvevq5v5GCtV/kx8np5afNRCYcVaYGXEDDtFKW9P6T3
hsyxgG/isq1qbOOxOB4fsYWjf5V3klkubfNZVDaWMsXor1FFoFWdlQB1aXcgdoBd
3JqTYnqqceERDvqe2ex13ljCZoC1cjNNlRQvyH3aLhVSydTKci/Hntf/ttjP7DMD
NpEmHpEUftP7aoLv8VhTNwM3+RjFKNd93cn7bTr+3yC7DdFvjf28HSTtv+eshk/x
5u0XKrnykTgQR2Uzm5B7+1d9SAK0zuUY98encHWb3PYkmgOjEjcUWIIk4pjklxTr
wEIgHp3nqmhkNsIdBJH53/NynM0wvTrfKuchghqVIR2Pu3bw47L/z3mRZv3xDc/O
k7cXqSXdp4w1xP/32+dC3zvsB7FJRp/5t1v8+38SGy5zUhT+t5PmDnQW78dWudP/
SDApG5oLbK+eolFNkKFXqhmtpoKKXCC9taGwh6Fht2LV32xRNn61JLz0SCgRqRvi
Qk36itgbXXqW1t8RXuJ1a7vYIdZGbR76LTowB20OSxJBIKR6C5Onnh1CIzPEX3in
/nEHE5ozFfmoklkUZtHWq876E0kvQeweggo2yo51TWCucooiqWJhT2hjTtdk1ddb
/9X7a3otkOsbUUnvzVDovJv3BHo8E7TkzcUe0PpjpJ6QNMMdLa+H8Rq+1wPU31gE
LJUV6x+GOWFwGRy78p9VVp5Wfqg6cV30ZDdlQN4mU8nDorNFLLwqTw+dyKt6ApQD
bKLpbGCpY51wPtlMebjsekf+WU5/p3v4lfjGvbz7ckwT33vWqNZIMUtYz98K4FFn
mH43wOgroIiOo0X9b+uI1hyHSU666TAmeXKj2jRmicpKRtcLSb6jEzg/4fyiyfLd
lr+T+mVxarGRrYyCpKcqaX9mSS0JdP3jtEbj+z+kxaX723ouzlVtwrexyP//9Pj2
+uHSTqJ4J2KNicw6QWOniFTc6CzAfluaW+R5HC0MEZGPjDt6XTXDRAd66zQ+k85Q
7o6Nq8AUG+aBhDH9x1q6xz6F7N88H7xGRQE2f86uoU80po54P5Z3jZmec6iWg5Ab
aPuGm4fwb6gIzJOdiZTd12777A3QKuJIyxnFOcYln/Z2basRJiI9tXVLG8ngjNCd
o/YWftEpAmAPqPu2gll9VCGWggbNIbUP1jfeheMh2mUmQUxY9aHIbVBOWWyRf+ZS
jgdWOJp96JeU/VxdXxOS8w2xjH4OU428tka2q70mbn6QmbzZVaAlE3EelaPhppBG
TM706LmbgXUxxSlWSMOlUf0KOxRfi5tbHwWuPZZwJPHtcuDtbC52qoaMVETZhq48
8XVpZ4GtBZl+wCwz/2cyy4RUUM0/azlnugjDrOCAeFL0hz+nvIfX4KlnvQZYlA3w
O+p+xRK4TNJ3/Y9UXnDAPq+yEVBAMctd+mQ+b1NsjmHIWU4msnvao/GoGIEIxcwm
tqFpLa4wPcG/qbfEVk6M3DCPuNIUgUaaVMzSr/A8xQ084dG1XWIzjAuzMBy11pyv
y6RyIpheZ0azr6JdmQmnO4mBkgpadbiCSXfmUM7dNIGrbRbbHZYc+k14QHM8Z04K
269u0TK2VN8KY3w15Pk/iF4n3QQZddUWmgiJ3olELEE2vxCdaA4maCRVe3rlb6lk
72BaZKNeJyLIX3MBT+sPSLwuKGeEyKNKOI7lyx8fhq8BQ/D/zFnlCPR4Z/eok7Yu
nBj9+ur4bQ1QPFEPSk0n9Hff8Xpc63j71bfUKq4REe/x/i/SJnqJCMSzexVEaSP+
ouZTDElGqPTk+CLkbhBnkaNOudVHqFb1un0x3Hrxn0els+rnh1WnA0YWo1ic2tfU
efykVc2vVTRkuHxNfWRK39N8LlIbsDx+csA5yBtWb1KVAMSQ70fKGOXSxNOgej1l
v90Gd1QcjKvCImgVf7fD3GjJiWjq51YgiY5qPMb0jL1a5/liEFXj3fU3e3ykq8k3
QtsSz+3FRT0RBlD3q+XtKUSqVvUQOoXqB1Z2/CiJVAViHPpIkeq1Lxc3mOm+gY4q
d5oQUztgsV+1haSPh7pa7wWWXtyuzMm4WnNyecwGfCFGd7VDwcKs5l31GRw4nJ/j
71vfJkwhIN4+w6cLvZw5vZjF+al48s4w9WYztnmBrCNQOk80RGv840u7EyYbXB5e
K14dTGqDzyBUa/aAeW1m+psfw2wHnE7ZD1CYO8B+pSlb89z6BiuqYTm+HEb3/MJ0
rsXPucEkoDvqihbQxN2SNvkcm3LTdGCwfVYtdirjlfJfAUTqzxUqMQos0CGprV70
2lTQcpNyJ+4I3p8dyMmZClcVwYBFBmOrIfRwkh/vMQljAs/25E8N/QLwOKN74qUv
oFuOm/8ayYYdvVe3bwWK7WD+aBN6xtxp4mWpfUJ1Y+0hI0sIn8bN2KpWi8RnRlrW
fYqiW4/di3MV61rBmxdTrNl/PxM4tqR6O4qQI5CBcWnG7S38aF+qcIfdF4AohvV9
5BRHoItG2IM4ZlZzA6mBJET2HnHBlgHLy7BWpi7pQ1HgCWTPKpFpne6G0gXj727h
xGHy8Gdy/FsU8JX2Ymz8QD6j57juFOD3QLZnyzZ5wMjiWQytQMN12JxiAkq4Xhht
TXyA7ixo6iLpi2mKm9Ai+J6bQUOY6n7bHazJkRsL5mQ7Y1287HmATItXrFuXOc6W
g+3eTrS/13Y/nSNwLLcKr5+QHlK1aApPPND5/RRMBnF86uZzMHWglz5365YHFLA2
q7DD15SuzEdnEsUw+ZNUH7KDHUarFRt04dRKiJktt5GlbXWwtzzA/jPVwTPFIFfI
9gBiet/u8ea9RLGT0en8rjdP+hxji61urUAf4SK9Pc43j/ajWj01WJsneRl5844j
D4/JPWUNHxZTFuTxOCExcy10nFiMSDDHcuCmUvSeAh5fYAp192jARbbJLZ05E23Z
25bj1FOHuKL2NN6shX2RD9XupwhSZdKIOHItEAY28X75R9/VFNmmlROnP2K13bGx
5d9ujv+OHBArqHMjY5PRLV4vYt3ZoQJWcd+GhUkpJLZ+SBqzeUSeX/6qD9MYBvXD
clsWtgOZ78YMju957w077pRQZyCArTznsXMPZsAmDpN1MkxMwwPZ9JUNQHXB3Lks
VG91xUtSYYs3bfxxOIwTOvIkzW2ckLonszCAFyIhOIZq40VFWD+xICabmiHJ/M9f
3M6sAO7llgUhca9/kIfIOzKAMuHg/F7PMN5vANrCIx+YrIGlNqOdVic20Kwu4FL+
p2xzpdAy3aujzTHriR6rwN4FFIuZly0ArK0GTMz0ZdW63Xx43pEQfBmHjWLgNtJM
e5CSsamTe93GLBjIDBX8KGmdueJE5Fde3DB/7iY6BWlnt38iTpApfUmtOLK3MpaY
rq7nSgfRTwlze4hFjRiqBLv9VHNV3TyzQJ1IUbDpHbyedEr00WHRrzyy6jlOCgyZ
dKVpjE7ug4uk/aAksR+V7UPRzqd7cn/lv+dG+zALQ4uRJodTirYIhTSWmfjJ4RM5
0xyYIAQSTAYG4yYSPrzduylVU7465tYhsjyPmahkXPwE42RgcTJeREbs8QIGQvbv
Y7QPfPdsw6b/VjX9wug6x161+/WFDfJD9JND3hHibVokwlsCBHboMXSRjJ5KAi+t
9BBIK68/ANAKXPGhWaGVnqDrR0mxR5xw1X3I+eMEJeWxxQfs6TxLytxBDnZci3c2
QGu0ernTbHx0O+FcB1W3JIGMQsYOk7jM/af+PLA0s3vNvt+v4dLOBPpNFMVC4qVF
YYpORAukzybxWlnmguEZwQW88T1pWX7NkYnL3NE/2CxHOFMkJ5pEZVSO6gOgof94
dXyco129lvpAgYjGklk+OJJFuDSM2Klx6mbbvN30onwaEJFtRvLTGo6KayMWnTrM
ThCmqyXuBVTE7khj3xrqw6sCp6Swd/Peskt+5THiXNwB5wRxD+eo0cKDue6gqk4M
dLJyobfFbhTXisKoLVfal3QrkZvc9rM1XsfBUv79/xu3edAYgsQ5COdjL9ycfWpI
MoVWlRJMv0T5zQFZvMp1ry/7nUPifKQbXnEbFV2ypZRuiN6SjcgTYJKOKn4U33tO
Ju5o/89aLHy6jOXApZTDJg4oAIGkD9kDVJK8wXp37P142Hzl87DBDq5U4WS3te/U
3hNyg8X4lsdQtXrDx3P98x2YLyt2vXB5WCjX0zgFavxQPEUutErEMlle5FRB+yNv
jYO8/ZiUeihAav0dJBYhhC99owG9k6zWJzj2r4CldDfXzcUxiUeekiAy0f2DO/bS
0rwLEtlzL8aPl49ePZrF0INH3s+rJkGb0zb6ppVN4wq1ZV2+QmS/dXG8uUgM+1B6
97iPtoOMH+7X1LIg+fbeZRFAiAur+flUFqiatY7bHY8JVAHjN4mHxvJXCL9k+4Jl
Yoi9ItlYBA2VImiEi7GrbVMuUZpuvb9acgMelYBka19gAdP0LDdZAkBk5CswlbH4
13MVeckpH5n/aI12KJ6+lWOAEurb0KdRU04zZ6VWa0NfEAla8s0m5ebLhcsZGMwq
XO8uCxjPKL7B105BtryrlagtePCBBctskFmoQNgr73gAczsBuNbQkGOPx/m4kMAs
kpfF1ZB8woEosv5+IUt9GS9AaK9mkeXl0yZN1Un1vZRtjPihTfYNmOqzC2qpEfFg
A+7CXecfxBDN8RKLW/C9OpMhGHHT+fUyg0K9PqDemTs01EUbGyjIu4ndFdMzd3Hv
1nugyNWcDg9VllGFaoGO69QG5nLsb7atYDQl71hhvmi/A/PyCK25NYzRkpTibEAg
wYkGADL2KIULs61RSAkFoX4Q5DK/5bA5uL2+HQO0aUe5xFYMbF2MwzbOI4Q2UUTL
AJR0UMSRkIEhHN8XcQls+2sdXTxlXbtkoPrlzkaSf18Tw7xLlEBBdkXFt6IDpAtc
pjeLLP4A70tA5AkPsJiZnyWD+S0Sgdh1ut5TF3Czj/dSIcDZul0L6pS5f/LH3Dpi
i/jlQYVjR+2r0mJlbbV2XBgMjiq4qg7fBLy3fpBrfPMdpOQ1JsH8bn2acY/T/iCH
IflXtY45QVwwwc18chC1W4fuSrJuLcUO3bw0Fepw3IpalWvxTKVb/iNJIyQOn+5r
AfTU3Sq80VXQdNJFeiGpdZWdwddPF4wzNc3ChT8KBRO74ILaFYxj7dZGfifbDCRj
TMAwRO/5pkdpbwgjqSqaxGC2THdUQjFVdjjHlo4c+Q9Oe7c96LMkiYtaNMNYqAJ3
aBcrgmjfwxOxC8ZDw5VMEOhO0XGNopnfjy9K0MM9cqGg1zQjMMLQrsgRZsRKD5V7
iRB+LWW6tHLz/HfWLmr+MUwzRN1A+lt/pK+O1i5BSP9TTqUSxP+UOy9VzlCkJCNn
m15B8LDCBHFwGG0qyqhtzyoNrXyDaLVY72HJTvdL3gbvhvxfvkNnMChqrAAlAztb
s0MPf7mIE2t+cMkwUuIpJomHbUgK+UWcDEJk4YuI8mavtfoSlOc458N+EX+qQnVy
/0V+ythXskQiurYYlrTQTcV8jL0/dL9ZUAjGYH4aYO0jm59J9n5GcpaCn6guFOA3
JhnnHhost96/gkes/Gf/8c8aNU5ZROh1IxVmIhqfcjrv3gn/hT2UKm+iYblzVa1d
pYVhXxhG5x8NxiIQRdORqWcZO3vpZ0cjUTZMVoZQEyfa15qlhsE4yNDhsWRXcsB4
uOvEs3ePCZzq47WlLFs08Mcd8RzsEOM9J1HUwSx0wyHjpHKhMgCWDWHSgWusmsXS
Bvo8P+s+cf5qyAjekeWZLI0zjLjqD4aIO+5H3OLcXKYphlxCl8gHvaPAlmoyBshv
+Mv9pjtHpekm7zixRwxGLtHL4a5h9wN180NH8xVX4MI9xuxCt0SA4on4bykZtEkx
xBhrvrhyEvKgp9cplY4vkZdOkW9f6UBmyUh5EZ4ANTc4HaDSnU4XqnnYD00Ck5jc
IipkHGwVzEYdq0ixbq0y8WVeK+oNT8JiLC/BIYNuH7BH7GURt4wp1bIhwid0KPDd
NmEAX0qk6lJ08a8MOcNQagWzMMe9z+xGxL80jvvibn+UgArJjzp87O+xiTeT2G/w
91gAI5jrVwy7P6/x2iSCCCQ7tJz6kv23R+XnlqJD5GplsnRBVR6ObwnKsVUGPh+4
4PYP6MBxQrAQPKgc3cvopPEk8h9I5jWihz9ek5dClBM1AN9x6S0QlrzKI+g+SCBx
wZoxh8IIn2UEcuveol6sHh4hnUhwkCsRxBy2nr/Iz3y+EmduydPa40NE2BTEO1ZS
ZCDJryGLWxHBbaPm4znkadTs49h6LCvBw51dQmhZ9DhAUe0AN3Hx6LEAQKh2imYL
itKK5znsrsXKOmfLYpMlgjakB2XjaSE2UGGU2O1gzjogHcLvNqoCHevDuadjf6y1
9x29brD9Z5RYg64i0tZvE1/yLiSwEKBvROrJ6KWbJhABCEauWCqFjr0DbtclzqW2
1GvHQGGnmu+PE1VRHFgSiFgTbIyM9j6w3jmjVzGzMLtDh242ixTDlavaWRpTixoL
cnkhFzY9Ruvy2bXmv4EEGHIeK+b5zwPDKDFkK+EDWo9a/3+s+2rzAiCIJz5PNgft
UYdHHxWrhYKPdwWhfJaAy71HkVQnPkcL0l+HpTHxRPi/EAY+Lgk57XHijp27sFJY
M3V1BOF/EQkYFjVu1V2dDyRNcm75kiFnr6d02QIW5wlJL3x0anW8nYbI6DzS7Gwo
d7U7oHoew1+gnuKjg+H25vgnLXI2TK8s4s8jEbAf+2L+Vf2qXCjvcYfYPTerFlzf
nxzatXcGQBfxb205rDLnHidJyhmuk+KciqSeKPKIbLna6FAYqqwE0/jIkG9m5OP5
NtKhZKZN97Gu0sWrLGZwPO+vdqrpjt7JcgmHJeZH4SmFv0vRa1ynmR8Btu7FYcYV
JxHJ/0TvA/hAlnHuCAgh1wJffFhLI0ZjK6LJnCYZEK1/mdgmodltTlPxzRQx7w3d
7e3BGnUhy9o7h9oOv+sY0CGOPgNfnbJ1i++jvI1kJR3TJ4UnQV6oLk0oVGrcFnnO
uf8gikvhd0t8fkVGUdjdSWLV+mbJot2FlX+2jaYRoynEB+C7x6A3vRgoXYmSRF2e
CAIZ4b5ZuNxPeo7+z/9TptSsRutmMNPUN+3eJRdw3SfmttsYdCE0YNrGZYG8bl2y
wDLQ8OFZGPKbi4asdFmTnJL7w+0Ic8CY9HS3If9UEFdrfFdcrratbXcCjdQpawCj
9qTH4NEwqoFzHu8P4SQmCutLjjKQds7wwHmktOxWjgXMm33UZIEruiPm7ommkopW
Ap0NCBd9fWJBGbP3+1CDnw+MI+76wH22MiBNyLoQuOAh0uY6usUkdT68si3fJZdx
YP8PDkvT20CM9IEcFUQ7v2lr47xK3f4ucBRPqP7/g5fFZAxxok6DFNCQP4aHQmNU
VxdTtcw34X96Ym/LTpAeYLeVSCQB7wo6ZHJptiTU9tg3S0/JMmj4z+lfTZNbQCkB
Sy7mYvuM3eMxR4WkQ5j1EuS8ZEKNSJH6DbUbl12TJDHxTCUx1g19Vgjltr/guDmS
6Wl90TLkglnaGRmPiqDJSkNZyUjR2ohuQLNQkKvbfzHu3dWVDvXgXyekJy5zQEDn
B0n8pnnOa7PypuoZ4NFsfTFOIY0EL7bCK+eqEvM6g5xSvXF1J2UvVwdLibjSFEJ7
523ON38MQM5h7j6aM5WbS2em/9kLqcd9sHhFc1NAPlOwA5kDE9AySR5BQlYb0kKr
MimsW77zThFMLKHSRe0Zj1vVyjvhOajBAJSL75k5Bld+PYt0o9weCGZeAeBuPbEh
EPA47nVfe38VlbNXLS8eb5tmqV6N/VtdN0TzM5jKdKJFvxcOks1i5IER1TZvpUKX
xeyiPdveCDc+GGaeV/1vU5trlHYKEFyKeHmetgyznhji1KbBSinTvUS2t1HuvFj+
fvjsKLR6N5SuTMcbmrPpMppi5TlD+z+q1odLeivSAeQTl3gf80AhK0qiI8wa3z64
JKzc3txjL8p4zqaW/EvOq0hbYSYPJNHRN4Yuz4+szfRtDsdFmZFZSVMTaAtEOENg
ySSIhM1G/fVHz8qEyxJR2PkVFjrfUx9W2R2Sl6DAmp4leoaBEaUKCjNP7Tpj5Ei8
yUCBw1qYf1xj94+t1zB2OxsyMWlcpocJ38KrX3GETOPHMwOObtMreKKLZsEeWH//
yj3cJagrXerQCs3cKQMfAnyCJQVpHc8gkxkEkKYyWRpoIgXHcyVP4mIU8rR1mAQi
hHB+3AU3+q5Dku1SJI9wBdqE0xRbLEX2MV1CZzjbiaMtP69nvULj3NkGwfnUtDNW
S4r7IPW6jOKLZOqJHYWMdcfYAUmim1jfgUnaizqELyilcNvnhs7g2zTX8vMmg0TD
Yhcd62LxzYFb1uFOOW7b/Ib7uS78ccAitKsw+TB4MbqoVzuhWXqAW2WW1l3fD8UZ
ojE1QhYWjyMPQ56v+s0JsC4nVoBQYSM7DQ7/P25Bihpd7vu2kvWDSnwksx+U4n78
1O6ObK3y/W+/4jnJofQ9UTqjv6298ZwcNmudEIm3HyNJ/ACC1RhByjDQLWyO6pdb
i6v5+KINMPPuo8j2PK/klcJw4q05Ol0dOAZg8+PSl9XT3feDOxq2LloCuanzmsUw
eVRabdlUn9pNKLEBUSzBRByhuSGURTUUg64HoA+RHAuZgGMokNX9wjVWvIKef1f1
uxUjpMCOPsaFVGuzquJq6GysigBXJd3qBfHWUWoIkLO3ZWUFdCU574Uuo0L82Quz
Hs+R2qBGT3yQPooGGF1ZawxXMIqAKO35YaVjJBHgFFgPfBTXcZ35zrZYcOIAtzR/
cca33fRFFjJGP26fZBz30WyGyxru9He+bRfebprL8EGgLQoq8/1vrq6Sxtxm3uY9
7MkAfnX7nkKKbeThwRvG4M6RTtaF6hHn0oCooAs44a/JFW0zhOSv7JVRBkdQukgn
ztPt1Qc0B8885sR2/YSN+C2mUi9bsBGrWCNNpl7M3Q87Z8TH3fKNH7eY7kwhA+Wc
rPfY4Azsv824lmqEDwtu3GmHyWAF04DCXU5OzFbub1PjPjbqKr/eNpII7IX0S+Hj
No9qdU2/r7zc7LErQbG+oZwPRQHKpVGS3qL0wZbyFpMVRyx7jB2Mz0knXgSxYW2T
iOlfasQhhrAQuu/SP+KhxkC3W0/opMk1EiuenbYE8nuJ8H/Y6hYt3uMf18urH8v9
g6t7CYh7277C3JejecQWXvKaiPeG6R5f6jlyTkZap4Ft4G+/uEPCya7G7hvMUmsU
+cnXx6HZGbhPBskJ/knalhIjxMV3j5EMLvXkZmHsHFXKtiMK/EtYEh19EhYPd8Im
OzeD0t4FzmBGS8z4grWsYXieWIornFwj5ovt53YqIAAWmwiddFxskAixuK89dh5V
9YcHlLRR1hX+ZC+eOZreqdGvVL+sBlrpmTbEKTAQwar/7V7Y/M2XlDNqTnvlUVTE
NhUYxKV37I/QCUDfYsH4i3UH1M1pNr7FmPTg2tZ2cM0jj0spdfqZTl5kzQxUAhBW
a+FaDqjZiy/p2Kk3IG6JxNagKIrHCS5B5IlcbsabUxnAS69rS7olSH16ndqIOVZK
Xr50MWd0Jz8LZhG+BcihJrGkyoTUdq+r3uW4Q6OmlJGSsHnO4C1mFRbu75xL6VH9
H44Uf5b4FfoLtujeg9gweKyjGIxRoeJc4YOQ+vZAsB/ESEf4oogjxxezUP9nPLQM
5jSIVhfCpI4MnDyNszydpDb6O70/eK+Z94oJMkvn/qth9PRS/XDTOq/KH9GzKLKS
rhq6dkftnWnAvhTw3Sd2i11xLj8YiKNX2E2GHeDY4+og4mGCtmSoOEt/nBRDSUii
TXxu0oypyl5KU3cXTVoB4r4ivxbRNIpAEVTqTkIQZzv1NgHMGxLMXn6W7TUjS/6S
+prmhTl12AO3QlGTBFDyT6Q8kcyfor3svJvpSZsb+slI5jtJlszOII0xXQNwdHlk
gGV+lVhKhfutUdZT0m2hfjq959nkkiz+ap5j+kqiZkZMk+a5UgqFcqHFWYko4DhF
GQACkMNuWC2PZEUYd8eK6csEJK8nxEwo0KVs1QofROr+Qugali0cTxI9tEl1Du+R
NPgzeZ4WPyrJPd2SuEvyM3uJWyiq6XPaPXFBb8UuBzqiWBYvkNl3RJIvDC+el4dG
nB/hj8pvYEKSA8o+wt8uyjxSSICl7hCwKajTTxzaOG0gSIRdiy7EFjCC9DbQlQbi
TJJnbdWJJnd5j9rZBQghrPeHv49SagSpY0wVqybDwpQTgfBrWcVxDlsIjEr2lLsi
c+w/IUF0JfIi0SqO5lwYtWaHlojKeGnEI1IGMINZ2OH7pRkc5nzHud9uz8ZIVCHZ
KEcWw1wfL5SJ1lFUA95bxpjbLoGG9YTMMOezDwVZ9sEgLKjdeBs8H07INIG0RimT
Utk3f8VUw3aTAQIrXREIyIUP2IAS+sHJiTd3UbH28yppEiMMlMSVCQyhdh2XHrrO
TDVFjIRIor3XolapFonNuhmNQnj8hBG2bgvj8vPw7zDocYMyZoiPNF0pVVPFuZCQ
o6WGgh4GuE3cVLfHGCCvG/V3JG+qri4hB7TC8xsEIJj4RtgMXE1N+HRBJxnXHtDP
31+e424QH8XoVwqmul1wabF8MKq4bV+fpss4aj6I791/E7b+Eqjf6gM3Onhgm8/E
WkdjaMnkHy3wcT9stzOD1Bi/T9k+HhYUtOq6c8QnFK7H7DI4s8ywyQ3TtxoeM/t3
WRdvmnTm237/m2j9BHvvpYvYbxnfmSwyLG19RZ0IIKm7rMBVJbMXzHZk82rsdZ6M
DX92zsd1Bz68GK/bMfoqhGLVxfDTbrBCIYGgZ9TkNB0OTHFFTdwcVhS63YDQoUiv
elfEY0zUdAOYBUtNdmZ7tympt26/E+xn3tZRzblCdMm6BQB+svYi/whfqXKNKeD5
Ya8N2jUQTBmg7pQESCdLx0b+feXrJibbB30UEE30EykZSDC7wRXPBHDySLaGSule
7qdZSUK4+lLDQHdpN9vawRXY7Sro7dAWieuzqYrIJDVMFkf0QB7byx70iJPyICgr
yJJGLu+F8cY6X+pqmew0+eMvqDc3OPSFhn/JxNsi+4SMud+olGGrSk4fWLISEx9e
M4OOfUrFIJTjXSxEc8exAp06uNvG1BZZb5qPjW+2cjG2ZnVDI2tvj1lwb6yq9j3e
iAOEiHnLhFneilplyhxm4hV3aQpO3/uG1Gn/qVS1TGXfUj9NSr+/okhLJsA00J7z
XiCpkzVSmZx3TxYHe6olSdHrVaxAnQCTVs0yeeF0GScPllUuRtrdcwmne2wwX8dw
w2wL/iLaa+glsaeSq9m3MGUiIEMlBQzUImY4H+QZmIVoLS9lRRCcxHTY2WIFUd61
noIyVM1dCmIXyK4tJSt2fxuiPeo/zypXESosMlgYlxBYkpKoFCM5VZzk0pUOqTZs
/qEWj3z5+19dFyabUVsFNzHWjaCHgmk5TcS5SQrz+kn4qBLgeU8ss95LPsDJzyXi
3WAE5koa9B5E2AjIlg6yY8IhPqwGPMCZRizr3hER8A+47Hjosd6waRl+kTXlYqqd
lJ8ZqTDZYnl8PYA6yOz3Ke4Rrsd9APZpBNmq7U2GUNc4i99ASbZF1DYBsFgwQflF
XV/5HId0HUOxkv5nV172OiNdSRmy6pbN7a5dfWqK8631bhF+VEfzFV25hnOnmCc+
3qERM+aPNh+fHIKjDYOgpWjn2dRu2KZcx1yAtLf0voVivgpLdcVmzYdIG2P2lDl8
SAaP3eqRxaU6zOIWQoieI2O1JthNI/UIzU732xSOsFmnGcAwVIBaJeqEczPcE2Mf
JWICXMPJD1M/aoMYXTnTXBfQshEkAooV5JYPuvAzAImQKsEsf5XByYvCrPg+I0P4
4fmm42fBFIsZx2ErlzOvgWjnpo00BQNcLrUmZF6gRdHTd5PaG+lxgDhAFzAvEZAW
CPZ2bAK7OWrTA86T45//m8i0kquXgj/Gm8VDLNpHytNUCAIxUMiClOxGh3RY8v4z
bauqhG2C7EwVktqZ9jrFNDOK0KuhyMGGX1ElmjR9G6zzxI6RwO4o/xdkZtvdG/wE
hbhdk/kY0EU4MdLbFdFWsuwuSXpVqjEeNcCmNcdRZxZZoIAg0ArqDiCqpv8zs5qM
gjB1A1GwKOMMFP+ZbxsKE0FqHLrd81nKmzMHJVwqgjdVbim1wYcfW1djs7qy5wmS
apc6l8eC3eyezR3StXPaPkP2dr40oVzNe26atW6VB6t3stPgz/j4dehgIHHlEzDi
h0mNg1bJzJfiyWial6SeVfVPcMylP3WlF71cmmjqESkmCxD7ZH4VOcHuu5/ACYQc
6RDaaVpuFEgikvdf0pbWnnVILBr51oKmufTWuGMvHazKTEFDAXAgee7IvXZEfjkz
9GPL/FQvDB98D0NjdjXWRoWSXWmH8jKJ+h3mF1xbKWCCr7/NjeRs8L7ImelVqnhn
+JHsA/cDAo4VFEnjQDaOck2apPgxnsLMNGZfkFcAkFgP+eFhw+VqSQbPjg6kSIhk
Rm8vh7hOm5Bm/dJ3vUqiOFPUL41fmRbyAemzXJdePOcoTN0pRiiFZ7UFZd25u+OO
wenZSCpQdM8bY7eOsBskc66pFJB/5TAwzPaQDr6cY/QC2i5MViKhSwfxe8FZE/pY
r564q3dqC5Gy9menpuVjLzOoplyXKXLif2GLtWPOhitPfBS0QgQ9Px3DrMocY8v6
ECekcxSgETiu5pb/Vbe4h4hd1mNa8JSZqbb6g67j1tM9DqPGhjX6bHfUQwfMJgF2
mQOpa/IAQu2MbbiThyB+yWl3R1a/vIvw+SkXnj/CQT2fNNxGZnTqxfiqztot7uZT
TjNbjbOTmnSziqTZR619X+WLPhZ/G0Mdu7cbX6IcU8WTfWcMZqKnMP7YgsLysqGO
RCZC3H3oi2q+ScFHFOk42jedzCe7+/B0gEf4vwXVbEEt4CAofq8PzZQ/f/fN9d3N
yXyIT/qciT9IC6fVctEimk4JR5kWIsG2aPDFuqxksqP/INqEJYrMKgBFkSsPBCrU
LziKF85LhYCdpoq/4S/VTzSf4pbvxLOQUZX7VbsxW0iyGOYLdQeJ3YCjBVmKqwq1
qAIc8LSbA1H6evoXLO0Xe+B/ZaqnhsZDHBdMgCkAy25NZJl82ZKDgexmo8zs7dfs
t/N8RzF6utm/3F9iwBUqbBOU5cClzzPPaxkmOZwS9MRDhfzCsOZwfRy70JkJaygg
RigIQAwT/H7Tc5vFaiEtnhL6jXuUHjwmBbzvx7zQWMSVv1ezYd61LjVZKL+epuM3
PyeBycw003EczHnZFyvTQxmepFw+7Wo2dMMmIQ9gKQRGYa51tT06OkhYaGA39D8a
D+1b7oeF5qGE09DJYXgSaRMsB2A+1z4B0juNOsnghJ9Ns07+0K0E/qHYtJFu78VW
t9qsr4F5Vg02TBVGwO2nKcWlzs34S0rzQta2Ur5iyZeNhoGhRViCo2ioY/p3bT5y
q/+9v1LDDoq3IU8R2UpAMLQduMs1wj0Ap9HY44K20x6kvjMAwG/7SbHUdkhf47FE
RIYIoJKARZ8OrAeVEGYy1Lord6r7oWxzCGMuO4WxZ2jOHgrBkSxYS1c9j4P3ZWU6
jDYZWxHZb7703hsBTfCWBOjFxbHWAGW0AU7fHWJSfPXi2PTjfUeviAa6LQUlJg7y
NEbDzfWY3RHeJac9R8Q2h0+jeh1f50UP52ewz3zQfq2kz4tFb6TXruBnY46cWr4u
TgLkviAGUbW3xkQQL/TDEWz+SobWCCLbrOja2GL2bJkLtlo20k3Z7sksew0bqQsY
AIusfTYzpsuqdDvlcGkBO5CKfepQENWMIn1U4EQ57zlzQJVyJug4KkevDH3l4cXt
61Tmz2i5z93R0OkzF9GAx5OCHUEVi8JmE+GswQ9OIKRWT6IyY5t9veY+53pdwUyK
nfHqNhGXsHq8EgRFK3eHDms+ZzAFZ1yCFM8jKkpsrNvemZckJBYFkKQRBBiaKIpX
XqWVGvpCKW9eJilF7uoYh/4L9cpdH/OfPDAjw3MQme1njj3NOSXNlFVG7rpv6mS+
hl7fCF8jSEX/kIRvui3LBq8T9vJJn5p0FSILVn9Y3uxp9WJL6fx4bgDcugf+naTg
oZBJ5+rdY/3Cect23ReVKwDmXVEMfm220CY3Uw6eXRjIoIEDno8KNjgzxpceR6Hm
vjVVpfhv9xwiolO3F/rfaJFiTEICWcOGFGnYCeiaf1qQPXmzPyWYw2870zHoMaQs
XjDusKvUtjsF/Qc4XcIMmlYvZCZL7zEppyNmHlxSYGlv8fDKE2FpiPrfKEKdJyCu
noapFJUdvPMNEvSGz70h0BhggbS9YG3yTQSxAlcf6j0IJGMwUJQN2ww/rWZp65q3
3w4Jl7e2vcQMgtSjX7rKUQwUIvErrd9VK50XI2swanppadmLa7DYkMJZGyUx5ykV
YdY9fssWpORQr9p/QuDN/IWtjXchvqoYj1h26tvYQDG0qet0jAaon5/YEPs3vycU
4F6py2ghnn7dfhBB6zD+Cj7lbtLg3G8nENXyH4jdOowcg+eZNeWmVym3WP2qHQoK
hDEDmlo34A+mCu7ZIElMSX+7xRCg1Y5VYzm4kf9BVIwe5G69yEYouYphhAw6lX6s
dKGBgguzUxxR4mFG9oLO+eR17Fcunb0FFsTndtBy/7/8JUkDysXQiCgnQdgchu2z
vBaYbk0sDgBwT0yxQY59giH4S/lSJISm2vhS6aOyWpu59AE3fcPZfNrXbNiOUnVG
JRLvMuq4GBDNX4/9y2qNe3ay+BLVf3uLQyAZcBKivdU8Cke7YuETWAOp2XSgST1F
cdJLJRuagd1ajot2zcS7Ad7QEw6BtURaDCf/aem5EeYOq0zZ73AeYWX8LG2q8z/D
MIUPhiIzU7THna4My7B4IxBlc8mguG++5FBAY6PHY0HLXqLwf8YbSR7grLkMINW7
i3mqjXn1p2p+jg5DQHIGqj1jiBK6RdoDDdZLZsO/sA49RoYgKbZCA3xCcVPHmUTo
sH7+QQpZ12qJJBV4hZCxf2SaOKl6/zinX+cDjw9aipg4Zj3rFvOHF9Y7DDx2MjZn
b3Zr1LQU/ynpowSSiccsWcG00R+ROMiMT5wiLiyt0Ui9TxA1bUApJWWPeBO2yBh1
Xn20Y78XwQLa1hVY9vUFB7a9qBUr69sudpQnbN4+FSfMHge3bIWuRWgIniq1LqMn
RVFDcb8dkaQEW1Ihw9BRulGShcFWzOIsolOnsYL3Qbtrqu0uiDn6TpNKvnZxfuC/
Yg7QwPs0yLRQj7Pla34o5FJZ8Q76OV5NcxEshK5myZijSqVvoUdsYUj9ShQ2FCyf
Cw2yWmuL8hKX+6SbKEkA/z4KogrU5xQCud8yviFr5vZl+nB7NYSn9xMe+LeovKa0
Uu0szYfViQL/43UhsX07356Xi0YuPYaRMPnNHlUrnI9n3Bw69o4zWjdHCBG/akVl
EtsFG8b0rmx3uBSIZtzWTzszHuNEg7uRxrcLUHdwu2n00Pl6eT/DQbgR9a0/B8Hc
NP3Z+zU6I0Z75VoG7BptZEY55wahz89QT0HPJ+goqdOKPYw4WoVS6rAqeCa8OHkf
WHzWbg5IwiF0i15mtVhW2Hn+NJ4/JBZ2b/ce1d2EtY4To1PPf9BzYaNy/nhkefto
Yt1RSaAOPPOP21cNCMkKDwfGKFQNMpA43O3xlNCbWpmjL9A2zF9sucdVn+q2NoFM
+61MgopJzE+7TUAAReE82Au1Pf2ejqvzoRhsX8p8vFCDg3LpQiywMsQdbtifgNWv
rjmk0xgZjs9DQc4MY5KGGwn+hmnYWe3DJERaelQzdrn9+GV3uZnOKotEjyk6Nsny
ofH87/JEvYm81fz4ukGJzSYe7lr56YOWhxmGB1IekgUwXvpFUadUeW4Q13wUOQO3
JN6aJaABn2cpgKFoq+H725OJZ4zuFD/zPf4/Nu++x7i54EB8dlt5wW58oadm9IMw
oxnQ7RKftpBHfIHVbe0+b1fXxBFz5Oj6rGlzP2wyXk4tcFdXVP12A5X6nPhodA93
zlvmgGoThNQMTknTNPYvO9YG5BJPFu9rXbU+PGqVdSDn9wgJWi6JE44LKXfzcjNe
p3vECKqXIZBB1YuFMLxa223btPFuDZWVv9KPLF2WOZMh0DqkrkK0ccZYeZNih3xm
9zm6PaqnsovSAipa/tcbR5X7fW2kA4epXAt+aX+s8f0PjhuoVJE9+JJIba3zqNIT
Zm0jEi5/W7qkbWrTNGKUjKERY9XzAdD988b60UXmCyL/8+OgRD/65O8uM2Upok+z
W8O6M2ZDwXeExq2IDPt9DW9I4bX/DiwxsIDHq33R2KkF4FWHiBcyOalmnVdboZZF
73/yeU6S6DYhuIP8IyBo/ZF34AHr3jTlJyOArVxGqt5MlLh9nezTDoLLOBCtsLlQ
vkKQSIZfFJcGIeWelQi1H9DwbaeKtKIwp0JszIeqgXhL+At/QBOS19QPjUqp7zDb
gB7Q974v5HDcsf0cZh790paiFC3bnriJj6d3p/5royFzxUTD8OHQVYxHQhBJ84ga
DeF5JZ5d7r6BjCDWV15VjAu4LE0yWu1rOFdkVRNxhjYM3IFRt8jZktYmyC270N9k
xV3lIPyqeFu+VHyxL3DkZIv7XI6yCaQ6ObBAfPKlNKIxUYjZUnQbl6PAQ0E19r12
QlbH5g8o1il5dbQ0FvrCp1MC7Xu37Z7wvMPBnrDsRoiRLHLeQuXBR6JzkgmcYK1t
0o+lFp7kEYXy8I21o1O8UW5GD8wFxOf4IVGQJEJ/m0lTCEPBzsjk/Im5gwGnj1sm
hwhfN7NgmzYYt8X2cpoPT8R0/UM2f8POKQVzZpux6gm4oLYP4RlfJgxi4Jd7ywKE
E4G4ZtniKLwvn/FSzfHNw6xfouaiR6mn34qIdB74URFVRMfsRbcX4jJUpfokK4n3
A7ED0Vg5tNgZaQld1coV9b3eAAPi2tNaczolJo+g6ZcEd8G/jHNKSuag/SbgM8k1
piYSH3Iw7p/9EpfrSIDcbw4zgeVyiIe1m0WkyKbzkefpb6HjELnX4f5PMOS7BViQ
jpi1y9DzdbXo4N49ZwWqHbNZaJR/NB8UkkSIz809LeXb1RLY5qDH7wK2jkGog+6f
4Z7UXGbcBmuH4KGJkvY/pcULDymArIWG7v9a3S1awqH6/FprrACZGZPnIfWbvTB1
dcaFKCebeQRBqNsEMgHNz8O5V/qqwD1jAzrePTYeUmYen9aXjA75hEqeaIli96nR
HzREhyBupnPE7HHVkW7zmzGfjm1tNzk/0eGB4GwC7iFB2VlUJSmRL48iezGI6eex
Vs7Z6M78oayRx/Tq0KFXJim2DPoLz5Kh4TNcehv78i9pQ+Y3Zzjrg+/KsDuHO2a/
ypp/r8NbiCKaG2A4AicwORlOKKKdQh+82Kt587D2GW7xNxoEsusxgm4ACYpakV/m
iFoYKVPvtRCDng34HQf1UlpUsuWoByfkxFIEAUcw6VlUxp41NX4c7R860gSneQob
PrTwAO8Nou2I23FxyVF455vyWOVujv4LOwLidg8A6/FWQxbGPx6yV/yo4AgIZFTb
SG4WRps1ZwQGGQZEW9EH50YvYXNZxzok33ZToeH9SY1hMnfxTg7MHvzWaYGdc0y6
EJdPG0GOCKRCSb1ths+vlKqoeVhG3wldzSqhCWyx+7yDlIiBHUsxEq4NbxWngjdT
XQpj74MTMbUFdtS/2pomVXNh+5YLpzLH0AL4hpcuZQRcaqdkF+WAT0XI7maz+eTi
HoVPKNMF76xrvCI9VcjHT5lPD2EL7ck6zsTVN17JSciyxmHrgawcb7OnJNOPQ37P
RmROn/9SsjPdZDMAikYqH92YEwHL16h3cE5ZCR9fw5agVI+0uWsOmXfKe9q3aXFl
ORcdpVcXVnKQsgyV0BeyXcXoWEXf4hDg2izT946+omAC2m/1RrUfSRbOXGsnGZrJ
VLGv8rtRkGnFysz8jq7YOMOC+7VA3cVSYC3tER977rDVXgIZif5UCqW5Oe4licaZ
YpE16R42csdxT3HyE3e8QJoqobaNT+sN68W8yXKNGYRqg7AZjQJylpKcxqGx3p3W
Q5s2OKtWaRcXWsOUQvfRF8eCREbBAjI5TTnfwwGMtZaTHkvF497PjjfURVm2nzrc
mmGnyYDiflyhMVU9W+RvT7o/7OASUfpOKrykNFSWRwpZFgb05dIbWSYZNZ8QsCH5
ULALBNZb8as8O2vFOYAf9SPNKByJZjUTEqqq8G8NWTpefaMBum+V4ZkTg5Fr+1BN
Z6WG01bskZyao9XtwHi0i7XzoZoLk+8+3XEJbCgxl3PXeDzUS+nXURLYU+5OEciM
GXMq4hXO7WOy0F6i4a9ps0WKvskIu2PgNIPaNU7FetV+hA6bnwr3oM1ts9Akxx4+
BF/RD1bk9cWQUYrSn0xkMODh69amZ8++NHZNZg9HaDpcUMTJoxJhkxSETeQxMNmw
KEKohcsw1RkeTBGH14WKqH2D3mO9NIQfvkuIL6R0VZj6oJB8FzqUMsRQSHIUTA0N
zpBFSY9JGA/0SYS4Qw+rt/mT4Xx2YfBq9c+HPIBR7iSo7xDdzgZF/HLK7fO/pDJq
ckOEcU/hHF7l5kZ0xKTjKEFgQ8aTftazGt90AlTbWeRLTyPXSnUHKosjO1iUfc92
bDHp9q1Nze/IJe+4F77JDdrAnhy3TaY8Z1knKSrGr5zm7UbM9+7Ckbr9BKhwu8Ju
dEj9a8wVtnOjSs8QQMZc0nX8YZiEZmp+XIdw+x3AqC1is33LftoANFRu6GhiOlLH
/Q9z4mz4UZFFY/YbXBjUsA003vz1+skxAJ/q727gkyCA7GFkSEKeQZ/Kzk2LNjUT
5Ayc7yaY7qsT3XkzrJdfEl/kDhhpNi53x+5EZ0DteUfqMx2LkB8DqFLbw+NkEVA1
Pjy+3yerQMe3pP5WBgYoqRB/e+aIfGbziBwguts94exbAEhhEKY2AYxdEBAV/SRY
TUnl0W8FzQ1WVblm5DttrLMrX+4hNOTQOU6zkeLRaz7QiGC1xs910z0delHpPXhB
C21eGZIeG+Nc3LGIoW5X6v9MFO1Ik1jSqBZfS4RxDU6M4d30nd6wnkMwK/kFB1HZ
+8Xiz0kxXV/49K80HNijlPCHc+DflUQDLUq75rf1OnsxWZbCgpl+5be9Ix16cqyf
qUluwCNGr19NtVyFuEEiREmrkSoLMIOnJmV53abdAMDyxxEHZKUsglOmimEJZt59
seeQ5F2rcg106DJJzpbIJyPbJSxbBM5Mgh9gZ/RbmwIdO8uWbVE8AXizSNtZjviM
3SG5ItIaCd8k/baKGDl5PAKo62QBM5hU1VLUIaGglWWjfWmJbOrHeRc2NKPodTlc
STBTXANAprDhzdz9FD2kCwLO83xrBay283GkHqZtVWeUdBCJwFXl0s+IabK3R1yz
FCdPrBJTOT1i/WZ+zVbK5R7bVLJizcbMoj/ebCBkbht00zjrsBexN51/DbBSFj4j
TlQAnMF90yKGSUZLAYj5nPD2RRipO1ozpk5M+/ixXmRhsWt6e+wRvzRYU5BMCEIi
thtLnHM7ftFZ21pAW1Sberf+fz5lrtsQSra6dehCsVq265z4GcHODnTKo/BlP/RA
75o1SJat8K2K66IPrbdrT2GTqShjg0RKOVpyTB4Hhl8ubdP7tozCJQcvXvhoby34
mVcHCvOtMAH4nihiP0VSyvd+BxR8DaWsuMcEhntPq3L28JAIa2X4vnb6JwAZ8Yu5
8t5zpLwpCk12zS7+mvf5+pEEsy97ZZRcdrvp39ty9cs4PPZymQiJCloj6l/uhzCM
iIjlVDZvpbZd09rsQScQ8zuj1RQVV30iiZNno8OIo87zHJTzBj9SRDhbyyC/XSsp
lCsgxyXmvAgYaJaFhoN1f2zk4q5znvKAo8e+4CPWST2D0IKsLbGf6GGlmk7DothN
iapBk09NnczGw3d1sGt4qRRtbHHJRl6ThjipzPsjVd+aBLM/A8PBS4JLIQ9ZVaI2
PkPu7UuCzfC+BlNZ8HtWxQE+Ejjj9EymniD8OELbvarhHyd31HTTizljYE+XLEj8
G822Ha9k3ufvqvGBOyhSlS0QacXkaVZ4d1CDBZQwZu+gbnz0rfK6NeO4zkdNvUZY
5m4heFYGUt+aH4oPN8xHovXHoMQrGkRuVqNzzIk8af+LIgKav13xOx7V5/lTs5HK
s3hx0AZY3kIrC5gkdTqyN4dxWhKpCVXiHP4Jy3pnYs+nPUrnB4F9SDK92Jmv6mqU
JCpf3oe7uyy/dKcpfCQN44TUAdSiQM/0SwxI9vU3HZ/M8+labl2vWjpwhL7512S3
K+1B3JMrLiY1cR+9a4oSwkUhLJ0UI06/PTBtwyvap7lKBvVHJQ43W64uEXOzQUGi
ZqupQRS/FRF0aHoan1XJQNFuhSfo6cHZmKq+Qa/GC+pQtz59Zv84dvpQTruHtrNM
930Ij2O5dii4XznRBgRrBN9QTgJV9EJ0AqzfF8TIc/aWfWnjWCxDTjRUl9d4jQQj
o+5E3zrtdLnQJopJwKdALW9MYmDGVLrc536KIpLMsEB2p1NuCFyBmGwledy9wZaT
dRFqIkPql9OZVd3Cwa602EgKAdeICuLurZKj3ghdP1fc9CRL7UjGM56AJl1x87PX
2yuN1krDH6eHeMQGe+5qI0zgW+1s4Nt+h7HhZ4DB64wGpotT2/ZnX3GBdxzQr4v4
8y0vL/qjxoVEQvvFqIUPkAXC5/gv4sJVAlE+o4ykXEQH4uJ4sAK2/LSy9+dUKoyM
L1cJrvc4m1wTnRIyC2E1rpvTnykLFWw6HeEr6cXtM9cGDPcq02Z5l4BIpMtQDW/v
LbzWqwcapLy5wBb/klvb8u5Er5BN98sy5vEejVVD+4ZRuGp23zDTvn622WhrSF78
5ArLAl0HfqlIQsPaeL3td+l+YcJk2OV5pcGmXoSf/VDZYYRgOY6CmqWQieYWiynh
8c2/8imaLHa5V9R6zWOHGaqBNs5cVxHERh5mNtPmFHU+R5h+LPwptBL+ZKp1BHjm
6PJoje2BcbYeJJ6K17a3O0d7rcXX6Rjqig5H/rA+KAzKeDOcRAMAqZ49rrFgK9t5
WrbgLT6HZ96Rq/HRTFVfeTOhjCPDHfgWKL0nCOAvGm1aK+ghepElbtRfSSj28mam
hK17JdNJPe3hxacUgCg3NmxmXVbEtK9gt79WJvmWfLCdl8EroQJCD2oBMxFTVa4A
6/CS4WI4Tdm0Wg5OI076SrzjneEuVG7cDUI1cTAYjgcmABAgWUxIr1VewTYTDIho
sXNUg3P+mIj0nnEmlJq1c0TaRzkmQkp8A3hnDvYfSzI1xt5OPHtRI/wzcmRSOGWr
hMMFBAZSmQnNyog39CyuT8tgt/baAqqi/WdkY8JutloW7Wlr22irEi4HSiqya0gw
2v15c1W0JTDnhSiJqmOKdKm2JcNh+ix5pMDpJ8JR0tIZCXhJie25F6xKHfCOgata
4dUhnxCNxk465XY0t1/H51aZNxt7EsizrRrP94tPKgyFpD5wRN6M5i1fyqWm1P4B
c9ct5IWpZEDbUxeOtWcttjWcGBH8ez2zUCTxpV6AJg2ET4yyt4zF8S8drFIkFMke
XB+w25wUmAWW6ccwvKYe4PFWUa4KNh4vXl5+NokLtGpb6tESjdmCF6sTqMfe3KdZ
mAntslfzp0ojT+NQUqdAi2wHwOt6w+T0rFnPy1cHmdzGwu/zHfMiSAYgOUa8oIry
8f+b7gmAXi81PHTRiVROPOHJRJL4crIJKRuagxfHILuRGgaMRbkHzO0Ty65ie3oz
nkbshFxQGkQRToZ0frIvyEV3qV1xWTcUYdWFj3vksrMJLfLU6Du+Ulh9wb7BPGYF
3DLNnBMpzdgdODYKBE0+RqkD91jQIjnA6Oqbtogcqre6bEda6OCSslfyjsz2xNJi
qCtGre+4oyjEUUZVAIvE7CeLksrTJsqXdShdw2DoiG7to9Q6QbAENAozl551Pzke
376ZKejZYipSOjafHPNdPdEBt7J09T9oAD9HF/lNe2s32i+aL86W+ZYIN1BcWxU4
36cZFE0hvUwvnPTHHWZBZINorMCtk4TAQKT6QYKcr7ZY/jAysSWWs7KV7GPsvBRU
Uv9rx8y+pXywWu6UylXjewhzVtqaaqRXi4xrQFWu0h/9WLQW4n3EJL1FWOC2Gb2v
I7AfHfROkojfvEm3cxSFogMX0kCaz3RL5FY6GpRdFEX3OSG6I9C23Trx9y2XH8Ez
YxW1tXnpmgjLSWpTQLRQQ5v8PQoLzl3wb0mck5OS+1+aUP7iCd+BTMMyYH+jpVI+
SPjsbfJqX3Zv9tPwbiy+6gyZquuTSfJQWXATq2q+fHhCi0DrPiOr+qQVss/YneKA
A3ZgAcI+dRmgP2asmHRnzmfuOYkDIwKnuweUfY2hW9UZrznyd+LTal91DzbBPOwl
98qmfn6g65WTXZYQ3FptRbMa06uVqfWabZ59zBgloNuTDxhd7qR0jSafi382ikfd
uB4bCXObQQvrWVdh8W3Bpipve2geVyReY4UtGRwWjIqFgh71tr8Q4Dc0n9Kxevt1
Iu1i6hBSLFUDzGHHCa8+r1Z8/pTLMG1/zFMzYEyoPces180yXMmVZieBU3a43ucV
5VBRStES4roS+lIZEYXqZrYuS01nHT76HFcK9QNBShwdrR4Hrap6otJM2G9wcKtI
t46/xkhUDfO1KJ1oMT7XI8cLMzmfewtEirT94fiXgR5qDKyyMArQRlo0DBU1/3VS
NTHUPizTIy312lC+cTGRKbywm8bacDMhTEkdbjg27xUaVExzIbJiTQvWegZOdHq4
Q/h2sZLyyZYIH8xwggeN6De61378vPyCOnHACjbQ3KEqvCriix/6r1YvhGgKyLtH
ZsCKbIR4yBbZwNT0aXG7dutun7bwCPZqGJAfobedizTXbI1+1E2b8uE3M7vlFoN7
3SSwphjVi5fkwaHmhrpdOomK47cJURuZEqcUn8XpmSyjnp5DtCbIyeGWvs4+Dj06
2Js7Bz5muwa0B7/X6mXOetDmxqbTr0IgQ2y5k/MuLyjWtcDOYQixtg3vquXNDbFn
cm2PEtRGlE48enabVPwp6wJAwnfcR/SeeFd6bN8bSB6ujPrl4gK3hyMtuMryKVuf
BMA/j0yzrhHBorARV8w/C1bbbWZ/5yKJOFCsnXcioaccqQL73Xc842qDe1V5Fff9
om51exAU5Uqdg10bLTXzaa/ZZUJDqoES1sLtHAnJBcxyUH2AgozvAx0dOWkplxAg
lfNkvesNJJCy9WgTJAc9rWdBTCIhjYTyTE/og/+UC8w6u0D+ZQhQuAcTAsscXwMh
Hegt355l20w3x1py6npHCViz0ZATnW10AM9AtCQda4bQSVLBWnQuLBQY3RpIsm7L
lteByEuDG/dwMEH3c5HEahH3O6gxGAS+C+GogBiEwuAiIxKmiVwbMJ2+nZfY7FZ+
0fBfV3ZLkYhNXehtvQbbHUy0cf+6ZnfD9yVMwtK4vfw5l4bdTTNiJ2QZLqxJgMq6
ixhkmYn/CWb6ur0cH0ssIoQU9mA8yfe2hQL618KitJdwwPCuhzxCvEFgV3fUIV9b
JPh84JSBcIvN3d2Bv6vWntvVqmP59CT/S6IprNDRCJ54pV4TRMr7Oy4kM9A0Rfap
TRms0SBMMHlqtOUTpbQqwDAGQq8U0cojHcOMbQzeWQ32nTcfbdZOzCQbvoSwB+E+
4lQh56YWDZlNEDYpE4hT/Cf6Pt5U/biuToQ+0YUrIRtToI1hngjnShKxN2mYg7QS
B2z2bZjkah2C+d6+7/05517zp3dBPBogS8LP/FTsZhd+v9ASfy9DuIEZxztrosAp
kp7jjdtC47qnlj9gxWqHBmXhHO9bjrv4690CqK6Dq+bTAXvuXFE4SaJ9kPbaf5OO
vtZauBlWoij1P/Goebe/4aM4I3vuO4iT6OLuB+qvXwF7Qz1ULSuULB9iQGTMRjHt
zbKR2hwooiMHBEGAlmToSF+BnmdRV41UzRFYiozGDrL9dnEiYNWCyVoXmZJNlOCt
76JxP+za0h83Et/pIjTqYuFVLwKWcGUUxMCirk47NmS3INQO+86HiCvgwPAw6CrA
ycNCqoWKYrNUSNhKhdSpQKGv/fhAzLO9NT5nOHd5JvjOLcfL/+zuui4dHzCkeUQ9
agJEc+pod82nQcC+349AlUdvFoDK1PY+Myxg4Ig2HNnHTItbHX0jLKM+1zByV4Lb
PBnyoMWQ0o8OVs+gnZ9VmdAv2T8vrrTEhIJ/OFHqOA4cT22gX7Sr/tVXqGczBMOy
AF6wp0bwmyEO86qWoD6jbHFLPwP27QVEDiPEPDuWQJIyvlua8IR4mXqSqvaoHR3B
jp9nC+TK4HNmSCpc9sZ7Pagf0mN64O1ZLabDyIa6d2H5REJDbhuJRApxh8LFng61
HKTUBq3w7omZVasB4iZtTjKPcI4NllkVx2ChN3gIonhGZN4QSTImoB+oE3jfewpl
54HYfn9HjMg2oa2jJGyA9eCymfOkjVsUUaS+0Fe7sGYYa2Mpkl25zktojGQHnsh8
2u5Y/+UooGhxKSfmKomR+NlWXZgEjES3hp93GCvnUByUfnMctffCk1G8Lyl8m6Gx
imqmKXWQx34U9bLEjOfW7l2tkhIsDnOmJlb+NjfJqvud33O3sTI1HmOhTkoyomCc
4cfae8SYITzN1kld3SiFEXsszO+wOlIKiDFS/cHZEk7GXQSd7fuGEmWXqNkd4AY8
TJLDzOSfLEHnDjr4CvVd4lu/RWpGPoohoduAnf4NjLquxW6bSI5/lWLgU+yvzUkh
NiM4qvQ4MuTnuN/4dhDvQtZLaKpD7+a2J6yBRge7FjHtoS//3WAMh83mdyGfQ61+
fa22BuKct0ptSw8n7uj8dvh8w3SKeTs1mDuKK7JiCsL+1LfMIfxBxw4aibKC01J4
cVgiVuTBU6QSOi8FfWiB7e+52UaHcM1/+cwlSmxrnAY1rBybRp2r/nrD36DGVcrq
INrnMY3MmLh8e8gOvDHYJGSJ42rS+xtQsx/2j2TZ+rNZNPTb6+tGJaJiICILinXf
tvxXVU1zcXzN3dOBt2Zwkir7ZZv8jQ3AVGSgJVOuHwCCkqIMZ86sa9JSaTG56nKm
nSTIylPSZB/e0bZiMVmGWYCuMQRsceyXv+Wd3yQ4TTprvmHbfeM6FlXHlO7AmQ7P
KeRbBVXSOMTNlFkzoVv3CHixRfM3RyQnAn1eXvIJofs34JWjFft6uqBxMfojf0rD
8RIMqFAS7Po0UptsKk5mH9Lh6Vo4dc5JAAUCdKjK40UXB8HGO5dM3ztKQFeGK6fp
gLwoHGZkbu8vYa0WAixWIE/IoO54qJmiO4bAj6vRG5in0lBaURL9FkSFQmdQ7/hU
Ae0ZQXy8W+BJk87vbyriwMQc0wtRvFIJ1hzrBoHXSNXkXcUlQwSk1V75j/5UnGcT
DIRXEIGqzAvKo2gpfpEvAp0rmnLW/cG4NDNElN1AOtGMLoyDcm8qlE8uawuhDzWs
h+NGD9tW7Q6bk0MPo95jcozvKCn+3DMonj6uSmfMyyIxuIzZMxQMAg67p+ao3KIC
Vw/4C4j0pnUvBTq7Wo1Js1FMhhJilS4hYR61Qbf37ecbsL0KLp4I3W0k6ygt7ipN
aHORdjdU5ACK3XMNrzUChKHKsPEr4LZHboBEU6C7PfxxQlhSvVaX0987hvOovvEC
IZcroWWCJPjz+UUa3XugTk1oV+Z+KT0LD80TS3d2qC0j9SZNRLf8WfFW3VqDqVb8
e1vmNMiTug/H7RetdbVv2FDAnwJwWBM8/blZrqaFc13dZ8wOf2/eAhcE9vzF1xrF
YYeqCkZn86HCNhbKyovA+rg2BjSe6tUgkboOPs8/scyJ8Kc35Qdqrcc4JzibEIRS
79iFEwMn9ioLpX9AJOT7fskUse0pXH7zaX4dQVvPbZxbYWu2fFPJAntHvkq9ywGw
P85S4way+2984P7Z7h6n+tweApOtr7tdYn9CCEdKh9vcxt2W1QHAAYHm9yGiwlxk
VdGYOyZ3GM1QD5eDwkdiEN4If/OTw5caA/zdBJ/kWlfRdXMF6zyI+ht2tws+oAdd
W51U7nMksFKnjZAA1cg6BD3g/boH1QroR8cAt9V+A0MRjVF2f49TknsI8sQjWrET
X9ZoJISU5Aw0lZ5ZoEqteuAXTweeX0XAW7M/jXZaBKyo3N9/SsSW2Z4EuhnItHJF
vYMMXXOWCi7mrYeLwLARtyCJw7zHr8TTPChnDtPHx2C1/M3+XVmeQCA06pWYz5vl
jFxfVn/oMMYoyTfWi8efMDqaN8NQSmefZYwKz1qu/q52cxeglm04r8ELInl0Ygnf
5xs3NSfDCf2SWSMGxFv98bim1++JU8/d3sU+MF2Uz7IPZDWKLaSIMWUckkbCKVRt
OHd8cc+CRNSTaTttyBT3Y7V/DWfIS4bCgf4qXSKoM4QHlcYK40fRac/vbBSI/dIx
25teGBToM3S41kP6WOBu5mh1g6MbS1I4FzMgtMCWRA5Lbki1neILDVqCBeDeR0/i
O1+ShWfM5WeulP+Q0Znfa6igrj0iRFH/WYEBHd9u2trS9I5uzFIgh/rIAQZeMXUf
tctYO3XUMgP2BRXTgnF50/tWKWmryfE5cxTuIjhK8gumdCng9WGiMHVpllvEkp/U
bBmLhXmJHSiObtDK1UhdjnGJdqIWKAAuIYSponR89LXWbRbO8BhX1zumudk6fXG/
Xhr4FVjJNkIT/Kqg4z6CBCNW1hWmL43U29n1pxj5jR2mT36CY+U0DO/a7QjUTb+Q
ByZceZ2S8xENP9xPFHboOB+5thYB3sMm8tMlqlaaw6duhPzhpga2oZDPrkByJGMj
0fqa8MRooDlhOfSFJpkVTmAcvS01DvunhJLP87vtCAnncljxLt9beOENoYRHM9gb
KC7V1DId2GO/PvgP14zc3iaBRTwRVJGv5eGiC8uIQ1Hp9MvIi3kzk7e6E8JeyCoS
KRozUh7XHVxeynAn/GC/Tweq+i6lc78ogWXZOS6aqoU1RMt+YpMMaXIl/uVzFUKj
GlRjwsXE6jNG01VnhrJ8cicewYMgVzsoqZxkcYxGzkdweFbcCn8e9W+RX2rD7J+2
Yro1h1aUJd3TEK2x78QOKpvQyL/Tq7M3uZarRS0K8pU18uSYxYHnZWHChg3uULpj
M3N+oBrOZ/nSZ09Qbw0XdDk3p6GMeAFaCdNVWaVovPIbrnhx0CO6SfnFfmUOBDuq
0duEjgtOXTEpiMKmE/D5apmvgzKQm++nC8PK4vtyOo/NsO4xoh86hIa/6kOScrPL
9/7abaDAfsNpnVmL1hCG/Nv1xJ6plytvVQMqzJ/+KXtL8Qw+z2sGRdi3Fdo9EfDX
Mp8k6xeYzZxUQkN4AVYy8OgBWeXqW1oY41wlM97jaaXJaWfl7nmIJCpwkbh2Zq9k
ba/izoipas9zcOw5isyjfj6Z70Ns+62HvSVPAOqrOkvn202oc7EyHE6KdrfCYz3M
qMALjzBCHrAIpRruk9jjSKbu1z5c5JZXl9kbi4biJ2ItPyuPqDF5NZKpSJdKLa1u
hWgjEsaMiWmL6j+HBzfC/wSkuyz7RKcyHKt2gc0WugYvFvHK/jh9uefpvCHJzwMH
QxcitvrOZoMXEqlqDp0fD65eaR0IwvSSdHYvKqKSlAv8k4fmbs0dI/iSx21AlxUc
ylaLFBlX745yRf6mEkCsGwz04GV/MiXH0tQ9R6HyRhvkZ/kngcr8QxHgeKUt1JDT
11kbDMBQUfJ7fnk+0LLzUvnzz4GEM6UAWEdnt1nR73765AsZW7Md7zYP0pJiDqFa
1B5tOllbhRiyqLyVlybERXnREtW0Lra7pLB0kISB7/hBB93oVkSqoz11wvJfRYGA
OPutkEB+cSCXDUp0Uw3Dm+tBKf5Cj4EXE3JUzQlzchugk/0VJqedDPjidz1MgqS6
+xP+EpQ7L9zu0q0MKHNWJVZp21nm44ueo++WvAomghGI/vO35N+66pBS2ISztMIw
Bhp7EYE0HfjB9oHqBSLOtVGe+wT3feiwdsq2hwUlBvbIn1YoiIdULnkBDneR2tGT
XOTQ8JHuDt+jOMzPuokxSksDZnq/bYy40swThgyGa+2/hnbDBN7nEFRX+PPpivsa
S/y2PmjBFwvlggZWZZwkwZY74mhMzwFAS77KRT8gW/Ga4B9ORfU6SrcIm0EmfLp2
IoMFmZbf59ueKJX8R+QSBnWLzgldT8l2Bet0ng9q1iVWuqAQnBW5VTSnFmBa5PXd
qjKRCj+knrfVymcFeDOG6044QHbNxhXa4ueVGJUuEM+jukFvkTPStTb+hCR0GsOb
woj+Mx2GXibA+IsdJFDJu02AjnLbF2jetigywP4jPKLFUNk5b9hVpX3tEou2SqLg
0xXQS4+L6iVYqIu5DWH0Miu+THDVXQvJkXGRMT/A8IseDjW6bYxYsGy2jcskpxJq
iNLjl23kWP+D777PgJ3q5mKEjQnJYk8oc5BhQM3uhOpGByBv0zKFrGZlowFAXIya
fCZ8rlzW9QZepUNdiKxuTKmQigvtm1USuTWe0x8CgaHrFGEaHdRTk8sCxAzcUGcP
j6cIJrAaLF8wtNIz3W74V+JJBzCcw9ydNpvz/DBXGdx39cLFjytN1oURBgyVvtVi
HI7ACIX7thaOHKgBUJqymhUKpUBNkOXEr9X4CXhf9MZsXy5QmrGLvW4iK3Echp2N
Axsk/VWqXL7u4c+hWZvIELcKVuXqnJWH9Gf7kDhnV4RFhInS+/HVS9fqptA0IM9q
pnDtsVsemGdgSOqoy1lBZlUnMPCd092+RrSvcsXdJgCuKL1KcIOSly99hSh2FAET
1TW+jBzLhIdHRDxsS5b0aQD2kDs2PoxGCNrc0BlJh/Nm9XaP4MkNzk6qjuR475++
jZrVxi2S1cM+9DUZsmZ/+QKvkPKZUql9JI59VKxMPuDjDBB7WZ0XF0pTCPpPeRMn
8xnoYUD7x6Vj5on9a7eqLxYRmD99KvTlClSzTlqkarlDKYK5t3NXQADziC+hGo0t
PyadXE+3JIK0LarHZs5Z78E5utp79JK0EC/1WX4L+Kapf9FrkMNDfrbyjM6fQNYa
fv7jhFgoyFyED5YIeuA0VbE40sb394wrqhOG3U+PcesEWe3ROzpBeC95zPw2r29o
RQWgAjPXMs9LNoSsqzEaFeEI+UtgM5RTB6d/IxnnRFbVBVJHUEWYdHA8t4jelKJo
m9yfIuiFTzMJYB1EwzjooiTIgj+adiZQXT1ZRCtZQclOzbLqluCJSDyHhHoCAyS/
yMdFpgU9Y71If5QQM589+qT6ngdLOFcpmP8mG3W0Qr9qt/oR5T6Wj5L6U4dILlEO
AbqSEeEvZ+30XDxDL+Irvq29sGo93hfZXkk6/QaFUIc7V4bEkmMoy3INBd4FDhBE
r3KzyKzcT8XTgGSjJarKt/qo7SbWNOtp+NxlKlKzjplhERWuMRGEmxXAMfHLTEvA
PTxUZZLtf1CQ3RaGBHgchns/Dg19021uODIQoV/aM+XbLjhuQ1LN66WeBouVcDwE
1v3c2Ykhbo/Ldauh6bXqWl6ibJJaiWgTppvdNtqXNKTAdzMflRwNIjaE//o/L0qe
dFDaUxUi5Q9VhIvyDY9HLhwjMh/htIhY2mFvgL6Y6DlwsixCBPqjI36uG9x21vis
5Nri585yu8biIVFYpJ+L8zAnoi07ad6j6DQn0F7hYu6sVyen4JHydeV3O70PjSte
Ru0FcmqcU9NbkCj3pi/BMfdWJrqRFdtz9Q/A2JO95wq+H/gyP1rYhTE7VRah3yzN
JXUlTAO8msPqly89DJu+AkvoXoNcBT5o2JRHXFMQvl2KgrxPiIuOnnx4ktDekOvT
K+nBtTWFJu6L66DQkHYPXNOv4MD5cbV54UvEscT46CUgPyzz9SpeTT67/tFkYEXf
iW4igt0rvPJyB9GIYHXmSeG5/Hw5yMjdJkH5rPFiVw7hxObh53TDZStS8Pmy9UXg
5zrjhlPa2Hvh9OpDHJIMQ/DPSvO0p6ibB8J26w/ZJrK8Cz4Uafm7/ceWWfr5eXbO
3OIpSM2ia6PUGJHo8fNDD/uJSkl8t1N/Po/eHlF+/U9pWELPwIvPg63iRuA93VFq
bPJVxHDOOWhY/08Fp63hXM62g5uam38abao4LRWdv9/NZMjy0KuzXZbWwvmDaDIK
b5p8n6nHU5BfCNzp5Nqglfu6A7rw6UAuImGr+WoGldnvcnka7US8pUuY5raXDEaN
lGGfiSocI2yeT8RxkFlC+x/BIa/C1rHBXp7LPsGg3sU+1rjz9ra+7dKuZYd/sRqp
MHpyiVzDjfzLug+B/5pAMSB5JYBk9dYwhwvRVXcnq/2G2ORBFklNgt9EeCGLhx9T
CKx4TcrTfvX1LzsEiB/cDjZqbeS5lufYWFvlrcXW6j7knLGjlaH+i1RJnIsTgAAP
m557KZO2ln0F6GU0kv0LXwS2BfLA/DymAwuV9uHBMj6+4XqNCGzK9QFhpISwAs5O
bldqpd4iO3tuaKewT8kDNbVk+lUAXPSUOZAClXqNmzoaZgTzkX7xKwzf13pgVoVu
ZvnYyLoIB7z/9Yu0hxnI+ZbcunZvLJPEOhUt6Mn+wKEVn2kKcwbG//7DA0X4kRUF
yFDeZFBj522hDleLSkCr5ajbvt5f/x2jcd0lpUtI1Bhppf7GfS8Sur+AaqwzAZsu
zAzxerEKq0m4V58/mbP+HzeNmzHgqV+Y6T/ULyGcDOe0THDjbaLgMTsHRjosVnYU
lumT9THDz6OMpMnf9/6695mlz5srJs7IRGY7QP4RDBZ03DD/CBA4NiZRM5YyEdYi
TRllGyDMAjKqZwjgiJwf1KyzYhD1YegbOHNsh5Yo2DUB/ddo/79iVqUbcm3ptHqz
wsi/g9wYnjWmOFCArLpmgwbPBuIUe7anJDgW8gBew0GyHOBdvlsTAN6yfAi8Q4Bz
8zqXdSrm1R6wt4DtBlGIe4SDs0JdQ8vh64wWzHAyEv6D3tBip1dhjQwScmzaL5No
K17KYb9ofJM6vuqA9DC4Uxb+Q93tBNkVucz+kD5s/sMDOnvc4+WZiSVRBfwxiWZT
1Um9neTkAvdW00a1Hw7eI9Vheb+L9ubZSSwMu3asRRJ1fPEmINGj94tj0XRjRKCL
ShH/akCe3HOa/LHaIADMZBw8nXQlFhdry9mzRd1UshLBBbM1J9nooqZBSKPqLxYa
PALgN/U/8+/kPHLlXaw4XG9ox9twg8O0NUIiVOlqsQE7oogomdRUhtkexIq2FnWt
kmGmI3e71jV8vN2SNNXNbueydXKUVrapyVNug08rv7e7gbFRIQa+WAZL7Z9kpOXM
GW/a6T2Z5DiMLPHC3fEpN0f0Sn03NEL2DsHhKq8hDFOUCJ14Lh+MRScvz14oBBmq
kSJs3ssInP7x8VwZ92Ot87y97g32XYwW7oTvcV1xQmJT9K4eI32rLjI74musgDoW
ViybxBbOuvLCRLk0CZHB270f8t02MbVhFqFYX+t+0yL+kMr+hFDIyV+GDo1PWwIL
hKPlSZ0tEmAWRt+U1GmUHQ+OEJ6acKzWMI8pHQU0z7/wu5tWldvCPx2AddeQjHbB
YjPsMCze2GjznhK5R32vbz+GAcIkeF2rPoacvj0r1a4tcrlrPzcOMn9Zp1AkWxrk
Sq/e8k92UrpQ7ZPgMw4IFA27Kqn5v9cwvv5VtGukQTQ3C2E7BjVCdCYtu19qGSGy
dfnpcVfo3yCUVhgX1GrJnbwKKzFZeLBF6+6lcRqUVO3bY7s5JJGczVTFTb6DlWMl
4ls5K/a53MLMS5XeRHPWbA8gVRJF82s1hZINnx98T8LtRYd/PX++vdM7E0ntCsDz
7IFPNMhQAkVuYiqAl3STl1VTCdcgRxV0i25HlUeNYBoa9svenQGcrYkejTFxpXaC
EBbqFe6ISu2B1vPs/5fVs3kke/D1KwXE8ftehaNAHg198JGN5CzZ2FW8VQ4RaOHg
hvokiuzuPUGTIOm6Crym5zhdVFEp+SYImMbIAL4HkBjw6fkEW2U9H2nI5w04/OXX
l0/bkZ+XDYDxTRktYAGicvRenNvjHCCKtuj6rrB36wovoeRWOeltiASqR/KvGeF0
8AQxqZI5WB3DLZgyNV+PUrS1Ps3j6TJFZJoZ6bM6MBjBZJU2yb+853nfo9T5PNYN
664fB6vf3DjgJmBLcua/2+DVifVN+WwimBg/+jN/gRjsik1Hr2ic120IQNTPWOrh
IsqtMh84yxEQNiK5s7SfK2JSB1ps2cKOSf+v69QHbU4WWra0MHRMDkWHZG7O2bYL
nMFHBlGc0DkbVWbb/rlUbsskwdIcMjzN7VbrCu4jAo7nWqa2xClu373BQarBK5SM
pdTgbiieDXdaWWOlpgf/m5K3ZGyCMOl4KM6k8AGSDikeT8NbGdBJ+6XdvQ97bNuy
N+fHVSqvzFNfke57xWAYx6FdE9P6/4lyEVTEqKhheaPL03oBTq2uVNiSHJt89796
AOfQmJ+/zaGxt+WmZFKLeYDj5RcnH9u0XbJmHe3H7vMQIb1EnHPrYKjWsPi3WxZx
3jzeSIBKoxJ+lgEndyt1nSzjmwASOKIa3sspW5VFlazgYhgWSKz9al6tGcoyluvl
zUuvZCr3OWNxB4PkqWlcGgpEbH6j2guGnHbtuwFvZ0nEDEoF1kQgrJpGptIgpl4a
Itkzwvz+VqktIeSxraNbgbr9mag3cVlb/H71XJRvkANBPxkke8dx49XDM0n+RH0b
riZCS8qlrZnwo1XiRgjqIPcjjenmH+DCuz7GfFI2caj+rzU78SfzmmW1QFsB0EPd
rhNeE06Wnu4DMLFcIe5KN4bdblzQrH3MfWKTBB3Yzl6Ery8LAXugIo8UZezuwEdc
psv9mT0CbkIeQ+HmfRito0GffyICntXNsxpAfPxgjPY8Iu6lhtA06sniaw4KGfK+
Bbgu9zHDMp9z0QW9wjMih6Xl5p2pbTY/8g3FbPrl6biofkmM8XpEUjSmlbNnRsHa
MR52CBkjJ7YqcCR9Egmo2dMzXOrkJS9byC8qlGzmJzsQQ2R9Sanck5siENBlhZMk
CkngCBgkZZIBsog5EduBCSLy6egeTSoIz7D5+6xcYGU2DxoUAnpiW0VUWyy2qhED
AL+o8XptXKrYFmf5MtQPjGCUKsBv4HBbamTxOIcnbVoM7ItY648Wuq4phg2SB8I8
ulyyyQJCO7czUebATKJAB1ktLsrCG0KJV6rAYodaGplbqgW7THO74mXGQBons4j6
ch+eEnj754WW8dTttq35D8K7ZSHc+Rwr8DvY4Y1q6KWKruC+GCsFH2Fi9LOdTGHv
1ObWvQhXv+tbx/i72BmVOA1lZwdrTPH0TBx9iGHIMYcPiXlOY5AN2byP5i6zRL5x
2A16ABnKhiaBTaUyBVoeLUeZEH5CBFOc0k/YQWwEjk9oGpIlA3CVfz763g7AAv/8
kvBjDzu8htSrm15fcwRwsimD0smU4i+lrk1yLsNWPf9GkQV4LEbvCAIh7u3/POJk
Xi7x+eWQgNYiNcsyPyLuQDlvOUq0oEskQC4wbKlQDL+9V7G6NThWN/JgfegU1ir0
aPedM7KWAyut+eM607A9pC4+1EabLso/Y2OKtjTEfJFpeACTCy5xZO5/X9mYc5Et
BHuFcEMRmair3RxBjrNaEz3SPGrP0Eyn5Dxl/LDh/f/FPVH1+DmiaPKgOv95J2wy
opsNwZWp+Fx8ZMcACyO6IX/GpcZtsLjoLJjgwJnBl13arAOVe24uVOiLPcvHkKsi
jck87jIa/E43f0q+UiUmIFxUhsYvizmhEY1pAWkq8NjuhQQLnkSEOjwUxX/twI/I
TnJ+cyGhstxCIauGnqczI/fsby+4OPcHCnGY58t7SNHqSLylmKR/d8p4FMYza0EG
N/claGIPSO+WsD8avyqkNBJcN94XKY1BvPvAwQruBHm413yVSZKoROhQzj8NNPcZ
v2mJzPW4BQxqUHVW+dYPfpfJSIQ+VTuLTmZjsMZMBvArmw+QUA6pZdTdCI7VVUBu
e8Hv5mCpw9fe+um6BV/nmCz4ShGxeIhOkaapBbYAjJm7BJCCthsTkC+vYn2KOpTu
nvojqPDNi86iL8NC7knzNdAmFsswLp8hAR6oUmtZRju6boz23T6bS8iaCHfvWHbM
QmCi2P3AEZ43fBn0MQUoY9v5E/wIjLG1Q/BnU97bpI/7zOtGc5ARfCix8Ztu//uH
dH1J4pR1AopNZDQiGl/c8FnUSoFIYmk6cyCD5ZeesKGWTGrehL3yv7p+NnaWiutZ
xFhZb27ExCjqJeTYvZlEUoQW8L6DDwgVkUK3RNbPzxEEJQTaTf/4WBrgQAYfjT6n
JX+RNhxxjy52EkLbb1GHg+djZzdApzblXIZ59nSZ6cJPhsEGFj7o2k2BlKDvBW03
qnzyQnlO1MK0Xzk6a72uZoxvqhff4WvHL1Q/BC6joe4EMKBwbjAwcYYJNEddkidG
MyIy+nInPBHW3Vdc3Ph2Plb5FwLwMFlNvVeHSpGnxkNcT/Hpw6aJABbWAYo6eavn
HJXTdPB5p0670Xt00hTeEE7i2geol+Hi7yibWVIRKW/9XRG278HDT45mR5HtXvZM
JwrE4WYKVjBB35pdHir1Z6X+dWaD8tFrUzd2gYh09HF2TnCt4JX3b0/AfzjEnT8Z
9nTe60S5A/+BaYPOLkrrwbJUAFA3IYVnGHBHVdzO2CJI8qlMCoFxWOkcY6OMpj5t
UylqAnewxLhmRyQSTU0syvlM9WF8npOyAliJhxybeDuZ56QAc0DFxMqr2+2co2nw
qnf9VRJJ54Ml+nW5uLm5UQ50r2DI4b5ydXwlaDmemTfqSUwGIcw0+t12VE4qfPMQ
wG4Sq78zlD9dVISK0ouCtIK5Y3tqKo/0A4F+cJ2qwh9oWmnlIuNhVFjNyjx0Cvg1
Je2DaVkYt652mUei7gfIT9TigEfBS9QinOQoXpTs0c6j/SxnjzXwAAeV6u2Akf3s
d/gQHhYqR9PM6CKpitCEvvE15a2jiuDgUAE3b7m6R3ytE+s4Wge6CthBcgY84vCP
jhouYI2Xsm318GlBE/99M/aJ2P1RaQLZ5IvMkKj5rIdbBFUSMFa8JUFfSYklxUB3
vBHDoJp8YlSipXyuZoEhxmZHb+XOLmIPJkaa5y5RAcPbvzDwm5udYejYwezLMNTg
2Mxk0pMU5o3/Ij/9xpcWVRy5RzBxyV3AEoXzGDa3UrhX/DVWhcT3HzRliQYGv+IE
1V7htWCx9femV8L6nNBlIfbUofFb56PcoAWhtOhS0w+4w1w3+jYJ1015sxpmwSM+
R19+aEPI12FU/H0xe5w0S9yMrrJUzbgFpfXnSX+IEA6t1yQuT1fGcM2C1kbKagU2
SLLgA3y8In0Byi1S8akKZ4MYpz0FDdrqShhKclez5+KD1PcWtk9oF2k1QYdhFKN8
uOwigETsJGVhaShMTajc433mwVNMGvy9CZvYrPme7Oi1RtT+0v2oESJCR0A3PxVt
6qhVls1ks+h+ooFC69gqO3anGZYj3YPeCv7WZzccfVo7A3MHzocczUr/z5JZzNSg
stNjyE/F2/Wh5oaF8AWZsvt0mnj3lsO5i8in3h6ZWmjKlQjk795feP8/isn80Bcz
Hk9B8EFtN62wNUIgJUi4GaYaBK1D/vSVlxdUbjf00mieF8NJUAODko3bCHpW1BEs
zIMt9vCmGsHV3fimupdM3EL0nLQadpR6turb07t/TpM9ez0Ah78UZe+YAAzPj+82
QI+5XUazS+zroUI1WtMZErAa9o7PzpMpyUh8ppqZeZACZuzCauXSykrGe+nmWp0P
k+WGa9Deh2XVDtlQDA7COd53PCxkpzGYbDfbfRBeb55qP1rikZ4F8PQpizp21b6u
/q5zgI0UsydNL8D39t4DLx5WDIs6YuL8ajEW3Tx0LcMTPFAxAId4rBQs2l74Hbm1
vTwU7Bv2rqy8Ms/E/mRC7yENmzeG6dWe0UZjtJ3KEpCAGM+MHMglmqcYFu5XPOcI
qczkNUS83/9fsMwfZ7cIa/f2sb2mpM2EqSq+Mh5ur9sOqYI8jUhT62xIwyDW/C2z
TIMM5yQSWJVsB6jLp1O02tBn+NSydzrQm7AbdljAFwWUo5AVh6XX4QgVJTvdzWwU
TaJoNht/QCZG+1wtDZGH88zIf7z63QJbB5CNoLInYrhiXJN/l8yREA9tJvxPYodu
w970PRmbfeNxmYTXpSGvS8nNFFWv6BetSHGIAfFYILPox9XKMFcUVgffc0H/xwC0
Vqacrx2ckzZY1uMSOFrbPBbzHE9Nvml1T8gQJoDu95akz1BlcAHksxZMgOVpNKfE
JmFHL2Iyvstc5AIspTYY7G+QE0+r+xWINY+wbQ/rCnTvn3VlNS2mapgrbJ0WR4dE
VfDM0naw78L8qqtbLkFH/9OZd1S3aJAiJeHyvSlrlunhjczcVh6AJrZnTI5Kdk8Y
tL9jR/vuOvgzo5cYjjYCqmtFOmsAXpJZYA/g1gFUM3UjPOysNtJ0ayodC6k4Ag6c
/hpZM5BMsNVU8qVOPNLkTePHuapo71TOFnlvNYzgi1LUkMYCZ3urGGDL1Yy0X59R
ojsb3wZHF+pS4uM9cEJPum5BwratCgwjAvBjrTI9XEXvuZ/RwOtUkpk6E7XQYGc1
dIPQIyoNvFlY9H8X2Eg/AoW5WyU4j/Nl108z2YiVITQG74LfKqi5Z2F3JrQhQx53
PJtLf5126JeRW5z3QJL0Kf4jDfGYpZsI5AlZ4cBiV4nmSLDkVyB1XKuExlsVNfBu
ZqHuzQAudFFiMRO8tWCSiiXb4OZuP01ka43xpzsr/tKWJDEVHRkYYB7tEo5pQ9bY
4c/Fki9j5/pe4GtLkORSK5EULI/r3zU9cWSic041aMDFlT8FRPBLH4B40LohI1Yi
3pEJyFjjxQcRw8u6r0EMIatqcOPnCNskxqZPLrpn0SSX2f1rR3/xCV2jU5j9o5ox
SnQ3IGdqU2t9lRfzDir4s3QU+k0Jaw7xaH/S/+WeNWYaCi1wXJZZTqrEBIWieLPS
RWYD6oWq4UKfZiMaoLZFjnxs9WwIpHxczYIitEJSTMdq668ovfyHQNtUfXcWIa9X
rRSesk+vd3/czrzxTh5IyrxWo1nAOQfxrGt9b1Gqu8O519hxCvEVM7QmYxahWQst
lUNJsDA3986w+ikpUFM67ihpQohZ5d7COlKY14q9qT1E7EQNbvagxDsZ8zqWMxWP
h/22Aiq/S9Y9/eCVZJIlMaAlckKLGLBaa/6qAj6YdW1BvpCupJ4HT8Au7yygF7Ay
AWmObIrfccSQ3FNekCtM8oZz9u+IHS5Z8XfeNg+xPkaeeVm/VnVlBL37BLGv27Ss
CETqxPUqCpYtmfxac36vpMeDBOh6oGxJa9d2WoPaNHWYDUYoyVdCbHLFBkMxsUCa
BcF65bgWH9dl2aIpGt/B22FO+kBTISKpwmHp8OXy5qfg8SOj2O31KGQMXCMNiHsN
YhpFiFr2yDB8GzKyLn/QspCDSyyyUcMj7nrhraZwQWSbfbXNOZSpDrQNext01kUi
C/qyhxXa4Hf7XMat5kDzb1Krs8dylOxw8cR8SL030kiiOnRJTZBXcDmlH6TnrGAY
cL3Kx2TmljPCq+kiH9aZrSxlCGImqvKaI+9Ny8jgDXhXamzNKvwbVIKJshh0TZ3P
Eln5JXvJ/8SCS4XAIPOXrYdGMmP4gSBcI6n2GxJtbT7zcpggHdKdbc8QRNhvLBow
jDQai7zNy0asbLqH3pbEC8bHRQfknhLTZGq7KEvLWmW/l/yX2o09GtkPFXPlbzon
YDt2UBFkDOXZ3EooU6sKpdCStGnazLgVlysvTw4rfoizkL0ov0r9anzGO1In8afM
xXdVsCPuSOCqx85/RawELrw8jQn/AWvHTX5dm6jqCn/cn05xdi/o0Ci/syt17nvh
QJ+ojic2sTh0//KlsJclR4t4c4sHUKESbMiK65FNu6vuvgnz/f0KsnYeITKuOluA
6rzJdYzZXB3uXkj2pCqYGXYLKt5pq/O7///XUgZtCnn+OLDPu3UOUjw1Ba1YP0DS
Kc5bfn9n6t+PkfsulfjrtlN2twCDVRIxqqPvnZpCqHNe2w5+fMizp07EJRXFZV+P
wb5Odf+VO1edJa79So/e4By0Tzve0yfD8Vg9DV4EKwnCBSnYkRLkgdy6sGFKJ3dw
3eY7RrxNFL+d89ARdENPcnNixR01CxS0iefVUfHQFp5yBHCqENYDWz3ANHGj5SBn
E9EAKMRu+HbRdSij96NkAtQESayfn5J7jiBQPkHNGlzdD4cJ5KLJ6mJES+oF8EBX
T/coR21LMxhWRGevq1J/I31cQi+df9qa+3iD3chkFLMG3dpaUYIcgnalueWYBTwb
UUfb+dOZ8Cw33hiIZ5NzBLTyjJBaxNS/GYsXoznM85aeKpcP75kBnWwIVWxXLKqx
r/itZxkUbnba4ocqV/dg04usN3c5S8LPpJi/9lsAWMXt/dEvj4+YqaKqw5mQqCvh
3snOCKRE5YKxnpLDxX3rQwVI2XnKZNReCTMZESh62Lqt7sg5F3joCM6uPzgU+jY3
8rPzMjzNy+B4jgRl3DzkVaWP9xA362GxEOQuOJYPB5jglRBOE6jau+L8hClIucj0
PxmCUaG3amcc/ewel+J8G9dKGFHh0ksbPkPT6tz9KnUX4MUToC63gscOj7zI56qV
JmP3BEyUZKd60HLbJE0d6SmT+j+JHk8XxzOHIMRo0c5Py+pCd3nWX3Se3M0+mFLE
15zGyoKB31vkMMTjNm6q4sfF1TNf914bNDmJCn4+E3F/21ILodNAL1NsZ8u+3Gmp
Rl5M+OnUIVdJfwJ+HO7RtRYYDk5QWE/qRQyFA0TrwR7p7FgYN/Pv9pWRtsBRopYK
m2wp9BOA74kAEfvdweHYAk9PrNdTK9SkcdesHjdoANbxcjcWLto7q9A+S/oKJ6i6
A9gGdD9yG/htxuijhCUKlTi/f/8ow12NWB6ifMuSh1TO1nOrpxedNqsmTJijjW5H
LaErEgFFM6+RGuQIz2bMWIARG+rfOCM6OApBmxNLsmMcyRnkytEGFs9IZkNxdTRw
ZoV2G91/tnYY05FxuCRrgT2c7YhbkKn5Eo/WU9ryKqrnCk7n9GT8mtVFNj1dqNsK
kJZ5TkiZ7ZCEQ1fI7rgzhjzK1ai12reR9mHoWN5hiiUpQ0NWhQtUxbWqy3hR4WhE
m4YaG58bTIhsBOVs165Um+VQHp9XuTIORnDdsXclQILQabtfE8hfGLOtc/8KnvZV
BQJh7MAQX9gbU8kZ/FI7WGl78SRIHRB9w429cipQF2a4mf9nBIWLYPfJYPGwhC37
dR4HcqLQV87LUUzO8rtQrlO14zrD/qHYcWgv/zYn7205uoWlaa7Hdu07CFdLBPDP
/WYLutvw1AXNMJ+AARLP0XfV3/BlrtXgjZm1ckBLGay081Ikq9qJS3WHZGgHZeh+
RB+6hf1s8kBxVSeGDrhE7b/solSj1oBa7ikH9dziYFv2IHqHGZpOmdP0csb55HZh
h90QJu0UbTmx8AyJVC1KJSh5sl5dfoiEwqY1tGKvWq8VCEvh/m0qvkOch0x4eToD
nnYmJBU+EbeSkK9NUUcrjyz78ySLCOHIHEBzgKstxDiqSri7zHN0oWeMdai/msrv
DpjhV/y3qSLouimsEs4c7w+TqjaOFzE4SyuYljDjGQx9Lsh69bF7u16qGdI17jGv
WGGM5hoanmDpyVBP40ZCzdLaaYvhx3N2M8sjkc8VX9QEIZc7yozJOPHd3SdumQz2
Wl2TGioChXxzJSbpBypq1N+w+diB8yYcD9f6kLmoYQFVMnC7Z8CEcuOQQQ3t0GFg
BxltMIxvnhz3CSpZKUJL7LmGICo0QXmXw12FAeM4GUXDNmr2DYQEPJpou2+F5ul0
3zbuVwHxNmH4s3pcOqAPfFL0GbbgykLHe9uNBxLKGM0KKf2aTKG9r4GPL4z38HVW
iJ8/p1EUWTLnWWXtfKY0qwCZvzHIQ5Pa6d6mkrziby+V+LMCDKtug3THurp9EAZ4
7ItsfncrJslljvcXftm62kpRzKIjYdjQk8q1okssvow+Adz8AE1pjX2bYvba48Oh
U6XxaHeJYwuSAZzy6uwdqq3rtwlxEVjzlzY5gMoSBmO/EG4svYGw3y/yzyl6kNiy
sIIiKA7D+3sGdwwEgWhSEvJW6naCnRD+QgCbFG0ZbSiHcaR7ernUMslOG83+WdPT
LbeL0zwXyHKTOsZI3JxlBzUct4S/vynUW8IVb+j0jqlScs4oXGpwOoxZGd0BMwSr
w4gg/Ow6TIDomFE4jFkDhCNzF4OwNqqyiGW2qQ9z/u3YO5GWE+MhH3eZ+h+rG8Vx
niBr76A79G8R+3yAweFqvBzD85Ei3ifijWXiAH4UIYkOblT1jFn5nUJDx2cS9z1P
i3T9tngHNSHH3amRP2wwNDSyNUFrhqyg40229rSzt55Pr84s1OmhhJo+fIFrBGNX
D1j94KQKkmzfcN6q36eYQiEY+XEbz25kVHzn1jluBOa/RrdzobVkfqSZqFFGuLoE
j5OxmSRZ87ZBFNEI8/zul1eIU3kWg9wwJ/5yLv5siYQzX37Mo7bqmkOu1B6du87m
7vpgUm1uTFjbUTfpXL2QtJplrEkxGBjjxAitugJVS8WQ3Kw4Fjh923THQBLCqGSk
FJf2WoRGHJ2mkcFbZsNgiS3PySrN/zuJ9FrdzzCPtLu/p+LRROMevU50LDq/xmG9
viXNP382MS5gtL1TBQxxFeYFE9Y6B0jz1i7po9HPCWaM6zjYEBzxBLZST0chsDu9
YS+QQK88xauZS7u2GCQ3X4acdf0aO7qeo10i/2yN9uh6WaXW1AY33szGqeu4/Nvw
VJ912/3uUWxPH9E0ZK6v7n7am72f7EyJKqqPJgSefZvl4Wry+zlAyRYq3MkCUlyV
izzSgqf6OL1DQwHh95TG1+hjk3AzH6U+UfHpaffikdYfygcBNzneKqXgeMsb3CYR
ZQzCSBggWNSHOyAAp0CK5V+/i+Z8venxP0HSMqfVUgg2AUd/lHwQ1IZ47jladMA7
4Yarfre4y/GLXZ9dbcr59i8j0/3L+9cpRkrB7JAK6DCVchyTvfjpVdwMnskHpXgt
OQ0q+0MdT8ZfkEVkclIWKcPvs/ZnUV/kf2wOGcnsdM/n/GewMEvOmqp8gDz7Hktw
bbqBCLUfeZCWUvXWoOl3OcXYS43uHSlu9ZOC2V2yepSX8cYiPvUqG1Lsx+g3TNpv
UeTRpCDSqa1JeCQzvslChR5KOldLX9+wrL4pLsUhRPub5vEIUzjkJAY6Ptq0Ich/
IdNwujOjtm4LaBJBxtsH4nsleM9pXEjmcSJp+DkFbFmDydo9HlO61yRlC1LSplgX
j9HVd+GorDwStZFT5OpJEq7Tfe25SvKMvnuRIB4ykfaqs3a+lXIGPx0PqYVwtMw2
ZjTtdOX+UmVst7/TBAnhorcfR3X3Ck14OiLQXHdXMI2EVRJ7vE8XmegR3jyBwDrh
Fnoh2CbkrF8eCJhj1DaWctJbE0wNL9iJ/7+BeWK02ACedVAh3KQ+vPKsoxRHmthE
0scfyXILuEtyUjRI8Ctgv95PHMEwVmL25SEp9nwq33DRwMODbIIBh+Zm/HuVUZjd
VclyMfP4mp7VfPBfa7G4y587Z26uGxoJpGWzeFSXWG5sXuKdSogrRriPyojRvZmf
aVKRmOxP+XaGzZ6puBp6aBRfAzPzM3znMLCpUyTUAZ2w2f+1+HJ9SLIpQzUmHznW
sxKlPVrPA2+YNzaZMEVAvIviiwasjYSqjhIuG6+u26ukttgO+DOBMWrh8417eNvx
x+BlpZYkia3nAc0pTUPpAXT3DH1qU3rlHMCTj05Lw4cqUguO5jOgMptBIqCVpEui
A3gWLBO+6uDqaq3Dbjkb3u3xWpEgdGXTK/Fr1uPwni1CbXNcX1t+R6VPuHRg/Lvb
kRRAGx0pny8V9gz6Q8LjeKY74UuFvCFxLJEcoy+glUxbqEaO0X8InR0vfz9XLvXe
hM2kkxwPqHxOKGftsRaSe3CI4ZjV1pLAWHw70r1h1KqcMx6F6/IoqDX1aNEIin+i
y+OgFACWrExWa4joJ+Sg5Eamf2wySJm++DYAUjRrDbJM/jhrNqaISn1CXmOxlQmW
QZGyU8Lw/ouQAs+DnKbfwrORY2nOfXwxBaB1FyI04OA1mG2HCiPhZxtaexG1Ndzs
GBMJju2B6R9nHC5kqvGjcgsmYjolmXrNBMVEx2X4PT4hP2A0Q0hB99t+1dIqNlCc
xgVzzxmzdutqvvfJDR9e4tRT0OtXdfHMqNLSRu8y/GPJrkdhgHMJlWIfO4rMPg5o
NiySciPFoyonY3SW8UFjF4OcdWgwOHubFTr9pk8cQIexIvR1uZ5pVIAl+a0WQ6IE
mzTyiEDlk6I5m1v8sPaN2ZzWpqoUBbz4hXjuIQ2wQeIvlfgjkoIHGodU45HO3Eq1
Mm3gMBeAsvv5CE+FTuHlwp7jG0uDxIB3rUGrNREYDsUdVOF8cL1+9l1DwwU6o/s6
ENXQ+gT5gc/KKh/MT9OCO8JeEBP3hGU8hbn6M0GftOLmCjgZ186Ko/PG/MoJw5ni
bAtLVSRJ8IXj9Oj2Jz/Bt6spB3XFw36oT1cRHhiAi2Xt/X41uNDgdMuPmWOqQI0h
EBR80zNbzHxoG0L9DAb2RTFpgUDp/w+OmQIVD5dsx4i65Qzz/LKGvaO+iJ093r3I
+B+6t6EBWz+XR7MvwZ4URQ72keSYHTgqKhAkHpYGnvN78tkw9c1lluIi3Waw3V9n
0DOlN4xDVSoFW9mLgToU8tR/NiT3xkkcwqKRd9kO9oVF38vB8bIHfV3XN5BFPXEO
Lb/EWn7qYQJpzqHCT4LP+cAlgXgfTHX/casWkoTeuXVoNEAGXFuoLvvKc3XEnnpS
aIoaA56jq/IPo7HIiiTRbOcYPas0mxfnO+1MCtdcuBscorC/eJHsiaXkeMkgswSE
aMjrSuEgaBJqvpJhtQOrHCIXAf1BZsfifhig/iZYaA/CCR/yiH1So7j9mH7kE3aL
/Lr9DuSytjG2yev1PgJj0hHXerSqCYW58c85Xer3a5IOrmC+PGEH+BqJKzMksyA3
y/M3ZBtpHSW9iQoCEZABCBxhUcUSxxgYFyevlcGugD1utQJeIQB7Xc4JrCidPpdj
n3WPkQIA5rDLqaD08rlU+vV8evxOJ4runUkGgEoXG4gz8HboxsEef442MGxrzKMl
SwN/BD1TXkN5uRr9r73HUn+BYMitXBlJ67+xLC/ekJ7adEzx9yhB3agmzwBEWATU
y0JVf4F4yMjknWZQhBMB/3puzfcTqMftg/9yKcxB7PN6P5uRnXHLeFQCLuHdFDty
98D5SI9cKc+tZdH4G72bL/jPazVY0932RgEplFCg6Vf+5I0SStqBF69CWT2NzsdO
Gl1Cn+w27dqwAYMv0qAz7JslowBONbbZ8HiMFWReXnO3KOLqUWj6r+5Lld2Rhk4W
ik35k/tcc3MNhNGVUy/VX0njeruFFNq3xlMmUIwW7RBB3Pk1g26tIOKmBC1GC3Rt
fPwJNOmi3MpXcmGWPCVataR8DZ0KpK8COUTir+sHtOBXhWcKwAJFoQ86/UJev1E3
0mVhUdKC2sOtL1+eXciEHtcAML6RRJp/qqp2zEoPe1UJ1eK8SdA3mP+Kse/T7Uh5
s++5fSrC/hyNaSYWWjKoXxWwt4xzypEwv7U123Ot8deqSVHXV7E9WN66gg2ftGur
ui9uzN3Z650kM5MBzxwBbu1d7t+jk5ork68+EtGg8ONUIjnSienEAnmMMavP5qTc
ErqwM1sgUziZdsQMD9euV5vrQ5MReAqLVgNFU09dETAxhVFy2rx6xDwXVhVjJLMA
f5QxDOebfWpIjis5sm9HVByG5un7ykVGXuyepKd5siJr4abQAtQLfa30wTmrccC+
RqzNzY4iuS0k9bVFscmVAu6JaVF7C6qN8wy7Qhq7ttwEm2ZoZcpjKaYyvtHVpxhr
KLzrMK3y7aHoESjfdDsCnqkCjbHXoas22X4iCVjOMyPrDtFN4vG65pvDjU/YaPKw
yfTMRt+Mt5EYDZQETwPOsoTfJNaxRbkGJ96GOzXkjuMYQroQxkl3WZG3w4uslg64
0nM2ou9EH2V8o7M4JNW+JnE+NDhXVY4LeqzwsQrWLunQfmymqsZ4qrN0aP1AnCyI
sqBtLVRaH33XUS1oGvVtHs1W1brDJfyfBnFXenz2v/hDnOIlhTdbb7/ZWEu3Cfp0
6vmKanMbCOJL7gFfzY9KCrMHDYECHOTSWaK6QlHUz8aBQbIU/79LkrTNHBZ6IO0z
2EvDy5RgEotEpdCTiKxT69WzBNob5icSHHUYQpzWn52WaIDZn7CmqLHhEHW3XwMX
xUIvB4WeYuk7LL91P3Htobz5yknYQh2Opp2YK++kZ5N+mfFZnqvN7fhzfiD5ge5F
65wVfchaxl7PHp0HgAXMBMQehUI1DHqd8QWUUHJrDiUWPhSE1NZA//NbAicaxMId
F9NH3g5fi2L2p7JVNQluJS1p7oYgoVbArAvuGcuR5S6UDWSyL31VcaRn7ehfLufg
XXeGTtXqAYXqmJGltbdY+Sc/QVROJ9AaEBFAq8f9CjpOVvwHFmvQjlKlUEVZnWM0
zyiQR7JaF7CFvtmOvzozlhcctF5uPXKPrHpb31ZoVr2t5PurRDwRMsDxCt7qnDmB
BLEHKBsgnyORniIFwnRoxvjGrFHWQzasUbuSdWhgIVDrFdsyg0kqQ71dfVozDe7b
Ycpi31urnwUJvGStVZvkmA5Uf8/episeK8WrPeIRIHeU9eaL+GOFvXy5PN9ZIKqe
UExTwELR5O5hHzHN0EqrjK1RNmnLkGVmDcf4vRLkT6dJE0rkxae3dgPdR+JRxf+V
oxLII1IettXsv4igKe9dziFvKarWR2wMZSgX/ai2djmZFLqHkSEuxw0EF2mnOPmn
pxXFUI1UvuGXSToSN+whe3nHSZ2W3LjPy8bVh0qcfNl2lC2I+NUdMh+1K/GE8bFM
gs2u1IfJicA884AMYhwt0H6xQvXiMd/Xu+secBLwk4iAOjrjdD1VBMB/TVE9mMcs
MbgVR5OZt+FnYOFQXWDJ6yojYz/vhrNPvIs9N3BP6o8Io0uAQLnTi1Ghhe4ZTl4A
MLl5fQ8UxjvlehXHysZk5x8rkc5GQN6xDYAtKZq5InwJI6J8IP0rPzP/aA+g/Hqm
wP4wyveFxx05NAUWTIHQc9PTHNBqKbuqcmUdlJffr2AdB2zVqm9U4tnmBdjRXlYi
K/DPfEO59F5imgApX/40lJZpPC65eh52b59lDXtEFQrC0evR6FviqZ9MBOvHQaKM
/WM2z46CzgS5e77pC1H9WRZ2iRr19300+HjyBcXfMxombd7o9p3yQDH8jxYHu3Fe
kXF/i/XcVoD2Q4nldy1H+MZqfZqQGI5Bz2xV0XUhwrCrscJJJW/UufaGQER+0992
BxsWHKqG+l6TkbkFutzK2Bhbt8GgKy1HMzqqfAPMCZ1gHj9wmtbYcvFpb5vjjSYm
EbL/sO56Do02CFaSSuItx93DLN8YVlVSuKSVo9e+AhjR07j8R4SGnlp0vHDzx3vX
2x5m8zFtWWCk+BjodGrmgP34xCvuGlV/XAOCcBoAXLSP3RYQjGpEh2Au0FlmDJCN
tOZ5yP3H9irjJqfPRkLZha5wKco+c2F8BrExvQMVpEmr1pQC6M5Vqp90zHMshwwj
MViCKFrZZchhsK1JIbWJg8F0ISQbZwkdG8RqQuNzcFenSzzQyE4aICHzt0jUKjEt
hxnaYm48VJuTIh+BifBVhIi0xZTB6Ia3vIrDTDwgM7x2Y5oYMi4a8Fs75i4DFoso
ibycHRxMU+Ph0Oc8OaCcjVtX7qoismjj+hRjxb0bIYB6Xgj3E01bVGBxsXtRxfQm
Q2p19Ituv1XT7l5NYpYETMh0I7Xzy9o7JaTzfLs+/fx9OPhuvgeW1w4YoI1ju7g9
tSEiN6dOb+sUtB5U1tqfqdRnj0P2dEU0wZ1224EzTh4yommxE8Tyh/L66VajFG/s
EdsHSarOf1JF0GRJ9HuwRIYmhB6jB9uq88CT2SfRvlbic0tQvcViowRdsj7aGem5
ma4FVd3borOeVcr0U4UuDykgyRWezmhk/Ek4hO0Po6nT/fz5lz7+US2nxgIZrsp5
6hVwN3iwYpTD8FgJHH6YOzVu76qDBnoQfHEfyhnijQXWzJ5+wLRZbTnpGqzwxjoV
XcoQPKPYBBddkscRDDiruJZCxSKYUOjcm5n/w7/CCCHZJ4tirEE3INsmJL22B++2
03fM8UmFHS91qF+Tyg8Co4v6KCKWUbJvw0MJq6yaf+7rZjGr7JBAP9bNRlbXyHoP
So7Nxl9z93HHNNysfAs/Isbmapm0b9aGMgo4X/9zMb0Jk9ai+FQHQAMTp+DljOiC
KRhtAUZRBFwk/Wy7xK6z4gdBEhwPZ0raIFc/8XPFJyBkoMP3G83YFp1RDDlDobey
CGCoMZIVCtmrSVzmEHt9h1oD1Yk4V+E3hfhoYx4QYuyDQ3h7mmNmHnr6t6l2wQLf
yH06LGioMgKldjcZMnm33T+8u8Yob9gl47T2dltMbSbnGs5FqRSH0J2S63k8hqFZ
TkcnlkxUOlhBJH1fHLG0qbBAYfWaBe7qi+jdcYnwPLDmPB9tW93O28Xd9iS6+g3d
Ttsd3+WD4M9OoiCN6FatLpCpShsFz6Whb0A6QBlqgpYL4ZdoWYPHZdMyBEHmnDfU
Sj2//9vHADlY3vDY4ruGca1dn0j3iYha8ugpAkEQL/SLaqiaRhzPa7tgEm4qiQlG
3wo39TSDjFh+2cm+Ch1KfhLnUxhjguC9jsmcYeo74mQApgxta57U3urDrhD+F2AZ
BZBDl0Pr9FWmAdhQgoGRMzwLbcazVm/mAVHd8OVI4aj+D3b85Im4vcFPQt3PbX5e
IPJzuN6CJUpmCk+6NyYHwEuGJDeiaUxn2X+Kx/MyzALYfq75gZ79Q8a2Na9bYrBF
4FjpjWjZift6NSkLp4f+N7mB0PT6OSbfeoDsEaCYFVh1Xnz/LjaR9OwD/9OJmFcx
fdzg0NKXWEA/08DgX6hYuNfSYtt6s3I2gdeG1m4eJDahg6SQYm4ps9XT9wyneriu
8+GJrHFrIk6BMg/9c73mUvwlqANBR9mO3QBAJePs9LIr+8mJbDD41eLB5s29kWYW
MEWPPbax2uMLJAehs6fbEz15JcmyNquXPY1HVIa6xRje3QgKJbnOPLdLgLHLGIsQ
UEzKJYXKS41/rqH/X/zVFsQ+YByD2H+MEbgxB3t1jytwvGD2a4fkwiK5DRaZZxef
VMAV5wI53SX0dDTnbNYihNTQ4+qf2wGqcgSUUNK5dWPNZGd2phyMfqPFjqk70PRu
9NTE/nbThL3eh2ilZUoxzHjubGKwCExnqAo7z7z2ULHjyoUJ7VdA+ZjWaLQBmNdk
njMXvZPqtvyRR3IiOfuLDErD8MTZfYG92P3LPAi0V1q4H6eD0/Xblg7XySQ80N8V
AwRTZTkXit+iAHKMKLmzrVVtkxbnL3LbA1PIhXGLxmtQhQv7nfzKXJ4yVBmaNKtE
dK8SukuJ75DRkAfB9bYLPBPSNjjpxGUnNjrDPVLwdtf7J0y67/e4bpczNJwl8E5W
Y3+ia00BozhFk3cAm6skn7C9STbJmpdMjhzD62E42SFYbeD7oi/Q3Dpj4WGYKRQi
Z57xcAunogN+F49UN9CSWwrndEFxFffTTzrMS/x9Z9pxTmCMkl2v3FXuW2nXu68A
aodGtTGc8rBwpyDdcQq+MaupFUueDH9kDiink6dKb3jz0diVEXaGtCA65DrcOC+f
MIaqfhvlh4hoe2Hep20EzQZKcQgw3UGgPx+Kull67156mXxb9//1pYa85xvpDyjt
WPyKyUZtuoMMjvHDQFAVo+JaRRIVWPPM/8HZVP6Sz8uHo+Qexyc5s6JdBhlrb3Pt
lZQAkGDn+u1P0GkiCiAw8ErVks4O08166mfvi+QRK+0LqCNiyG9sB1Icheb7qVV0
DwcqxpHspK3Sp3n3TSHc4X+0cjvBXulFbGvWokBkX6LcBATRAWNiHCzrslWEKMH+
aIhYg+FOGTjRUGbntVPo1CUDJLuDcqo1mus22oB/UljlmmHV45IFAvjCGJjwjWjR
EbU846LY8b4IC+qFmnuLE/AKqDzSs1VpvMrIwBylmSdRLl8pWrTtuescWNvm8oIX
mIvh2ZTXPLzvB9Lsoo/hKtWtJHnszeXa9l7jojBARv2Vb3hmsOuafpEa5eYAXXoX
Yw+DzEbpNcIoRoWBp1hWWwd8XjuKlBCA2bx0r453jSvyEePvYY+4XIhQ++4EurOt
PMIH7OTQq4I6a1CtVsFt9KD1/EqFULGsANC3qhlPQ0yAOfn4qwlXaYUYOwszR9CK
iRDcGxqbPgz5bAp7ysaFLv6MWTOjqTwbg23yxaCTJ3EqF9hI72I0MNl9M2szyA1l
+5bp7CZuZ8UFTiuXzWHKeGQhEPidH9SxbHpj8Oir9QM2p1Ktw3f+FdNVWzgYdXYc
uWnUmDBbUCl+liFPrcU3zXJeePedwSsQta1ixsRumkU2MRDaKeD7gfBYXCv4TT3s
93Tu8aJuuW5gbr7722+3wPxBjEVBp8C9xd6bKFt78SnYlEqGXfmrfilK8GPsBEGC
XdKfea94UcXfCkpuXnA8CPvJVTnii7re9GY7CQm2CWMHagk6kQ+GHHOE62qBPQrQ
Kia4IBsq5ECizyyo8XGCdYZFlynHmn+dUzxsRrMwL/7vD0EWFYZbTa3iC210eKBB
/Xq/NI1nVsXHN5yjEDa+1USdonORprGc0rlwOYmafoUExazBcxNANWgLj5Wlb5/t
nCSfiree/79NHa6tqWJEwOtgF9Y2aldSek4PIWag1adAbZxEWE++Pccdq6sCXWKx
BvxJXv0/lwDwwqVgJCU5bKI5n48NQDXNA3DwIQjY+CPfP12B8D2iLp0VBV8231O8
oZESSs2QpwSvPDugYA0lSZuQjtljw2aJue9gO80nb4+Nl4pUlVdO2vD23qMVPOn2
gW6MBZSqo2WZXHcR91Hrmtn3gFoig8ttE5ZXm8C8oMU1EGQ1uAND1mt4AGVdon5H
FXDOEAndHhcG1x5IrKVxUgFyfxC0V7EjwN2GT1qnE9kVv6+RkTcCn2i1Y4JXR6GH
GB3jSZQPLxpYc5WsHdS1Qb2LrxrWGrDdZcfe8Ja2ew3k3oMLyNaHEfgJ9xN1tqAT
nJxV3gXsnd3tcBxlsz+UInWhMMzMq+HQpmv84/p7tl+87GuSVWsLUaKc0cOkQtrL
lnwa3uYV7WaCYZcCuPl4lXujtVTOojqs+s1iR8gNEI2ftsmsDgiA4a5EVCCtTCo7
H3YqYyLwLCkx6MYcsChm83byUnoShe3f3mq/eCaSwiXuQEIuVb0v8YKHFitmLAJ0
I1781FPDu+aakKOzXbPhhQnUGj0GbKhDEe2Ekb8owQI+kTt9VPW1anu7AaxCnjXn
YcC72F5qPjucGq4Fhn6nge98ASUHKiZh99L0Qgu+g/nV+jFF6z+2xkqIfREdBRoR
qZpX5oIAg9W4ePO+/hpTTFV1FzCLF029L9KKdSA7h+4Uj4igjH2G+ruCz8FuICXX
uXZhYKaDYK/SyPDs6kD6XO6PXTSGveTdcGUixYYeZ8EMzH2cf2v9EuOPNW8ZeFDy
o6/SeaTRfoQBngYwBDtgwwbRZl/xldNpGsn2Q/Aiv/ZC8T3h9AjrFYwQnbjzzD57
0z8qokQjTm1RETd3DkkU/TGikK7TQhLWkez2KynQFNe/NlJEAxShSTOHU3ol3kU/
2kxlEKiDy+/cWHeDUKb2y2Wml5Jtz/DuQ0Iw4colW6fMZByOxrXjP1VoIcS5ef0T
qEihluYTkj/ajk5B14rYOyBHDAvFU18vJbu4efrwzFUYdzNRElO+vlKQO3nsh7/N
oYg+hagGKrp1uOPWBk3kmVDwvv3lSbiVBbNfWBkRMQYyf7xnskeSPCRUeXg32Y/L
4rTT/pJIgJfIG6SEiz1M4f0Rc51SdBZ7Do8oo+bewzs36vXuRfcIf1AMK2tCHBDQ
mX65IdQ0poSyeSY7bOfR52FHcnPG9v6HLeIn7Fss0E+0V0oki37PeX6p5zhBpMUJ
ZP6dVJD+XyRSAuPIROoYx8HbiQHj7acN3d9Q9jwlSnMQGfAwZ8NXZr4hgjfgcocO
gL/9H2qIE8i58ps5yn/Kbs8oJDbkQQ6fLlvWOoCzP/urp12eeaVyxKqclfftFa72
og+YBybY2D5T14tSVq5BUsIa3pQ/di4v1ucH8enOVALtGsqc0BDLvVQU7Akbycjf
r8XyaJX3G53P+R/6EM32E8rPpzvZVlYsBahiqZ+7vDWO5x531qw+c0XFd4EbjX93
zlBIwKMAvoboHqjbPUsolm7yWv52iG7jSb9km46ZpH1E+TRsA1gd+FQGcdoCm2Do
/5OXdED9ruQsJtB16LP6b8YJsw6UXyMG1tevUhQ8M7gc610UdFax6TPfo//2qCgJ
tUOZf6st++Ie1HbK+VY0Yp7rOXKkwHCN6rw+1iKDvcADd4/MVFMprKFn9+yQolDN
g88G6JdLLCaAf4+n+Gt30md5rl3dYF4bhLwEHH5m5o+dVoV6aBSUeTk8CdZ40yjv
rdGmlcyNQHnowDmDCrpr7SLuK/iTLZB+KexEJrN+/g4380fFjAW5HM4nO4JuQQNL
ibujyJvrfoG82uEzRp5MqmErxJiGXRgiwuhVaPggPOthvEl3DKfPmC7gdU1zbitW
httDnJ29Lqd3Ezk/Yk944xtKkDKGlIHp9BIFDFkYPkgj+GqDr7f7/7q0xBEQT17R
T6a4hsLtCwGiuzsziMgMrR+w0wXV3PeKaKZrLvFXy4s5YG6gRGY4QI3JQoJwXuKk
DHcgHEr65n0cnVx5VSksOj6zJB7uBgmoehm9+6++l+p71OB5BWlRk8wNuFri69Hd
jTusRb/LKkH4CUxouTsF0AK3/zGEzTleLh+zJ8VM+jdt8bl5qwu5r0OOXak/xoRa
LfeD1X0mRObxOz14FjTFJC7qYYEjC65/nxeWU7UON4LkbSoF2Sr/BRVk3MLqHq/E
YrdjWD/CGWcBFlZnEi34BaazJwLG8WCw3ZGCgIPrEtsl46SqtxxYGw35yAqirjWy
ESGwlVkWvUiHZlJj7f9aBMvsyJsEgyHRDKN5M/Gw7ApYXw3BFWFtqP26Lw9KSUOx
HmSjOM3D3NLLS8q3iMgE4Xmy7w3Qbi219D0zHhKlpX5NsxxHSP2Ip6x9Ea8LOyJo
TXCTd/+NQ5zRYUfzm44rNO6jrk4pyFxECr4PzyC0dh4Udxub5Dg2MJ62PlCx9ze3
is2CSQTgUuqZqs6GOUToay3wxIWD8BOHhO4McdZsWc+71t0/ZbwPuy5HrGdR8C6u
00C7tEwzbRFJw1xBq4+r/OukTBCScpu9wKQ6p9U3ZfU92ZKIRyeqaXHIVfOeIpFK
SYALUbi3pCMoQC4ujmtel9Cn0lf9okC5U03tSXvFOTG7UqgnqGOy49f/JXqTl3+q
EQv+pwnDA3fiG0p+7u38QwgXy+BPCi/LnC1lMTivrEpUaQ7Z1ELTSESt8+DxkLs2
E325z5WAj8ADDJZRle+u6y0t6qsyleABfItaUYgU4AJ6FdtfQ4q9c0HGqvHNz+ze
sRa7RkBmSxiOaHDJalDD9Q221ShXBusmQTw8yC59epEl9n8gk9E87ww0er7nZbWm
Sc9P2QaBc7cYV3ofcr3sgjC83lpSa6J0gAc0eMigI8AzqE1frt1TFS5lamyZ78/q
7fdvw+LK0jT+ss6UXSSOz3MCXT9vae57KK8LMWi5XvtUQDfPr0qI1aWKKsRGqRwZ
0cN/fzyrgK5+XtZZmgwcH/nwf4HAXy1i9S9rLc+Z6+Q4/MwQ0iB9end1wQgJO6dp
IDwRIcehOqFiM/9YeHawGvNl9BZpu7CZ4XYkUml2YTERrj365uV4ej+pu2ajpYSz
2z/LZoOTVA1Jvafxd+LDMwXmAJum5fAsAeAJsBPWFOQ3jHO5v9UnPKImYqIBcZS8
Xpow2RXV4xUouS4xhJwMLlBGz4ERdHOEyYXWaCX4vly/39tVClvViMXC1Jb2mkAq
cWQC9jMdSYGNLoq6Clrdq/rq4vfas/JDGGbp7rVKcI+eKsCM69qS5Xd7FKQHFAqK
7ZoUJJmoF4zkAcmDRyssgesPsoDy3/W5cPLS6wAkoYkw3IufPDvlQ0J4Tt7tvH65
O+ucwkbKbCFQZOctEcBXvlaConOAwLFt5UmAfQhCFslOahQUq8vEkHv5FpdFSkBY
9H0nQgBrna6bt8ypqF5LowIEiv/gvZNbD5EVs9cB+ZK6QqiML/jzbhqYKGHOL6UV
QVwlIPaWzX1FF+gMeoCLJMEbD4Gss/3hBW0ZjCz0nS3FYLk3H6n9gqzsGslNb985
t0O+E26CylvpfwJNlyUO6E2+pyZ4B+aFDw9O4hL5dUiF3f8BrTY+O6M9Jc/lUe/5
tmzpNw3HYp8SjvnxlHZiQ4fqvQO2JQD2Q5lkoXcfT72O2oHCbYF1h4jo1ygqEoTu
KT4H3hXpC9PmtFrhulYi8FZnQSACuv0bHUmxGrcboFM2tOLy2M8dz8WDDc1sAWhH
jeUxys/rw9XLaYdgO8XGhi+l50WpOOzm+0DO5RN/DeFVWdXwW4E62k9TDYCw171D
++pq3G1Qf5YNP5RXOLL6Et4t4TpXaiILmhdP+QlkXejyMLq6YXVqZn2MSOdqm6ru
HMmzD6V6wjBGQmVEztoZbveXdsZEn5BChve/oHbzbo18chRu0Cbwc6kwNISc165D
SMKZ5J5NmdHXZWQ6OC/6HSkHgnlIDi0pxR5EPTDPcn++NEInTp6rLve0jSiPKdza
1uzE5dqghK7NmMXK50PsFKhCjmj2gwHXXVQl+h5utFFDgWxlk+oEBfN50PIZmcfq
QHgcPAMrVnYHgz2l4JnydQD3uQnPk/wZJusmvU+1m1Qr9pVQbR99Jlv3MPyBlxOS
YtAm6Lxli2SEDOVA9KJ+1ow6ZxtjKjS40yWGJ0nr8vcbWcbdfoE8/+Q3uqNDmD5w
hkClyY4/lXZ0+0LPqvpp9+g1Bn9++bESN9I4dxyCU/a2dXSB0qsswe2E/oxbBTez
bS1fe5mxlPPTrgP2yc/HJY9gnUn+u4BPZrAdb1UbSLeetdyImPV3lgWrLmXR4OOF
DHR84c9RUJT/kkjDGSCdT4Fyl1KogBbVT7p2zryKsnBu1/x9kLZppqM4/yvvWOMQ
IYj0y4kbz6OsUEZz0+H7GOAH3IiHlPukCrr2UTX6D7tP/WooGvde9ldFt2kCPruE
OjZaOB2SHPhrqexzj32n7u4+K5Vs/I4bDTztYzdzTfKj9uhEB9/goFpmtlOdKpYA
xENI6Xbq/k6b8KfpvM+6CRV/n5c0lnc/eo8C9WbLbt5Mx3YZmyaN2rjz0YiMQLHt
DqpVDiP83l/5WN1E9jP7eArUmLZpA3O4xMzavRTtFFGUHTaeKuGWQ1RHX9X01p3+
yq9c+2UFIeoUhnkFQybOyKW/MRAFm/0DRmyCFrXVZWh9LXd9pT//BiRuRSygfzn4
zFrTAUdIA39awjzgKl6PAffPvYtRcp241q/kWKJyN8/FrauDzMxagD6HfTBFLneJ
cIKl9AtNEdpj6BRejU55gnJgkv0UWmhDxl/IvFwXNpXWeCn9NE2xvp5i5XYaQnrq
qLnYbuNJSNGwFDMcxQmW+0Gp/lg+oJCp7I1tDh+MTF+g7aiM+Wm8JUJb3AdcRkcB
fjrQQDmsh3Q/p+eSejhsyAQyXXoq2Qjvd2Ota2A+K3zSJ5kNBTk++zwYXmNIAwsL
x330qWt6KyyCUaOjE9R4TyW35CmlmZZINt6s12NW/9tKvaxiF9XQzg4RoW+mtlZ1
8dxNk/USTdXismETS/ygj+e3n+dgngqbWi1l8V9NY6AcK1QQjZa4FZj2oCHknUAL
egylkILv1IwufmbXsEwKmXjfI5jdfNRjUKmdRwWR3voUaGpbus6P7t4ozUzTbzKw
yZ7ndDAJ+nR/+AG5/DzB4ObbBL5WSoB/TqK44Q/u/LujFTYMmxb0Jc6pGf9448nS
y3btzG2JHEsvypd7g5/a9oBCLLFAIL3aVWGVWuwWrQoGjOV77LkIkV4I40GnceWx
MLUcxkXo3JpcblJXAdquk6njghqTnIkbd40LYLmhgJIrzJRyYBu50ilB0SIQEkRw
QRJ1so7LEgJWSZkfgp6nj8fTLgGfLFce3hJeGDfFQ2r10dCjpy+Zw4Ay/8S/0FbH
FHsMqdaxWpz7dQiD9I7MC73vEYUD4EOPYtcEQZGS7whGtL/qsen2156croTVDBlJ
Bbz8nSYfL6uKDpuZDq3LXAXB71ejxoF5c2bUKv9rCH/o+OUxuE+skpGjeJdXmguy
SYurn294J/XX3gbJ5Vn020jYki/XjGgCTP6s5Hmba2zz13aTlanTNGUkgp208rnk
EhLMaZakLQ3F3UGa4AnvTx4NmNDD0BvxcHfC3MoAXeXmXtwnVzIJfbKyV4maNx7Y
PWwgtMZiVnq4qbUlWDWVDbgNkMfi+u9GhctMUdWaGDBRllKuD+9GHKfgai3TI4JM
xqVwdN6C2w6vRDeclw8FCNbBdrGs+5hV+DxdYOcCMSbEXV+cXFTNFEk4QNv8OohC
7k6XYJiKqLaFdd4sSseAFfgpqqvjjXmHSBrCLBdOrH86CTLOXEMWOuCZkYu7UA+5
y0RyfhXCR12fJpByVDORlH0GSg9LDU9AY8c15B2sl2iEiUxcuFzbyxRvEWscZgaA
7um5WXl4Q4eITTanHlpfJnzwwn6ug1iiRehzBI6nvf4zwZ+s6EEzicP4lzXN75s8
fJ6yXO8yDEho9lQAoZEWct8KvoUXGsrkz90E4bCrWLQN1DfrYM0HpczRBv9uHfJz
9PbJO4XcbGwio2CTWkHv4tEK4ke7CRsP86RycAv/l1HnVVu9LOpar6iqK3hWmBUe
hy+/BTsoagGqSaMhqDLD+OeRHgXZ8wS5rguv8EDSgMR9UpLbtUAStc7C5ZgmXJAs
qxgXXpkTsJEZYYqZK153g49jas7Akz82XzkKK2Hpo9lpYmqpQbImY9UoGf6W+Axj
NgrwaeeyUy9LS3t6npV/72FOgz5ZbXVNIX6HLGDT2L/kIG1Q3ioN7i6o8d5JnU4f
3x/3PW39/MzI1otEBjnzRtfBlMHTy1nRqFsJ/6GkOBlHSHBIrauE2UysDXaRkaoY
Gt1kg1YtRU2IDde3D9XRkzI68xedSmeI3NXwci8aJ0tZRQTya91RfkK8ARUhARxk
WnZ4YwYsHGW7IwGR8IJtcLQDdJeCshVfQrsJusR9VaAtjthg3J1HvOacXbkYIs1R
KKPBkcMO6NGT/qeHt+gUCkLzvoWiJa9lbBdJR82Wa2PGdx6jAI//3eE68/Jy7IWc
yixtJvhme+mR+BStHeGbg8kGshbRtjcjeFe1rHsGsxBnEtGq7umvdRUuq163HO0I
RGC7HeMV45bTc7+bPxS3VaKdGWrubFT9vlLX4eFGrKpYDUAz4VRhH3HUzj86b0D3
z+IsjVpghpEq3LmddShWLmimxSMeI2zC5OiPwXs9neoqk5Dt3RhlqwQKvXsTyGZc
HKwUK28Jwps9YeIUIP/o2TyhkgsDi4yQL24lik2DfTps/xcDeKO6dvpcBSSHR7JN
RAAkSrJEj1yvStJyMWrKmHa0Zzc+7Fi1rco5QarijO0Iz96ZwwTlyEa1dHQHopD6
EJXul72ipfRphVxr9T+eln6E5RV634CjtG6pxrcP+wR9suIW1xAWP66gEeOpTpgz
CE2n+IEp/ouZOzf16YQi9cqg1X/wjOpSM05nomQ5/GRwonvTtbLxeyKqtUsOSWAa
uBgzfpy6OV48WQjknyGbzITkwkumysR6u7o3Aq9ohY0kTZSlM/Yrns+MZryO72xv
hXdHlmEbQJFeoX4E/AWJgNI6y/zrO7HeQzZQCP/uvl9YJTkggqIdatd6aedbmmxw
u1DH2OFThvdkDrmYkMFFvQbiVuUeNGw4ma3MKjp5wKIhKHgAzkKNO4awBV4RAUh6
DuvBVMbywbkU8jevgdfDKHO7MmMpKwSGiB4qIi+iXEBfLJItYOOSw3qBXanyioDd
v7HTLL47YlnRwFi6Okm5+IDX1IsZfLur59Ks+nqH/WQFBM9Yuo3NSh5+1MmdO/n3
YJG0IFRw5RR+Q6l3bGnCWL/pFr9HSbrJHfmcHKNKXw5uchG+UmPPtHdFexZQXYAD
n9O5ZyJu+1PJJs20+B0mxYPa+OBXSDVK/uLHPNNtzYdyZCimkaGugfGoH+Bzxfgt
rqKpcV45ZG42KnaD1AQkSX+EpSbQ0839Td6weYr0uOhf6cGNRK575Km9dAA0XLuk
eL661GloP8JO3/lIEypS38a1zkoI4KhTe9S0d9ZWL/pblhgg0f9wm3rdLe5vmkeK
38Q1W3xxm4FqRpR8hDayulQi96fYRzMlvZig+xttF6ig9nq88gNsPU4VUQ5RB5Ip
wJIXOgWTzaHNmxxcUwMIjUX11QS3e0eULFOhoa/ZGe+NLojrk91kjheAtifdTgu1
0JeTDeFlHYfCpUkbf9W8pzG46y/fRtNLMMe/etlCaBxkIpn8v0pEmQk1aHI6DFQ5
SI+2FQzesW34hI+O9b9Tbzu9NY9xoQVz5e6+jM/fGEeFC+AHL77qLTAqRMPjuAFu
2YhF2u96nIZr03nkSClrcoZhm/3tkc/zQLXF8zgrmm2ye5cxkf9AtbM8iJNO+fKB
VSojgTq3teRM9XDuEvB/wfScGLUus9nTN4vhZDh6boo1Y9sPMrudpylq88ca7N8k
gGzcLNRO1Hl47eqfYQVadt32oeoPo6BfOUMKAZTnZDbopQTVUYdQszLwR++qWoNq
y1qciRNE3HyL6E1t3ho5P2avNCDCRJYHbFjqqp3ArffDWLrafiR5hViwH3u6WTt9
Or+erG71z0CU3bji+l3isVmYZJwDXXOlsghqTnVyZl76NKwzbOE1X6qjyt0zOBN+
zZPzIonSJ4HdLYQTtStgqTuZoAvZoTH9WU+b0UC2Qh4k2duxbetxpBfRmhUikit4
5KeLQi9/8T1rn8rlZHWVz5dNFHbGcvxXsO39sDf16/l9e+V3PcPImtkI62TBoLUa
zAOO7wEiuq9j0Ne5G+5ZyT8QwP7Wc2DZCl7W3NYQBeh5qw4PMpnTvrAVKq3ALy4W
7pJrmhycOidJWgLhZVW2KO0nDQQblqBlYYBFR8kfeXZFW1gHUk2p1xtXtdmJJ1QN
gt4jthwQS+qflGO8BWq1a4aZ+Y3C3I6sF7QbpsthxkO0p9o25Jm+Ncu3U3SA/Kfn
hkl4JSf0Y0jzeaOz8B0Ql6FVYYUyNj34UOnKkl5CTW8WmmLqyX4ogM4u1j1sz2dD
PxVL02w1fJgVhZ6KbvDte1ZrQ9fpauKDyTlP1qHtxBu7+xKOWCyDzb4IyJZR0tOS
vNmA8WMOMbB1gftODmPuUnJsG2QXaBenrMKagldjV/5WNMBtk3BXja7vAiQlZymu
/79GXSPKFOlnHcuCiBq/2eg0jIYggIWJ74NCTjix2GdAMqDtN0LzcP8UBJAlBP3g
1RMa05DeFxUdejOJwUrZ6j/BSWNu1kF1nSIzhOnP99rXHCyMZ0g1oyTP0C5JAVFX
dnOFDRV0fEqJXh/WDsL0RZwLZV+ktiovBba5nrBGfBCEwJGNC+itIzZ5zRosaRt0
LrXR3KYzg9KHtjh1WtCrymLMNBdpdldP83QUMX6YRjPdRO7NhTcVgUawCFZDqCKS
ieOS0XO08/M7BXVv3DOeKAyC9OX4TUiW86Sk39EB1wxwnX000pHl9xt0YLU0Jz97
vVKc7pZFHyHGfQKAoBARdX1OEZRESnXx62FRlcO/t7gpzVyBUXLoAAncQOzm9J4O
/0LtFeqS3GE58Jyv8mv4LKrdaO9z3X2u/FRUs8aNE6nJ5DvvddriXKe5ZgdLuyrV
9IrrQrgU3vanCHA7bFdtTn5wFaQA8jQ3m6BSLrJgb3HeutC97aFBmh70GVe5zlf+
NZnYY0fw9Ru890UoeSlspgFYjF7DNDu7D42uoVl4qf1cr/3dP3wch/0mGvMJoNjr
v/G5xOOR0pscEKJR4Vxm9ti02YYXrnHC5Ju/Jnzq8AZ+Z7xpVeBRR/Luo6I37qyx
HFyIpD0FsApoLX2/9zFnxGRHIVeS7NBYStK7lnfpU8dR1oYr/zaRmjYBGu/yfarB
JhiaEUbFyPm76uOwe3VhiYqGrw9kEHjaPjmIFz5nbzJu3KTjcDE+gaArtcCCBY0c
UWsZvPiW74P6sNqYXzpr5bxupj2J6bYa9gQGAsmQSy6ElSEOtk2pWtm/2nhD/tIP
HitbxvU5JLGrVgnYXqkNe6qhf3Evek6I72vz5OPf5naf//1OreDvQdarpni6608c
8UiG8NhPVA6z791aPED8ozL5iCfInEkVKwAm4LKwfBwxP7h3dGxBu669/F0j6gzx
dwPim4kLO7s48wMB4w16UOyZwYoiaTJfnY8LdlL/Vf/xTp0cvGTLqVxALPn7l/cW
TK9E63gCltkxmIZlU+itTTvq7op6KAHvM7Rii154u1kBsqnBsdJwFyjKWTSq8ydS
p+CYlzSZxoPeW3bvIitIDqgUCfeKZuiuMgzxZMxlikPlwXCtQJiyAYi9L8XNU39G
+4K1RzeZTNWwXMrkrrbX36ufB2p23pPnpzO1NZPxNRCnLxAh8a5VflkHUAATmM4E
9XPoHduzX6qdbE34EhBfYr7da0kxuG1Sieqe+qbMFQV/aP3T7EICc3A6u77Lque4
eM/4lf19lCNKt/TqgAnd3cyFy7EyZYNBY0A7oYhIvA2ICM6VzNEfsA8e8syzqxMu
HnuhoghLZ5p27Hid42IP+pW9wQ59FcxHYB/O2MC11s4DEi/8KcqvJr/SvuQGstZ/
8b7dpH4NR7EZunlFBgxcV7rczFXFulLwTRAFh9ir1rp+NmWcmcoAeEKM6OuQM8KY
GpV7ZuGZvAkdHMFijPQc6f2NJfmg/dfmG1BlblRValJ+BnyYHVQpTC/bCr5UjIux
nAEaJ7L3y9DxSFLBnJnKThc83h51IWczv9O3b5cYs/TepxOX8MNZCQ6RzOjVSgum
lXYd+/TYNxhwWidayeiUD1v3dVaF+jV7wCWwkHTv/a4dc4/sc8fTJMycl0ma0w0c
xgqkeE4eWK4dK7jmwsHQDk3uuyTEWG/B/nmgUtHABczlAvx6RgpNuwDU+85TPt/q
A9E3QM7B7DXuns+dKeeaF3yAtHmxI7Ow/XQxS2NEWPqRrCYUBcaMdS+IE0y1YEcr
5nx6m4RidjRY4Do+zibxtGuMUvFqjFZh7hnmHhtfrZ+svO9CiqnKyXUnafs8J9XT
lwWF0mLZkvhqrnjgv+68w3O+Oda3NmocmSdnb7eI9eRFu6aj7eGUa9MIi8wqV3yf
ayM6a9D7oawZ3i9Dg/0XbZRDpT284oraHWCb5nUQJAPO2vzAxfoPYcjwhA/AFD5Y
CJ8S1RECxFpmutgbED7hD8L4SLHSyFb15+aGNX00Q5UcP5KKxIM28BkIdWJH7IZN
DdcmQ+i1jZl1NbpBds1ZjZPO0TXiH9kZbI73NNhSoLMIz+OxRawNqD7rK7trgA6X
7gI9wvjyxdKsYXTfllfkunmu0qDyuuojbaqrRJuuY2uLfDX27bLT++N7xIJLItkp
/XrRLPFoC0J9YNzQ8WaymVKAzvkrx1d9hLpIOy5hoj73FFvYnE3Pe8AWNWJydY8a
JdgtqgOIeS1fMUbLAydOvraedquKJuLePOFEbQkLNyNVBzJ/f847qP4EnckS+NM/
XZlFnI6ouf2LFtLDlZlKlzVDojY561UirCl/ugyRXSY5G2KP6/48JzrZf+Z4xbgO
hYWkGVvnNLaaLsVtwCu8aSdlcg3xwiWvC29AAAFmt7iNjUPKNY4tmR1vwbXgcUz9
sb+bUEEoMNFfRuWLIumhm0BYbFL+Gaqr6fNNS7GnwanbgKpsrxT2pHHRtvHWf9nz
y2l2lxCBfQBKbqnE76rPTEZw5TAyuKR2xikcjrWEV5v/HLS+i1tsPWhLyrfOAZA2
1guoMjJslg+HM6dvog7gU9+Q1zQHg5XTOWCu86/ezbuW0cNfZktFUmRUiwaADxOZ
CSKcHRaM0veeB9nFEJbRKV2f5n8gKL20ILKiH8Y4Stv7uaqDjEUMqNbsfHigGP/G
cWs0UCFaWZrY05YtKcmt8CcMyYTAgC2fF7IOX1ie5wWGeobU6wXcSqeVruwqadm3
tJdWnulyiDFMbfP8rCC9IrIqbjWEs2ujlvBYrCA0xsRhABGi9goWYvNacZLO9APV
rwD4//06LIGP+SebNdWd1M12C7kIGnWStK2ZS3lNfNNIEOAkvAetBTGnpB1OiwxF
wzwTF/SF95fkBAO03e28UuVEpLOMF7VMvSFEMFUqQssNPwBLlOu+iZUYasqDFm7T
tl+ZZjijZyfmDcRnzjhtW1tty+QGD2pRSG93oE5KdiN4p0aqvFUhElmzqHV7NDL/
3CdJs65LcgYAB5gVQllEIwrIdar06y8EHQo/vEid/DqMV7Ex+wXMub5y8GnF0PO2
rc4G+5DwHV6+90FsfrdUoyy4Lz1cTFnbXoLvH5l98hpoHw7ky/8JEvOWJwy4NBsI
rISM6ncIizVJz+N+lCB04fYnug7+FTD0w/MahZpVR3/b8jm5PfTYQh2sL1d/yOZT
2uN70LiwSxTwySrS+zkQyq/fhxPYvOlhbQzHL+iEz0BgODYASq+y1oh+32Tugy3V
03J0n+wnuAg4bSXNApoQ2tPOk10bsXWErK4jUfPj2YsgVv8RoNNlykeKxbkvSIbP
4pAcTH33D+nYUgGQG5PWSLrkrQ0yqgJ2zhSoh9suEhcY7p1YDxFum0JGpFq+JaEf
fGCnzZBwq/Oi/hGFG+YSonJJX0QX8KCVB2O74vXAn4xMDlYWx68mfe17XuFpq8gF
NROOVop56FLjqPqr+T6wEgywj7+yZcXuXJLUDihoPVfdFFW8qFhtwjjWP9uibYo4
4MhXAJp05WhhRWcneYMsHmxtwN1w94zkvr0CKU6IydxfxK9kpeH3jDGBJFDhferE
INu2WLGxeqyXO7y7R7K36GTO/LkVfpLZA+iIHfNEm6aEaK2PDouUJJkB+ngKVv4k
M0XtftF0oVrAfannaVFewX82YlGjRVuzCJhWaHG3SWeXjGOvdmMEiE5edfdc2x+m
jOkiuyrBd4O2wjWxPyDpaUpDHCLjdg+oOSpTAAWriq5eMVW7Vkxz/lVEgDyTT/ft
+s9Z0gqzS8gzTzNecQSKYNV16/S94i5/5Bivj/Ji8ujK/BAEWTH2im5zMZzckiHq
oZFesq2eATBSWLAF7Ae81Vvm7YzQEVDZ5ZfxQfSYlXjrHL/ucXso8JIi6TFcJqqf
Gel7MvV5khWOYuT91FUAw0NHq4uxzafrhMp2mZhx5QD2iGfp6RujEikg0zz413OP
PwhMpDkRM6GSTE5E16MDYYPAzT4OLNK0Bhcgkr4gjYeDoHYklAaJVbx8uBsZpkTJ
+UXCvXibjN54NtkzyM1PLyFkEddGYdZpujFX2fWky8NWN9R4p/FUnRqM94vWdOst
5ccHMq2Jl5z/F5s8fXdg+EiZTTCKzrhVnZFnFajlPokvVzdGYlMbOclGjxK8C8I4
Da7hxITaBx7U9n5TPg+0MI1kdwasHAf3xkvSm1xEzSqteN+2oySROuwI2PuXvpvT
ES0BkdAV5PJ13pA4i0+kMkKbj6oMeA9CjA0CPtG7pM1HKhlUJqdQBWytM2H4Jdgy
rFiqV8F33s1wDV39VZOHJlZstHdNbLfj5C8F6M8jc5uNv+g8DR/FK4/blGQ3dRT6
9bnU5luA0riMHzfEpy2mp0yj2/LROW+09CXrA4izGWX8tN82KFaT9Fm3kcEaOnsE
X/ZSg9RHBYz/EkWQLP87OuHe/byKeKb2rX0Fnraeisu/ebcVrWoFu4Za51wTu0Kn
88MNmvoR0hcK9/3KeNVnNqD7jjwslPcfHTgwaIBFyopTA0QieFrSIJj2ingpoW+s
a0qJmbmgfGQEfbzX36Le3FrRMVF0piP+r66G4SwoFkxp4R8dOluZIzDCqXAwNuE4
BrALRb+ihsYd/DBZNr8ROw79tHUntMPt6V8VksYhIdjL/4rZ9UxG4f+TCl6LBzzS
VeZ93pASlY6I91j3jpQuFaUhIjqHqAxymndmyMf3N+1WLaCXzM/1gTo+SUmWJFVu
tXVpVxo+RCQEYKYwC/3D0CH/iOO4xVq9JhsMqTuVmm1b0/9PVeunGOH3S3iHW+kC
scnK6IYZr0pQ3tg+i3trEjzy0XTFGZ0WmzLKANjNW8df8Ce08ZyQpfpwonmJlkfH
pbVeLiUn6+7IDx5vrYRXz753D0dG6p4W/roPsVmZDUELjX0/XAhaY41hzLSAetvU
ABvArJODlVqNt5o8/H1OYQpsffYorhalf47w5c5QznoHHm3vmID2EUa9J1BSguj8
9Q5+2WqbFRWRbpVmN1qaaErM6100i20vyXW/ptU126tJLhb31fQ83VqN+j6r+Br2
QhRgM4hz8l0wSONCglwvbOGaptTBpN/Bd9lK9L6/ej3PGVyWUyYQsW1T4Kc2mbOa
mYO/9MhF/ZA8FG7LunyDJegoe2WOu9sy1eJ+XFXMJkyBd11MPGPQRYWlzZVSLb4i
6n0wdQnXB79NZkTJodQjCjH+Exyo4096vrmS9j1mo0Qyl8/EBeeU8OerogwDwzbw
qUo5LjKVKhxphx59V+dmjuvgWtDGhf19h4gd1wM36l/gu/f+LQlGZM5UN8ipNnwT
Suz5UhAvdR3wEJFTcJJSPQgBMRyjyCoHFCeqZRcmFzfSP4E55NgdKpeudIGl4ZuD
u5AFwwjYc0Sjfq9YVVXSp35RRnh2aUfTuFL4Qt0UYXr41NbKkLNGFU8JLXkerRB4
fPzqnaE2L0omaH4KNpY/75leWt3lkoCrGNwQseMB7TdXNkX1cdzuOXCiKV+bkZlC
e1BO1jICLOaYxvtPwE75z9eQFta0UwuzzVbMnuE0WV41yE1if20oGS9M3FTcnmRn
9ppkHXC7X0JaUB5LmPbRQjQ667Aew0GXLxxXVrThwx+8GUdOm5vIfnpIAHyWxkdb
+E5hSWlDXFqucVEdNBc+q3f4DSVPfL3BrKAQjAn8w1LkwIvPLTylq3mV/D1SeRFR
9YkLxIvkz7R/9Da/InxRs8FsK0CZiaI8HXbigvYKoz2ZKRWOVJMEGhQI5pD2FLhy
96Lfjyva3xvpfb74GYP0PDCEBEMiPinQuuyjG8KWUIx5mRBngNSGGbm0uxRENZ5q
MJRqtFg2h+zN0Xa3hYxKK1fcKbtK+nefqA5lv6/OtbvTcqzwyMg3vhLSAto4sbDo
pkfPXeqgjj6xztdPLg3aGv52XHBgFG6P19j9NlFPIRuWwtJsL1JRBmZKePofuyra
XYCb3tTw6sILbkxRRcbm+crw9dnwaGgl4obHaornqDMS5fetv0KUTIl5y7dWTw46
xoeoYqvO/kAMxJoUQbMngQKY75y+nMw+X1n2O9o2w0jQhF6ZYd9OKMtEVbxTcXRt
aMn3CaMJXizhMQLYFgcw5LnGHLFbeVyfCvmRRL0BtAJZaPDg9r13X3u+M0ssPuwk
yV4BHlUqj8DbYGratgTVwhgEiG09FvnB7UxyrPHOuqR2TBCJO8wdz4t/QGrqooBC
d/fn+pTvVt76+nZWqZN06sarKTe79NJjCR+jJfzPeVg6kgetsdmqLRhRzTbQT+g0
SwUFs3NNPaTQITJKfw1y5K3RFas/DMPY3awDpdaT8U/+EsUJjpGZ4daq21zk0aU0
+Y/MAHTiIfSc0CgHaW7USEh0T7Q7QQjkI6dJ4FSa1aBE/3uucMp9FmzSSI9j2Kto
QDl22swOBqYxtD/XtKyG4RtHgcIMCFCmjVd3Rg30+u3lgfuQn6tWKMji7k/QMlZ3
l4rnMZOxHqMhtCr+5qlSYg==
`pragma protect end_protected
