// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
imjEf0SZY+01P+3IeH8z/wurzcP0KTynODK3o4LRN2h6UnZqOvTRju7uMomiPuSB
/Te1ldxsK5Ce1/OVD+/Q8NdYvW+v88s//mO4SR+ek6Z0g9C9+8GVxYLma1d7bwtH
EBGtsLOlHy8BE3IqUdE//c3gmiZgLwOcsys3vX5Ozd4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
WmIKSJDQs5BvEsbGh8nzN5n4OW2vnXV9AJjwdFVX8v68uCM0PxYr9kMHR/Pa2qha
KejGNS1vJA2IZQ2T6sGOHya7/rGFkv81VWj9kgllFjt45E2FTlY/nXnE8FhKeIhA
NAN36iXfvChxr8cDqeePZmAFZ56V7v3BYURAfhTMzMrIO/qty+m1saINuQhcBP+Q
b5/67QDNHbzVxeeCzRrPTQq4SE6kkrTyBYVeph8XzVf5Z8GSe7wo/HAvdBZXbtMU
0ml9ZO17vgmm3hCRGkoconXQ6gYGe8y0gu+SXBc5NiFxPbSE36K1KqcBfUV/v88y
Go4dCXKZwAtO25ASkor0Qyrsbwo7f6vuB5gMUBHtcg8/75szctpvwy2UmVMVmwWg
6/9o8xXOVYrNUvUMi+r/YHp8u5MKW2UnXnFw6jKMSByr53kSCMXt7q/TfWgIgDOy
k1M8Py/Qt6skCVSHRmhejq6uPT7xASVhtqewgyu0TbypYBibPrR0i5B6DNYBA30T
+LCToB8Jmsfz7086zKnjXpmSd9eCRxnY+Vy+kvLD5K6Taj85ksVep8QbbN+7fWuy
4r8I0Tzfrt/TI5h+Leqsdiijen7SQyzDmQFgJnPZs/T+585hSJUoaVeWRgVsGF6J
9glgUWzrHEA+zpYA8umlSfdssAtn1uqrt1NRpTVsnnIKQ7LMdthecq56wzuX1IKp
U+QLYiqV2yVgqQ3p1QmWFp7VfNHHnBpHDogAg6XacZAtXwdKl+Y9Wih0so8/Ab7e
mRUi2OE6bGTfxFtbwfAGNBBxXmPwyzmi9UaPg7K3QI+cICJ9LH5CXiI2sjosBQwn
GWnRKrCFw6kXTxF73IRFU8aVc3zQfcYkM012KpSESkPCSj0uL+2GZfDVJbrOkXfw
H4kfW6vXf/mVRGCX0QFllYt+PNnAp3UipBAah9vg6z/wVV21eThG7tLTas7K8T96
5OXpRiI009X6glOFFoDb0S/Os6xW57zoil7ujCle/RqRcm1FFfPwPnLB7JbvbCiY
ZMXA3McuXQ6YDGAiC83CBAE+zRe0Z9iHkAlicfUSBwz0X0cb9cQ7VK1WA3VI7xdz
8h0FJcxd/jUCbQA8llsqtB46AF5voSZ9v1YW0MOvkO19/ZwBXNWhJhhz09UbV+xV
k1KCs6u/12KrASYmJ/1zX41v7xwHRvboa/yGfLQECSKxcXH2QuNqWXZ9wVewmP+L
UB7Et8eMEdl+Zu8qfe18Gle2ORR9BCYzjHBQfQYAbYdOOm250KkyjsXAser9/w/J
YYpYBLylpwvdm/mKm7c2xOz4erlttiatwI9stZ0wBGEFUV3me3N+w0Iux/8ZqXC6
2wVy88yoiSKR595L8EM/aDKRiyhB0vXdWm+2cXaksi2JoRO6yi1pERSh0xKil5ws
O5bTuN+uEnSQ487f5Oj+8+WcrLcO588VmFaOREgGwH5/RdVhLx5LAhN3t1gVkCkC
V1W5Dj7hXnB8/G7WkyWBqBBjPoRRPrmdTGf0FOoLXASZw/0Gt0bdesTNisQzPt6/
RH6l5UtbIbj/WsDdsfTgNuBn5d8x1mhld/P45v39CIOQxe5S2M6d5M0bVKJXE3Fg
61fKcS9XvkGCBgEOxrSjseKLi0wcT0X9SbKw1KTGm24JbYOrezR84pu+x5TyOmTB
eIjG6pQ9Dou34WInEiW8nNb7JjQri8uy9Ub5SSJb89M93sdjmy34ZwL0dhX7q+Mv
1CuaKZ/MGiTV6SyKl+L8HEKALeYRSU8YCsHNaEbkNSwb5sAqCtt9cMq6GyZjxLvq
KiCnY0+AwWOyH7JiHkueU+/o1zEpFaQjIQ80td8ycmahbveKblzA8I+Mwdp4f8t7
z67NYjskj5Wl5/c9N03mXMfms4cOqM25CfhWU327qWyrgs/zvNhNWp9P84QMF0zq
enOW7C6RPxAVgDAJ/WOGvU8xWutj6FkIVUq1HByL5q699wSjZuspqOwB5idpOyw1
6CUEX+ORB7yD7qeK2tSxr3K1u0mT9RBUijHc78lCz5EtPtRezoiWFv1GF3Uo5pK7
GMnwwgwcZwq+0P+j3fM4JrNgIGBzq6rex3bmpcPiLWpcMHqmUJuy/zlyxpIQ1Xvk
c1f6yLHIObQ0J+5N4vVGezmu3pt7TWqAOe1RzBQoA4Clb3QC91ZEr4tLSFCU91zZ
fnhKYYup2N26c8EavoVv6+9uCaLb78udEmiIotEB7G3vARSdZjmLbWSnWy3w6G1D
zt5MDUsTTXpnufgK2u/FPlbclRzicbS+qtAucFcAdZtaUcOu+c6xF3dwf4pE1Q19
RacnTKONNnKleSz3Naf5NNmI/SEG/6UBdOLBmwc97mmRo93+wOmlBkOLTnILbv5j
5hmOxYNqIVTFjghkz2HQpeXqdaAl++47bBivUab/18usG8qJ4F2qYFzhtF4sKQdo
8JF6EkYP5S+3DMGfEdIJMdi92+t5fyB9yW6h0THyzKX7YZSIco/2EcRUP20p3uR3
JQ0p6CwAjiaTFgP6ns33OU/maRKTEMQ/WwfNPcNpO8ox2CMB2VTaureQ7Sl32xkd
DjyJPdiegZsULVX4Z7i+mocqUcaCZ6vUIPeRJ0eA2Rx6qcmmVSRhXc0aeN9gqnob
9kcFMi3U8vOrcBkm5yu9EefP9E05oiuNGz9AEsiqogk+8Ef93g/VLjlw/79oAu0D
CXLkaZdCvYiC71/lmIJx5ib1hJGkCXv1YWXOEnCR7E9gJ4WLpdcjNWYMWJZlQU6+
2gC3yzpIfuUE0JtpY9Oxp/yAeIa1oNHngQruIpmYZVLmGRKJykBQeF1qK7JI5Yjt
1nP3Y1DFvhbb4M2mTOc7mQsGJmzXbhHQIOhmkuT+Gz8g0WLnllD6nU2hdB5oYVES
DSDz8mlUsaPUuHeAcXMcCVo8lCiQlK6ICCSzKTY4bWxX5Iwh4VGuW6hqthe7+hqK
NakB4nN/FB/zMgu+sNrTFS8T5k39LfftaXghFH4mA9rtVNioXxahuXqL0tYGTI1T
uEZzrl25wPbADuEH/eS+hcf3urtGCFjS93EfpQWBYrPzt3H9YSnBIhFs7AgvWmIl
fBbrOx6IOjySUBtHirG8QjI2TVeieQ0xo2OKXwRuzD5GnW/WW5A2Nt8803edE18d
WMCH4R1SroZpAePv3NAZkVYsBxIBBYEIEoFQH7g6uMfSLIEDJJIeZ8ojkGlsKmnx
mbWycJS+0Y0xajZ+fH8P7aQyIq7iYFUtN+qLJd7Fv7zm1Cek4TpOK5eDVVopSCoT
CQJRlMj8DV7jhshgoy/Qo4u6bqUj9aW2k7enDggYM+Bk6nnCRuroAdWnjS67oMaW
9WfWxlm1jv0zfhRoRV6zacDn7iXit39nkrB+JQvr4i+AxkvOieMxWIkQXwoRcvz/
KTeznxPFt9mOw0PgLWrvE/kPC/QhkLu3dZ5NoyJ2wetOhTYj84PwZoJNeiltYb4p
MZkboF5Msu67yLQdykS1yvStQCMeTUjF4YCX2+Ry+ydCRr1doHv0UySUKGgSSYAf
Dpw/zlvGx9dw205W3I85HjYui+7GlzUkLJj2I+JG0osE0EjnJpjVtvqmEEbB8iW4
4LGslWDHXGjAChQBDiFw0OO+I/HDT+oF5TbY4M1NoCTVgyFHjVyU5tCokUN14Uhw
kKl0Uv95WwxBDLAPFLXOs56650ddRiRIuOWC6wJXySO4km02Oz6AetbjD08xpBph
+KbTpx8QfA8ophj2RxGmUc0PAPkZMz32WYLz5dJbm1n0I07mSoYNFrDVTLfk1Z3u
zaNmsn59jT+LIix/K7LdjIVMXPaL7ubEcXGJfxBtDASKOiqXEpo0rhlx75kWorOE
JYlL6I3GerbgNgiuqa/bis+WArRlWpyvR8E28OtftoNX3nCVG/ZYMQJhR+ZhHK17
F3ugg17qMGjoq+fq1sQANqYFYQn28L34W9kQDteBFL0pI2Jt0/3ftcBEV5AvyziH
EkHyPrYeg7uFDHntlFDvq4AtrjePAYVFtGgkp+n3QfHOI1z5LhHEpXsAUKBFrxtU
HJNZ/tF2KbTzOrnUSLN7t27QiCAIQBPcmi3Frdrxd+j6fBR4XZLF2JuEGdcgQ0oF
uOkClhhZdTHnIBXOP7y63wX9usbYEyxheTyMEf41YZag1RiuakrPuE8npSVAw1eX
cZMZ3ARwplCnxAWtXLAzQ4x0LYLgtL4+ZrCBOFdRme7PN7Pto/yj459xbVmSoph2
jo+VA3MnfECQW23PEVqDRSg18IcQ3505PAmUbjac5enBVCBGmt2glTz3QkVwaNuE
HrAy+yZ+5fRzxrtClw0mr0k9HfEzEdsatitCFRmf1lz2naPPEI/cPi3A/EI3d3uA
ofV6HyGXr52NkxMDtryriMNU2g5KeBRfw5Fs9ENFAlLspJAoasx3GpUmS3Pj5MBh
uS8IcW0fz4grCYZJo+jtmP0Mpoo0L5BNh54JB7kJQNkbfDhwQXVoq4TSRU+HBS/Z
xt/ZiBkbQXv9CcslRBZIPlt5tpV84UZDEWYdB6e4fc/r2fc9DMlMOXeZlXFy2CbW
mGuhNlQXspOeM+PPE6JM+pBTUeTeOeTEMDsR8pgyDOQRoR5Gc+dMV9UAOSu6VurB
W4mCFi30UfO88ZH6IB9yaxJZ46pkYuXJFGWx4xdoMi0wMODWgcIcxZL3M+W8NF5L
aguhrLHbuzPivWywkAx+Sv/g8ZDvI0haiopT12GwrcuTEmcbLgi+T9vOnHmztpsN
SC86XDkBEwKO8l9TFwwASasbq86IcqZ5rUBTscIVMKlgWybb0WcCYd/330o8QSqA
QGHOD3PFENUgrE6mPutpIUy0o0gEvF1AtMAPL06lZmcUiSCrmiQFbp5tSwwjvCWJ
PlhhB6cjU4Ea2oQK0ZO4+UED3ooua9gVNDkgeSIzA5CW6VEZxPANLFnY4rEfBjdt
jCPI75BQ1qi6RVlPua/hjaEv1RzQymyudsvHvVnYkFvmFpgRe1GLTuOlZz2JnRbE
tlVVLmuBGtUjfci89EDdFBdQhI7nRU095QeVCwYxByLZr17uvQ/7q3wMUD2KeUxt
M1m9nE6fomCgWBuUCczRg48rPFUpUrBuZlecNl8FU536AbHQGR9WpSIbwVS1rvB6
RBtjWDi5A+Hx/9eUNaU9sB78AJLipvn9333TKhc5RWpnBr0NnnQCUagfYCPEarQ4
M29dF+exqztAG3Mhn0xuj30rpdV8E+8y+srfpBap37QxOnE1GALf/7bFoMd/4Fvk
Viuwn8KgYMrT+o6Fz9hyM6MJu9BsQ2mQdV1MwpR9Jiy5ZV7qHmzT7HFFXw7AO5fi
vKJ0busXguK0mMQLHCsBnwJR+altdx0Cc3rlL4xm78xgqvukSl6EbsejdYFW241E
sludwZUWAu+8zGWeNBMWKtyuJwSgVnkQ6G8JfwpDP7t6hwCoitYbESVSwSRYcO3n
E9s0yhqDPDVYrdsktU1Cv5HX66QKC46nRflr6Mgb1pJjKlWROh8RCxAPwg8TcQ6E
rGndIncxPkUfwL2beR11ioW39WQw7ceUO//6C+f4963VdMZ0CyOAbJoZRMcEDDMA
gK8a2FNzSBDMEbzBh2JnEbJ8hPaiqVjfoSOPbrP5htNbRTPqKgpZwSY9HmQS1zew
/iO+5KK6cZs1h7cI0e5XTkD/y9xyj1IYKSZgj2s2FCqStB6FyYA37Sm+oOj9RCzM
OEI6+6dL7PTXib9zoXH8W1obtz4q6Y1BAyhakkNfGYSpD1/trfd6lYKcXDzIw2JO
9lC/rzwsI3+a3PrC948dNtezd4VtX6gfQ6m5xugk+o63cXr2MqYMKsQ05qDOsK90
E4kIiUoAEcLf9kAywDwguLXIMO8A5BT55yGbrTOZp/HdTR13eYygX8zmuDS9subF
y2xTn9N7t0RvAiK7wiD305qkaaTr5wuF2xkwgYddU4IOC+YlmU7IifvFSekN/PRG
HWqPk+KZfxrPMmp1oay4AfwvSb1Et0b8h9DzapHc680nKVtlhHul/wGtGajKfSvE
ZPlh49JRWcPOTfr92XxnQUbSFmtsV3oz4PrMFk2Xjx+Es9o8xeMTTgVO001f108X
+ZwhI1TdX//Uo2TLzd8OE+KxLCjIOUQb25zAUMhl6gon0bpaiQ2YY5hHBycYHp82
i7TMksUNX5c2dcMTGvKgFxncEJNQM8WBUO25xfkpTwV31mZZKJ3VD5Xe9Gf0xlFM
Gs/FrocP+g3ApovCEMhrmrvt3uJFyuRM6P/4WtUoGLpc8M9pGEyrmacsyWXCH6X9
CmuU0MJIn+KlAI7mRNaYLhFyiBpPP8nsL87REzG78baTwukAtF5OVx5RHA5KrTY6
h+KdHzSzBWFdrU6kckd0WOJl6xNotpYu1Kd3GkMLzJS/tEwqz816pe1dCRsewIGx
9su3SnPCByXltt51KDDbYxHGo7tVMeNZww0fn1ENLE6HxbqkxnUqPi+DH0Dxevk6
lfDD5QVyvFhw8fX1zbN06co6l/DEg54isoNnBzNC4e2dcTuXC2+o0Hh0Nwrl+YX9
eMfBBX5q86MUAOyQ/Q2r3v6BaJfMWlp0oeP4Y6rsYiTkIC7VXVECr6ui1jFM//nZ
Qry7KRV+vmUsFa/V10+5oknclRTJHCbSDd7n+140iK1fSRlPqlcXZG5u6FB2pj5u
jX6S/R2Dc46WH1oIpA/f7cYs0o1K3bZe2aobIpAZqcLAS2poYSEUb1h+5vfZAhRa
8vCibRYpGtLxbZubP6bLcTWsaHGauhIZTIe2KPVd+vdGNnn6B+N/Z4iafZs6szyi
5VlT1dKoSz4IhAQJCgTgLTyTAqXtvd3WHyQBp/sphhLuXZEVMo4d5BS3bhwQh6fN
OziT/ZF+VVBO5fxIH0NzarzV1GFwQzmvdYNzmd1ad+AOrrEilK4g6HC/WBN2K+0M
3cTudHe8enrvJF7LhOq4RPhmwaKv8i6If9W5DII4efnwUXxCIqC9eBxvxj223zAX
15JgDGevtnirxv43d/kq6hWvFM1lAhgtn2Slq36iriTclBjYrIHdgsqAa2w028ul
4K03urBNrChAR/BSD3KJkw8n3JHHTNrTWMDmXOFODTR6nwupsz/llkNEcKrUPq6U
rAkypjmjp4zZ6JCvc8V/xg1cUPY7XHudbBpaR/28hx9JkaX3sY918ThL5hAxmH55
9HdzZxhh4NzdmXMTSEa44mVqjtPDVPqkmllWN6aTIdbeCRtnKz+GeDJSZUmXOpv6
gMsPqJqjSwNGjof21dSzX2XciIDNaBxC2OpmpqrWLMmFFRAhNSKIQDWRjVAx9xlG
HdJVXAt88m/5SgoELL/3CdhnctoqCIW1xVdhQAoxTMCDZ3fu8uaxuYyhQ4SqPhfl
z7OslxDgMDxn/8j62sDiMxSkyFR+jHKWaa+GHCW4OdbYPexDF5j+NEvmiMPib6UF
DpYCjsOK3Xrf6YmJN8P9yBndSGPrG746PYq8cIWwyZuLXzZdZ9+146IyBoxawv7Y
aZTGACrGueor1FJH9D8J8nC0zVJilyocl81sdalwbyZhFJEzELvVs27XA8COeWZM
E0g6SQtZiQhHXv5/uZDQkjfpK+l/rFYKxSwCeAoAZjEDYVEZKqH+BosQ8DjIxfE7
Be8uU+iWTw6AiTuyuGPyuhhu8F1t/3hXhQcvSmxijm91st7Begyyj5WcdPQEtzWx
TYTZDQgiqbGQY3+DmguVDDcFHa7vxTvYHTRPFAauHQpXUhtg8uc3w3LwlwdzSL8K
B8j8bS2gVpEA/Qe+EF48MRHUGBKAk/6VrFDYEHmT0J7dA0B5IWKtZTzdWck7YOrH
QAYGVKm+JBcQRYbySGIFWiUiFjXg1cLb3WF9IH6vHaKjflJ+RyriaGGsPTOmz3Cg
Be5Fjxt00+ETaeb6uS9MdFkEHPInX/CpK9k8X/k4x68EFpjajL1juk4JJ5zXNmqe
GbRR/QQ053CZbRuFKxxFHy4dqy+y3I/6NeAViYrvR7e4pFwkbhXqJ2Bt39maELYA
l7UzD2IozsFhGzqWnd7XWvRA/I0ujPAktts1PIinnNMq20ibg1PCgZzk0y75ImHo
81MTdOBEDrgBFhbiXqUNBdIFvMgOGTwBpGbgCazaniOBTy/wAak5G0uK2amivPvX
0qsSNvLk9frU4cbmsWh7VwRYK7r/TWvsheo0irnTf3NrksObdSiKw6cNIEp7ShYu
CkK6nGNv1E9HkUgMjrWuftcKM+8OXNdaQj41RclpMAVpzJn099wmbWlxqn57lA6O
KL9YIxcQ8UYuStlgwXyZQYEyZmya7VQXFdsKkIQmJkJ0Mix7i2HNM93VJGOp7Duk
4S/ZC75K1p4je4aK4pz3msaS5wvMKwr3pLsshyqyEb/+RFyMk34LzhCv+jZ7zh5q
Yy4x0G5AFv9Pruu6XTxeR6IR4GiCn/uVp9+5fbr1zDVRgve4+9XBDvg/YSP1vubO
cq8ORR+dZBuWsksJ5VejRTlNduXJ3lL1CzJOvMwzZ3OKGdYv1wHFZbqwbxJUp1Cr
Z0xmnsNd6+n/iFEYYc7kevQdpQvoSHfUW0G14BemMUt2PqpgUzQtlsAgy2dhAnNO
vruxnfAwQwqFYRVcq/vYr0v0IKEHRvFpN2cC5P0QvWUJxLPDrAnkyvIpyEx0Bchn
wzXsOnSgqQS14WKkc/eU16h8Pts83se34Uz8uM4rc8+6G8Mk9GP6rWqkQ+g4LLjW
LPSDQGbLZBig2Q3y4UbSiiS7fCVYm9bM7awsQwV9t2rDc9s3ZK8VB6C+8JXFpnH8
WnyYUzYubvm/geICpfOkXuXlR4vGZV6ezH5zz3e/hh02lx/PjeT3tC6DmVpon2pc
262QC8AVCPHr8uxcOqHJIL5d6QXRdG3rTAt8TDL6CSh9pmlM6wdcRWO6nxYJjdFk
6IEnGf3RwDlJGSmpyExzGr2Ikwr/ns6+s8mS/y0oZImptKRRM2TRDHFM3ZEII6ml
taB3c6qNQAgUwGaosL6fFNa25KT0hREcLlzVxNBpskK//0vPJ1dC4Ev1ziR02Qnt
oLVQG/gDgveM4iQnaVHlf75iZdaV+FvPSB2xyXKDDbJ8/KbtuqgB2yRC6s0HfWhV
zR594+uxMHpgX01nZge++1BVU7QpC41cLfWnb7W/MypZlw10WjJBRZZ3B1sHvOlV
XabCVluBu8JF3tIEB/BtwzQRCpPpIeNiYJYRNFXUot9yIHrI1Qf2YLjHLHazU5wt
YyxnPtWjYzUpmo12VXon50Evn7vIKDJwpZRr7tAodXRnbfb0ahezyyVYVeyV9in3
ufwnyxl549JB4YmmN/8HlUnjVk0GVEBNQttgUlYFxvuR9wCGHdwa1OmwSyqBMyyK
sRsBgt1sWVVCqv/t/MpN3xL1u9aUhenWJK311/iC74KWZplgj7LKaWUWEfy8pVOi
gC0ADK9TKAen009eJvWZBcexdejtffgy0QYReZ06Aoymr2uUOSAENIrJ+nIP62Cw
/YRb8VM9SX/o6Gn8l1Jlggc8bcW6rg9TS5gxQiJWJNiZPKOouLlSNtWNdoWrFAao
pYq+lcLnb1wo0zzjBH1eURdpH7UYwET6m9vKs3EIN9wChREVvEi+Bf8tFIaSsdC5
MOXhsCyIvP0h5EgXlgvwCckHRnp5R5qC3+dMENO4MLQk+0WVeodaiWg4j893QCvU
ygT1WzJLOmTSxEjWgWu3SDV+FreNZjRdX4b5P76A9zXgh4IQAdPoqum5MqLXXhHP
hGgmtWqF1tWiafmx47d3mLKnSvSqQM+AzdufFGVQv76WSARUof8WhijkUOJ4W2aV
uLv28MZvnlJrbr/VXtY6DmkA8hmAN43oDMNyNpIxmzpoeY4nuRwxRzjcyQMJTNsO
qwQ5pJheBpAgtHSMJFvxxSU6Aga/3n5w6giB/7GG2MPq+3GkbwGnc3dxIOabauBV
dwMIaH0/xQQwJAkcahw8zF3q0SFVwua8xJGA22Gd1g9OmastmPdWx/DOYAzSwtk6
DP6qYnAWvKItmHop3Jd4E+Ee4UC89ahTtxb4W0vbsyreJyavhryEjdalWQkgCuQ6
15fq7PbuoAf3U7w3ZD3Sak+jR7Jx6ziC0RFQlCoQ6Ytq7mTH9qTP8ZrXQWcOl/Zr
7Fa7KkaRJPzkedORtx96PxPgPLVogFHxE6sYhXe+K8AzMYr/byUvt39IIm2q/kY1
h+We60KWACYB/dKd/loJU8VPsKrdY1Kqlyu9tab1lgNKYZXz0Yzx46Wi/d7CJIkU
orOyO1v1orpi7HxDSL0k19ZeHXBrpCkDkR3xgasRNeK0qmcWI6CJcbUON7iE6evx
qlCd/htryafmbdARsHrx9ndK0XrJCksuOXvOOz5UZV5pczAh78xMisa6qcA0iL2g
8Cf3/1E+VwqMnsEgvL3tKCa966Q3xXWIHWGScuHslToCjO707W4zybGB80EI6B21
d7UQcKJMiAFf8btTvjqBQEIML+a/eDsYc8u5jl2laezHOFnGNtOUl1f39oL8hjrw
53C0SYRH3wmxeQFwY85hL2NOvmlwuu32IpS82W3xxTZfXRiQyChK34nCySNxaIL7
NXa/NK+9+0WbQ9qwGPFFc2GbYkz+HLphTcHi7Q38FI2cBEodoVzN0EwTTpxKJka9
HJLHNpmAXHBTDmVxuNztA2NXOQkMsVbQ3zrCqxVeHK57MNr+uLEQcDTlW9l00DrD
ck0digAuyRcNbUx5T01OJ61HYWgZ0mPuRoFXzqTOzrzmpSFak+7EcRm4qGuLFido
m1kdAaYvzhDaZUvcjzqUmDT6ZnfTjcTUYaJfwmJbuW2JOkyZFKq7R3npYMhdcGLu
bySleEcUKnDZ1AUbWu4iHwTYTfM/Djvw34CJGT575PqNHL1y0LyGDldvnde6X9sF
7p8c38GoNVLYJ3MbBfKKK4130M9kjAt3mQME2JkCRP8mNB0ckV8jl6UWy1Q6kQg5
0/QrE0ZUGwwEPrr8pMouWb4BlsAR5InUx8uZLyGPfHS2EbcERn0haH4toKYlMoeB
o3XrW6QHMvmRpiH8sfHWu462r5BfvWeNDBSZlAhHhHoQHBPCKz+2WbmtIl11ASmU
L4NgDUpGQIj0kumgXwG6zTx3eYRjSzhhh6T8SzYX20WdWuZ8KsgY9oMuLWIegGwj
SdFjzMdLTG9I6dwtse5+QypmU5mn2c6leAVm+QwRg2NmUvqZOrmRM5dNvZmfDvAt
to2hNHJbmVeHImY6SL7xQtYAut7Bbqw458qQKifLyTTYUSUPwn6QPBawNf+3GHMG
BVI00lytZwQc4wstHNbdcbDNafPZJTHDSzwf24983siJss4bDGZ6VWfYWYFoCjjB
8f/4ZqCRKhqLjma5OyYgb9cvQsR6iL52j4JUIe2LJTJ908WScdKJixkmzIKvTTD/
F2XClHzxeZHhzBbg7OiDkqtA/ipA/KmBviqJyZuAs9Vu2vVqFtpeSAQvNGdRDpX0
c1SP+xxyqqWPWpgW1YDk2gXlho52ZsNeYId4p3PFji3diSvREsRDUn28M5DQ246V
RHag0kIOlHxlmidPTjjLFdhRA55oti9RFwXHpUzLG8O3rcbm8TxD6FK1aTYr20Xs
141KBoOJLp82L4/RsueAHNC94ShXTrLR7HCS7bgm9+TYyHTgPeKJAJwwjZaf1ylN
dO83PpUTq5n6g/ikTX5c0R/jWal2e1zHmldWEJ+HprXUdHtek1hDtf8Pl/6ElElV
vdWzWj2YIhJK2ZNvTWNINKf98gLlTY2rKcCrMa63PmU65kDJuJ4p58MRUwCr7aBA
oiGInyFLyZwd/DnV8NcErlywkvpSXe5G+kzfIxh2L8f7Ai2h6SCyC+fckbyZ5+3B
3l0Ou3beO4al0qFz+oI46k4oCzGS5K1UHfEVqAO1bHHDLTqA43CWKuD7dSSqRWNy
bEbdd2fQlWK3OaWz4PsUo578H1Mk3S/xLqdI0+OHTmkw+ptrKcEXkd4p5ABkk6JI
0zml0yWwYUHYyWOtif0OycEtpx1+B8TjyBk3WIJErwAI5CdZmgJUjXXIdfTg8OLn
oZuprrAWaBbtY7o8OOSTcGx1ysFsYPuLISfNEeGd50bmVYnWVxDopvUuWE0ox5K9
be4SA0mkdda/fae6Xtt23BUeGAebSl/jSvVHBtcDa8LvJ+Bj8mv+8WHrguu2HYPO
jBMs3FJmjhrjxojjrmtPS7IMPv7OKPxKAr10IGmF8FrLjxpu5CDKDQf3s8ASwlwa
2cUCimR71eoXGmNI4u3o16U6FeI0qaCtgBbJitqKZrivcY1zwQ6RTSqcpgJMgAmb
jc2bWl7etX/rVXXM+r4khVEuAqRkSNB64wL5reabi2bxwtHO2ZXytufSUuerq3Jt
IbmXAw5CXMXPAFE9BmJWL1ei63JS3TrR60IJUShxI7G5KEbUZTUbzTmP9IT4D+Vo
ElzKsj/pFD/RHZOBSZBY+ZCHXxTJQmo7A8F0d9dhiS3akt00SauCXqrqT2VEmHt6
C/U15u9AL2ZTyS7kiiQk6LqOFkTRB+CqpY/nkRjlwrJ8rsCjvwLDNsxO/6OaV+gx
NEDWfAurFc+eWJ++GJJaOVWNK9bu8Y6spniU517PeVg8pU2ecIeEnO/wo3d63jvW
4PiohlCbpKOT/2GvAsQqYEd13he+0rpefxIyeCtJVQXx3QfIDB9of6+lX6uNoLQX
iHPQWeY0KBHYaXv1HPDFPo7UIWQvy/PpnZPxNXqdJ6FE45JrgLaNkMaXXndgBdC0
e5x1L+zKTR6ycKdPb0ns89c/uS4Uu3oql/N+jOBfqsMX43ikGICZc5Dn/KGFohDq
1q2GN1XIIOyqk/g46O5GV5qwQOrzyaSmuj1ZM4OqheGuiNjSjBD2MCTKmyUGb/3Q
C3lMcpejtJM+7U5fN0DH0jK+A9bjHDNwkEpvfGB4py0y7h79xW4lUwqjxSHPhhwU
vXIym8pdk1WgibLII7A4yQYG0O7Kyp5J8kJ9cwSlnqQFYkr6O96aDyiEsL8SHRSI
vSMaNYjZPRPor+z281PPHfIH8uk7ZWwaExbAzVRRlbeBG+uYgmzhJ3+mbY0FFZ3u
Y34xIOumtxynWwRkUQ+Tk82mzOvr67UdYmEuHqor1o+vEWxmj/PXMwb3OFZgLNKa
ftoeTyHC7tSiQ/k8igMElon7ZcpLts0CQe8X1yp29Rni8niCrVp+hSKkq0JsXWiM
/Teg6Y96WhU6OO5ahr1MJ4FBcopjz8n/0ajqFR9iy+g67F6/HMv5bdxB0ey4Vqt0
V3oGYYtNTS1Lobc5sx8KAPvMTieOsN5LuzYJI/myeJ7N92ggfwaWQYAbPZHyfuZk
C/q+SPOW69w3VL5DKyFIF8vJftnX9NJQjFH3+P9RGIPhWOOXEur+uRR9O9I6oMu4
CGSsMeqfwpl0l9qNijmF4Fy5n3hXv3JwRHPR2T/AsAN93W6bnrxAxLpPo9eoz8y3
P+Tjp54chc2whJf6x8YdPHs3nTusDAmG/f1q00Rj6HNlZo70XBgEDYV6upo+bGA8
0BphBq1PlD9nDyEsySBDxym8TWUE3JjJItih8ltDIq930OuZHVvMpcU9Kv8E2Qp6
vmnZ/FWkDIxRnZwQpXLg8Lzkuy0RdX8F8/og2NbQ93wRKjVuP5u3ZAWA0pt8BJy4
QdsV0f+iLg4Af4u2QoEY8MVrldWfhnCHDicAv/ALPyIlwS/ykNKGYAitYrc+Iau3
nQvPjyFChR9mtE2BoMkHLzpomORuBmULu7Z3nhtSSR2SZofnph+wEzXEoITAY0iC
5wziNG4nIYKpqUx8x96lBPyG7uWdwVp4yKkdKRNJnaIEcuJj7B9S5R4W4mXVflLz
MS4VQ//1d1jOMl5grKybCS0Xtq7l2ltsoRQ/w4rWfZY2StELMp0LrmhzDPFGOSyW
pbxMpaXxjqbuq5AMV5a2gBixERtNYUPdyP1+mhjoXJ2YEfQTvMPV7IcXjb+cFmV+
+sDxfz1PdmCiTqfE4DL+UbFs+8UJxokjtH398v7OvPYjhurQ86s//SeEMVvCkntR
432LWK3RZOSFdb5h5FJx1mFL4C3TuFfVR6Da71F6DgPLSG0sn4qffrR+ut24EBHv
p9UF8oEqzrQaDouQ4Gq6h8KyCc1ErGujfvuggMa7rCXce0Lx/ea8xQV9STOmwNYC
agbqkpUqrCW5mhckZBLdBNoh/o4T8C4pFx0QKzPxxkAafAWt2M0NmbGLqvCM/jIu
ytAXz/Vmc7KVhAhNnNcjTATQQ1b1U/owHNDHWmQ014MYMR8WxskfIw1zdQcWeQ3S
Du6DY5WuL3SNotG3DyZQEt8gqDWZfHkF+L1E7fNZe/NmLU15AJ2v82LHjy6LrvO8
0WjQCDKSw2AvieK9VBTm69su5bYjASxbEIHqj+uujxCwhxnbWpvGq5s8h0p0CGB9
aRfoO4tkDcOlNTYYuZZxfBFYT2DTiEOykWBaxhUHiFK8UhAO04PUsgTKSy1hWxFM
21tP0ZFR0FuYfUE4ESRzsA9j5QtwIr//zFLNoPvPjvqjwILEQm6dLybG1zBwTwbB
htc1XpoY82zTeZ3ztovXHbK2eGs1Gw4bxFIo4f8x9a5z2uJL4CN/q1TzLdEFr3Df
R1CX/xhJ3pLGx6Sl3xGSEb/rtDW9qAxwEaPDLGGbSv7TQQ6dUtPBs9wi0jXgtwgY
dNvCN5jh+s2qeSmsXbSQB/oYv2StgZF4q/pAXycuMXivTNzmgwAv/CYJ1ziATUXY
JS2ir3ygjRpQKY/TUnjd2W8P8uilWYLmCv/XZPlHX2JlBr9qbAZVI8gQ+zU0O4Lo
33Dzs9/x9ZLkautbFo1trsWU7khF51ztPfbJyjp0uCUt9TRlwBS9WygySEdC+kfJ
oauBTDFz71jKyyHRzUfTOSFOActTD7oD5ApIgOfKbtm2am6BkEz5/fhxHim2Ut+n
iBCspS+eIV4AS78VG81oqvuBllFY+ZtvNaM0FHaDv6vC4RcJ65GAq2ZFALkEvWVH
lvEtxTknUFdSvh0QUwLwmBXq0JRpxP7vPcc1yv0RnCDYpMvuaqP2p/gfu/cEdQL7
jStmv5hEBYfMDeRA3CoWw93FXlH3o99/Rg50ULhHC3/3/rvrBFrHq/KIf4+OY47P
vwR1aMudQbiWW728BYpjwDd5nUiQHeimy/SiWWy1J5ROeTYtas/KIoAYosAI2W9r
noFjbNwQTAUjd0se6/8fLL3Qdr1mvbTYOOPY36XW1Jd2xI3jPbl61qxeyjLmnc5P
B+HGv2L5waGHPUY61PtJ3x7DtxiOVVLfAN1I1EqWAIkJaXy9JP1A84RaHA01Du5b
ZZQOZ+79okkME2yJ6Numy2kcn2qpshg/1xi3JsAl4FmiaLHhditTIQemfDmBzQ1Q
uHS2HriXe0V0LGtjIlT4CyTXfMCY2opg7ToC0n3Mf+gbSwYfm5tAT/+JQArEYHZk
fXP7IR2dbNHoKjf6r9dx9oCHkdaBDufetQOCGQ1ue0ei69O3bN6YGdKQxdsVa2Ch
0PUg0wh86/cHOaHcIrumNjWyWfhP4pmB7NQeJWhbf0oH9M2qv62hp5Kgfrtj2vZk
3gKB8dtOs76Meb6tN6+KS2CK8p1UyG1rFL6EZKx+zP7eGlJ8yeo0Nx6Jspy0RxY0
DHCss9u5Wl5U2SOeS51NKFmMaDwU1AiXt5fe9fBMA2aXkgGoMQJshAUbeIHqMIqo
i2yKZCANDWruyMwsdTQzOVE1Ybs9pAmJ+J07px7xBGsNrmWdWivRMAmR5uXaoKgR
ic2mEwY99EK2hK6CAfBjBqf7+0RtPeH+2LdbuEf2Vjz6shkBOZNjboqCT3u0otin
lz3Kli5MGKDFuy3eWSjm4h/WernGOcxH+dGOyhXy6GKiDfK9cTwqCRtid+CEmwXV
4dytE3XaAXmlLogT6z6hSPMSTSpi5PuNlnCP6QqI8WM93ozZpSyJLmeFZqsBujgo
ABRi0IAIK72E0G0j5sMdbzXt8HaXutI8/+SE8LqWcXmWuDN+CBDodjnkEa8hnc44
WudgKS17Pc2qZK4BWK1UVYriEKedngOItThXOE+L2lO/WKOWGuF6WxaEsBS1obAD
dmpEP1H0KV+p9uXU/fHktyX8pQY7by5/A825g9WQibHcUUH/ivv7qNXKVWbuC8w9
KDA9j1q4CfndNdWYsOhHFcDJGLdqcov5RPbp7KEWPbTKroh2nQ1A4ILg+/RR2fe9
WKro1fwcK8fbXb1WpMZc5LMOH1Pz+aJxXir2ONIYdTdWIMCsMpQnFXetzYMLfCBA
cZe4bXxLwktalO0dPV5jWWhSAE+9gLMSJoSIDlHBAwUQk1I4ocyIfFUvkP48jyfE
vWfmhRkMKWoYU8IiXBo2QZS4pcYwkg0geku8Yg+giOOqkd5L/0+kgxue2f8RHRzw
ZR0xv4ZCKtHUA+kNwS6jnSt3lZ5kAchGko2SN4k4bjnp6/Ve85lt55ffLiSZyLUO
qdmDs9+MksEbP53ATCJnluwKkF1ahzWrjaumgAasBO3H5i/4FzC9NXgDrvSgwKMg
f50zk1Y6ErUhJJrKVTDVAnfOqiAAbFh+9mimth/tkSjwNYjAFNtGwFKBLpVv7DVQ
w/uIJYGxJnBW0fbKJ5I6AhJNCUcxi4isjhrdkOSUj2Y+QFvXzjml3DIxNrbEjzqb
z4Hs1Q1dkBemW6JAiF3WZyzEFAVSzMSM2bFTPq/I6fwG9WqM3XOAOQ9Rvy5Qsw6V
6V8cN6dab+rfZwLwpPaYdbGJLAhzTeyE8ziiXXLzah+Q78oIA9FoN6OTgWCUL8k5
yDxQxjL3eNViCGLxWqk1oxuCGnabAAPwR8y9/nO62op+BfdAZheLSnWrAnrwS6lZ
2rC1Heb8LPwPMB3+DoBtodiFrVEWkw2OMZmk61QC3seIRGfcVuVHryDlKbcnnGgz
iBfYWPJY83e1S2uzGjP97JM0MwwWVRB8H5osUlsw0cSxtfXQjFdTvrIpB4h4Iaim
sQh7o5iTD0G41uhILzoWsEiwe/PpPx67OICeUBipyuhazYcq7cPwfswOlJe+2Irl
h3Ac+WKgWiP6bq3PCPnkMF5xtSHgbfL8Q7qFO8jtPynP/fLLsxNIOAaGwXZ7403Q
sqCAiiYne5S7Ka83Pyt0HoxKw7l1e5zvQvKl4VvQk9kwGLKQrhQeWax28wVn8vJD
yvmKOCgvLUP9rjF+K2D87NLpBOH4d95EDNlqEOkrs6y1Wno6gK5NIi+kssQyNNNC
65L/2/FkprMFpW5iH5reKQz8rwaHKUOdTSHKcESSnHwey4WtutU0Mvhg3yFDKiyf
tniKb8h3LJ/jPuafDpDBKLVfy9s55P4ZEQWALkU0QPETE0h27kwm7eRF+qNAXHCh
/w817q7+j09KTXJ5bQVkRNvR0s4uv08fim0a3w4msnCTyq1dRh8S45T4reXG+w9y
FEn1dPayhA+UD9ITz7kGMQ3uxTjSUh2Vz0KtTsfYBz1+2JVUqZ3ZWwb2RoQgfKz6
RnUN0+CZvLpxVNkAw+3Vs9s73QaC+NFWNUvRYRZ2ly/nYBA1uDyCgS/teUPF3pDC
7oKeeoNnHS+izdTYP9h1TItXxOR7n/JuyzvHWPbJy/ylWp9EwOkWYFJzOXC+ph8C
MtK8m/Fxms6e3JKkkP0FvCpUWjOHLr8Tv9kzPegno6HtzKhw5tPZXMpcoub0k4AM
WVxkI/UA/VbGqVydx6pndvKZanknrKcRORrLB2NPv87a3MHvJ7UhxiJSQ9BG+m5V
N4sqMW6rslucMIpZxrfjACNxXtST1l5pRVbuU+3OSXVek25dFcAHjfd1FRGPr0rZ
cCXE7d3w+sy7TdL6O52MfgvqXugBvMg+lt02oxKybGW8yI88unWp0Aqbq2hDaDJy
TPM/HWpYZkCne4uodRMOiYY+9XiP9uJoWX6EKfG/ZUZZxk7qF8tQWePW0/qIDEd5
9w1mXK6hIDoCrMLhO76ncucZSU//uD9+29OL/1a4G42Kjsbrmkw1j1jqd4ERZXTW
Hm/F8AOrkdot0O5tjViyC3a0NFOn0D847VkV1iqxJ5MTu0qJovrjdVslrYhJT28P
S0OGj+C6UGppSgCM2ibAAbP1lbduh86D/dGCviXucKyAh7xeGLDKf/n4e8J1c9Yt
CrsLS84i+mG5yiXCLCGx3xSjS7ERhhfOP5/7z51cLwIWQi3bqyqHWWbp3CJCSbpY
aXu906PPyb0GyXE9+gXljhBbQr2YXO94oN9C6b5StPtSVGeJoql90PiiTziWx4Jj
7/cnYZa38M3aOxRFvKfupxNVoBTwNuwsbiREVrpcGsJZtCJnyYGIneLHigrtdOpT
ovMYL7hX5FMtozc/GOqVZ1YGQTlWSdtBZOqT0gdsttmnGjIfIvf8zcNbbFpE7yOk
O8Ha6+oP3HuBZu8x2+umMeSML1BcC8iE/9FNRI1II4KsOLx+xg9tfZEfIQ0Kov5G
Lygufg+DONUQ+GGApZTEeFiJfP+BUg1P0Z5tTyen81Ye9CyRWY0JLCGHhU4XHRZK
8+oNSMKYndHmDbPCqEcgjUtEMG6w4WztohNtsiRre5l6B03g8XSEcz9PSxdXJASJ
vDNoJVCH/fkxOAtvkuwQJ5QiReBI5JvoX4JNImojMXDz2d9b7LtxgOi9uZ8lb9fd
1xbn73fjXi6vFISPwqhw8hsSV+gfad+WSjf6fQRyPLRFvJJQ1ycEw1MK1FYWu5Px
OyqVC4Wnr+xvQZwrxRramQy60BH9qm/l86Ieu8sVocKfKwG+cM/y1g5zwvtfhddE
lxS7HE9cW9EypMP3xVgATP7R44wtFITgTTuyjf6omF+S3Y9uXLUcmlyZJubz7cVY
OMcI10m32b0wBV553LDZYOOcknTmGXDJTDIPIUjMxCkWOC0B7bJ/t1gWQwoav12U
4h+tL5aHCLRPa26lRgYq5itJHht0NEtaEe5SVFCHNrNWi4ceGzyDhOB9l98XV8+5
TkbOaYa6EtBhFJzFAg/0HxVpwF6fsaxAQBUqvfr/QxJAJ9tCKOwGDeiAoLHvhCi0
F6/ujTWtSBxLCvGWZZ2xMBHN7GkEzycCz7kmoxQJf4i3qeJ32tADhpUourMRhD+M
U367kkhslRHRize5aadCniSd0ZVx9iYBly+7DZzo73Cx0YbO/XwmQhuCBxhMvgb0
wdkvNXMCspAIHwzCDf3mC9R/RVgHlXXmkygHawGDQaWuiLoTc6v7YE+G0Dysa+j9
tDtMbc8VqEfnGux8ICEqDse/l1jPTnbl22lNKwgVG9hjGm3uDq5O9ZfUyi65kvrC
lnuYgMRZkehK2hiVCShk4P+Dd7jHmoq3fd0tQs3RD35LjGNEizSUvyHr/NYfWP4i
3cIci2PWaUzDIctT2y53uitQFG7K0hu+abZd+uH7kDl6gWfqsxTaC/NGTYHI7sCj
+13bwuffMjjKYbuya+wpfiU8319ZwXmuUIdH9TL8Y+fmQXupPQjZqeK5fdUJxrtw
RcerTvNm/9WQ9Uvv+TuqjRqvk50Qwxr2JxSy2ioeluSlmCrTxPxg+6x5TpSwaPt/
jdDXKDNVY7m64dcuTJx72nJcaP69/+YKeo1xJvSbYymQFciGpXkhQuKIi/ag9NMK
C2MprEezl8Q4Yqhpe4PSLAPEsgip2al4j34UCROqVk16YgFELzSxM/JpRnpSVesd
i4/Jt5dlDmaIsZADKweHRe4YdpSqi2GbxcCH6xFGSv/iP0O8w6wGB9BgGT1KVEMo
zfwivj/gyFMgR9gwwI3CjYofNLKmNxtpRqb3xsPVfdEYnAnuDPgmshYLZQcb0ZY/
tlM+nMCMnNfdiDsA7OjoqSJQW9AUpB2Ekrn+5m2YFdouWV9RCZ9Eoq524e8BD4SF
H5YbC3ETCWPNdCOuUVc8cKMuGmRy49cd5MLUcjseVeFthWC+TmCE5dRJFm8mBfk5
Uqom5bujFQDdxNkZ7BedxppcXwTYMoPnIdfhHK8ncZDW10tZJkD4xFsRRNnB+iJz
8GQOJHAcR57V1IntX1dxo7YKhvdxE0PrlVVtUVkX8g+1N+u3DtjLbh2lOXzBTabE
h5H30ObcjwVKIQ+OQ/pzkYbJWTW71BcToOntBf6CZXkzMd2biCSOI77W1HXjq4Dq
Ah4ocB+A8iRrqR+UaoV5hsXsCua84ty++P+TCKLYwM7QVOK6uaNDfvvZh6leAR5W
acs6+IOAV/qL2BeyF6LMCTEUH0ETG/IDukhrO4dtc47ZOUh7FWXaUVXL0c2ii4Yj
T0whCstgu0MzqaGXG3LIOA5cxfACtql/rz9Ezk4sgyC/tBGRx1vGeo4egx5DLuIZ
uI2mP4s234eoXYqak4VZg9kgIVNuY6F47m5vs7mYokbMhd/PpjNZEtVAVi5kayME
t0f2+JAFKM95Tm8ml9s2TyDgf41Om2eyB/bqkT6OReW9jP1UjfNIZ4zRdEo/zjPO
HUYWrTMeaa9tuaW+USZd9pkjao/2cqitZaKflG+wVWpUxrSLrqFmtJvaAMek00Fj
L2jt1eN6Ns0cTjMZT7UlKWjj1xDVtDfFI66y779E+M4bglMgyEH6u/9DUIWugUwu
zj0hqSJbyrTiFm8luT95c+krBPz3hORi4cogim5jPTqcEifywjZcYKNIx0STC6bV
ZlHTj3uwOJ3CtA5hHwFC48iXgmhNQpp+LXDjTt1X3I/mGe0X+tW+IssjJdDxQXAf
ox2eCY4+xtO+fvi58Up7jm1wZafwYZG773Gfbb9OSaQlRZi6z1Q4pCkIrjgUKyzC
avdIWSxc0JgMSL/mhdVSp60XQ+ixI98GIgNvMmcsrPnNuzhzONuTiAJgsI7VlPEf
OhOZny78IeT9ki5m9/JSVlC63lWPL9R/vqWI9SejZlhVYaRrnUtufml1gJUC1dc1
3OiM0IKFyIyNuyiawD2QSBnpv3Ar3+qgxQGSX4Dx7qRhjmVBshFAT4+D/gmUzhDR
KwlaeXFDoyi9dGIieKSvSSaVmc5xYirdIkFPMwhJtcMRWuMFLt+A3cv+0UcCfTnY
UBwjNww4XpiGX3s2UAqKemHiTvOROqv5Aotk+GLVK8lWt86Fc59oRHocuOYrzEPi
fGvATo5UaFsWgdTQmKxXbsyKxikm+KohPHsgoqHppbWld2+nOYyBIgl2ketcHzY7
EiWtwqvWCCpt3qa8Vv0gM4jXypJ8o+Rz/u3vX0cEsvyjZ0lA2lT0jupbB3KfEzwy
8todcEUtQS2yyo7DGMYXJpfWD1pjNTHnfXANtR32g4WtXrTqr49y11U8oRttBHFa
9APBq0PrczVpirnOgYMoaA+9wESwYtBPE0XYBk3fvMwQQ3tfQp1UakXseCO009nq
8iYWm8cG4RPIX1sEjIkw/59NjkO5tKDatGxH/epOP65QgUoogzbd4YF1O9oYKvdb
5iIC+q0Zn4v53VvnWjRdKjk8+2ey97hxt0DT5EhqeArngBdP4m+26ABCSwpsDXRT
JtPnNUxbVHKb2c62wxy/kJEzmSgpfLKzDNmicK5u/Mzt4qAcGMoX4a7oJ0HJIwRM
f8dBixBm4kC/PIOD+SF9aKAyJVkUiEZe5lIYouEvVMT5Rnm7fjJnImgUqw8qKpcH
gINVl25bffMfZoFaTUedx3GmFn/sZNpEk/cLcJQaRCw/Ef44Pl9txzNRQ1OjbVBk
0AUeTJJ0tIz1mOLspYj6BnH9vqp1Ycc+5gzUXVhJSwafR/BZAXjGWBcG2QaovaOJ
hy9uAoTIsBLIKxctWMRSoRZnepkidmoj9P0hiDlbNWNcTowCqEE0eoilmBADyQ6N
zxkTDfpquryZU4iOUAjhqASe/9KA+OjgUrrIqt92pEpx93uuQt5WKHmhBWbjs1wo
yp4X73PJEcYXbrgaP2FSOPxlR4yoBu+6F0hicAMx8Iwq0ruT57bJxFQ1ShksE08l
GDFf6djKhE1991JshioYeYxksDTIk0nBky9bjCrFA8s17EoQzRyJh1SKG/NcXpLe
dq5mvWo+jrGVUsUMgnbax9iPoAQpSlK4WvBQFw26CmS4ESr65hNgFow72+SMYCpi
DPIrZ2UyOmNsh1cq4o9Cswdi07T5bWZ0FRnyMXSiBzkznmd/6nc/A2d0dmmLKToB
8v/fJRUPwK5xzyN628Qrm4mAZVnMWHazbBwnzxG1081VwuYtU9VHL93yu409YeFy
rNpsT7oG/JlTBQt7CiAhmR9FEIcANGka0G99nQ74n6vVnhvJBIB/2ZbjUj03J0bg
kc6XO0F8nwsL+qwN2YiWBcE3ijh/fksxKq+C+wNvXx60wiSEwPJcSSVc637u0j5Y
2gHtl38+bQkjB8EjSBqTB5Dra2Yp05Q7YVv+k4wstXQQvULdzHxqhNXe6+0iIrqD
qThF9SlhBfGJYUA+iFL6UIhv7gk51MvRwhfUoJxzRyduNWpBVldcOru/qNh1lTzr
i8mVpn5hlHCsNsdpJD8Pepj1XLh2le+Rqug2x+fMLuMzD8Z+GFRhhy0V3FVV3dnG
0HKTzJzUY1eYNVT7oHoPnzO/m6xs3HgAVi8GDOSvgLe1N5ovndVKULWlylJeyrAx
TBJdNxBzkYvObA4xUr1utb/hSCS3YrKCDuWJqzU6l+r+wTl0ZQHO6OcR4yyV61fQ
Fkf4kvjNqq6TV2qiYXJoaapnbrpxW0Pi4sV1fywcE7Sm1a7B0m3Eu5otB9n4LXwN
1c/RBYwfZ6swVVeVddhdqwBgVqb9SfRbyXO/S24ceDLDKC6DCWopiN3i8UxSlShH
UMa25YQm4En7BnpxMHi/wmkHKYxmgHlHNIiQj+MmCicnt/UHTWKhCl4SktV74iSw
ay0ZFp5/56cbkMPCJ09fy7vCne2SGpTd0M8aqvqp/plL+c6xGh037+6OCDy6ShA6
EFNwqVzqU2O1Xuccj39UJyKah5UCk069rh89POJgwnPA+0H8bGh91Hnlvprekzni
Ee8FhE2mGOs3sBrARz1P4+0lc/E+z0GVCRkxJs2wCE1lcT+Su3+uWGfumDJK8OYn
C4yXhHnWiFTEZ5jLCEPS4Ai0wyNR93xTRI7RiEHxCnIuPq9Bb0C//oRwx6bKQbZ1
ksDK64PmsNDwrTiQJFERqUA8wApKc5WqIrtWzp8EMk244xF1Sce68wB+sPlB3bzz
NxwLGvmlAHJrk2zAbwi2PNdc3gA8IXcb2Gs0S/Xm4vVRg4PjbBglpCProcMApKjg
rSFEtXJKTpf3l9VxizH81w+EhdfHbUe+QG/HvywCo1uiZHx4ItCwFn3nU0sXewPb
3fmNe67fgjJxeQ4loTcFJoPKoF3j8S7uixYaOSp5LO7tTc00OhI2/fZKoHbF5wGZ
wPRkx53oLrQNdra0/ylG8revZx9FDDXObXDIg7quubZ5lIOcKnZYQvJi1R/lqZj8
RV/+EdzQBGdm5skfcoL62KOdS3HAFIAaEF92AiPGuwobfdRTTvQs9WSVI9Ehlkb5
kaUFqFXqtVnUjufJTmfcm7U0oERmuPSv33EK64NZL8AUHewSwEcvNdcn4VXBswyR
VhzwQ08ndrPa/3oz62WpuL5YQVCGcQx7nwXAqhEVXlDkbj/OV7fUuzzT4BWBQ90r
AcXxPU8TyzHpT69VmF7akZAOZVxX/6nyjGW3PMeEoBsFF37344u6mSCztx42xo5P
TrGL+EYpLxWG1BWPvSM72ann7I9CTLpc/hMDDNAhi+XWFnDnhLpr0Pm3iDLZY9ph
9gjRxdAG8o0hCdYleZYvmqtCF2x1G5ndnON9ndTxLpOxysd4geTItNn2Vy3N3MXy
9kFIrVLme1+W9nJ8e+7j4wBR8lE6yO0mwbyUdevjQsiL1auSyCdBBgTGEnRn740v
RE4aQFZXpnfUA2CEbgllRPfwyuQcDqWK2QLZRRbAmo+8s2Hjdmt7HOR9RX5COdNB
4b2l7psqT8BPeSSUXQGlcLqCLFnVADmErm/K4mSVcmYRpzI63pFSnBfYgr0DDnzc
TwDqmseJAs6lOB7701cfAi/6cyf+FD9dPBNyVYXrubj8FPQu++Xh4dtVOKI9F8HB
OPY/BaT8C2JvnB8LvDomFchdLB+8u+1j9jOzsIE4U1/tu4HUlKEHwj2PUMNYRURd
nRS+fNo3T/bk8YUwhaQU3SmqpxLUfcewM4WDeT49nttx340sR6sMmP52dcvWKR/C
jg5bigWcmDAl2jC8vI4iC/XyJzpJQ4XWINo5jrqf2tz/oUjIptpCTIA103vgkIu8
GMqEZTNYv0XFPnIv4zkWGxlXAwsLBbPWht8M3k9DjSMi1XEm04imNGOdf/OxyyQF
+8CtqLBFqZvht1uMeSeKt5P1fjWTkH1EwTASO9HxMeLWdAxU7y2EYQJxWWVzoVdo
p0odzl/gwqhZUDA31x8z0MMxbG1VGhFHxPwRQUcKktSQjaGotCs5z9d7VYWqjqzh
d3xUzwuMOJsf5t8njdaDDGSN6oaO9CCfNeMxmlHq1kBCVi71NkRglXNQNmGGdpiB
rdwgZK5KohCA5KpPUrdEh5wU04uchP9rDW0fcatwabp0w90sEb88WG5sI96DRkaE
vcCb0sjKMgAcA9RB3ldv4A+W0subV/KtswpdpSRT0q06iFJVvyVDtUu++uZMBSrg
IAQG6hjbhwhCH9sEyXCP2pP6nAgPEloAkWQuBdfLsBB0n3lWlDzvjIYFaxeXTYBi
uwCBASPQgwL3HPZYq5qdsHmzs4MicpvIoG6mIudtXAoEAN5DRsNZLjiHrfiLC+sh
XRi7lP2eggcsXYj07OfkO280MGjcu0DRTRSAlcrANElsT1qF6N3UnSULyw32cA0G
ZFMTWKoU4kZHDmEOIEYSRV4+/h5ng527MTdvEEiHXDO6cMRc/d5ACTNiMRpbYhRF
85e5RpBIbvPN6KvJdFQphTCFIPGMpX+dvDBD69Z/6ITJSc/rKheKDvf8lP762dW7
sRbCu/2AXjc0GK8Wc9ezs40ryJfCLhqtN64K6Ksf6TSEAj03Th4dbf1TYms54KZs
VpfBei5W55A6BVcBFzTEutuJw1lE69IUTjz9iUXgUc1pea2Ce13iCElc6MS00HWm
YPgGOWSvxuN2769QdkZ2rHwLLf8tii0HEGDUQ+iQK587rHM2ITHIspEbc+3DIk2A
4rBKgb+bmL+73yUyG6nz2P7MmD9Hv1IDSqUQ90K8W95NDqXrMnXDwmawmtBaKd8v
I0l48jhvlwK0Hs0d2BDUtelyTKGizpO4LtbOQNiO/s3SarG6ouB8DMAaK98cH1eX
Kta60MfTd1flQVV3QTWBGIu4PPABo3NrZtGKU7A6kdlCOGJMINeOcg44FOTI3M9Y
9KMNl+FtlfMADe14LIKpIbyQNFyA40HaVFiiGRv1PhKBzrvVomqAvIZfHHYU6NN1
XgMeOfxjgQK+Ng6myQ6gbxuyt6e/cvgM/g8VKMgtNUstPdJmyHG55BCdkBhbdHlY
Zd/J7fbuY2QWVtfU3D1nPaQaLZZmDN09rFgTx6zaeVgHpkOkqsekEJcRgRSKVND9
2LAiXcsBD1b0JVt3Rej+BIY0zyjSsQr7gkrxxfyaEviLUNrfAWpOdPcEPQP4Sqlr
Trpyd1Lj1WNG/uPbeL86X+V3znjjPsKNUvzwHA8FjrckewSMqMq2zE980DxQ21cl
fmIAdc3GUjR5t7RG9vAKwR0LzVeDrqC7RuoSJxFKRaZnL67NHDnW779Q0UFccrLR
PxV+FgAmjlbsL18cgicIO6JA/oVaH1+HyI29eIw4BySHZEPNRlILEEfTpP/spiMG
EiJfhQ4VIVyDBJs33G2VkNmSF9L+lo2S94mzh+8FEGuFWcPAoBG1sdUee5VG09Jz
z4W9lqVrGtH26eqS3RLtsIjNmHsw7jJ8r0sscHRNq6vrP1fhUEWCRDo5TLz5HNyW
Dekyf+K6o4sgV8zvAullCcFl9D9zj6v+nkjTOrJI6lxDV/HmwNlYTuC/JlYZkuMs
+NBwiqJ8mxCAKHcFOMNOpbIjx14Ma4ca2Bn+IMnqFyWchtiBV/SvoYUZf4JljcBZ
3W2pApvkm3UUxlf08nAetGGMYKjBaV+xwyT9zJjYSspQhGucwhjfmfHRPJoUbD4n
wzNb8iu9yzRhb9Ji0S8SWb5/EoWcnAr7CuPYaqG5c019j2L1urEIU76fbGystWGV
KMUyWNflrCSITtvUPOEM+FD33wxsvcMWmQHsJZpD5JI=
`pragma protect end_protected
