// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mJWmSObx6tQskw159lhQVDMfH+t7LUZ2iUQ+iYodJTTYw6X+4QpN0mMJafIxq3CH
yYSr/cYLBHgFOC+MsrQsQjRPIX8c9HDxYOQUIvgYiYAP+Jc7lqSq4i7sOoqwtZLh
r9l9kK3Id4cW3sv/M4u4SCLL89lEkI4nD8zkl/Wza4k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27600)
Lcg4b7hQDe+aKBT0KXn9DzYWExvokTAMKk4tiuNa/ymDtWvQ+UjpF72ImJTDYu/b
Sf9XP77lxhzH4bp3s42fqLR9xJ1pJgcrcPCYB6anrS08RQ13HzqLa6N8L6QzW7pt
dwrT6YeaN0R7O14ZcdyUpOIg6Qq/U6eY8eCJFJaWVOXVaFoo4LAX/SHqjbvZXwDc
6LaNiDYmdw/4V5Siu4ofhcblIOLM0Lngz3Ek14jnrjZggxJYs2H6bioZU6WOqrsd
ZgjpoW7q5jYfZ3nuanXNHyxjlKR66PUob8fnnTEhsalUgJEHE+W8rAACV26+siWy
Z6EqTiUtwjhmTpc1SZZlh4IKmwGiixg7omGnBmVLXPmb3jjtueJg0te19q2+2F9P
ONc7lkM56RS/mku156wFqXx63gk+7MZztiINzVWtZG79dCZEtGYPAiVrIFPcoTlg
zYiW0M5vXTjAudBfCiUNQ5jPbE/X80vcnrSgLHDWv4gBAuipQ2Mcwj0wXFhuel4c
gA/Jd0s941bw+CF+qaUws4BEL7AT4+mgjZ0+UjS/5GP3tsIGBc5QBh3VE65vaHmU
5Jn2ndZtUJLr1fHBJFYJJuYwSley3fbIZkPrkIDD11yyR7meZcy6IxsTT3ujVDa/
Nn9VBxUHTZRVLsTooY+l3eBVCMXoRcNYx3kWaZ5LBJwxh+T/sz96P2RFTI39Nslk
AUF66WbRmrlhH/ZlTbUs8n/JX/mNAAcL1HiVs0rkQqBb4k3IpaVFgzvxXThIGx/A
/d0RLW7x4OkkzYK4egQTUkDnsNjA8uy7dRrtRx8Vt7PHzL8GHT4ZXockfN2zpOdJ
Xefv/jsKcEhda98ZbsAxtd0faE7olcCgozHKYPxmIRa0rsrv0Kc9W3HPO3uhE3gw
mYyS5QEXQDJQpXEWcQD/vR6tVPDJ9/aE+ER3YQRfZn+Szdmsve6yTmBbQ8kKtDzd
CLjMPUuKECTQatIJ9Anp3AaDErMHSo4PvMCbv9gBuP+AwR7bqyt2PS06I5FVHj2N
pn9cyAi8dTZ6nFEn5x5NL6yI0+n1VApBdBLQTvgvFzDJnnbE9UHR27W4TzAA6jzJ
Q/KotEFk+YXA9Z9xZVlXRYTpcRQX/ov6lh8zB8NHi9wopRFrKi9VvrpRYtJuPqes
FG3v3zENvNXuXO2tPOhOufVqUtTg/L5VnY0QseVVvPOdGAiO9ahA1Y7K+FAm6CTy
2ne1vm5dsbSTh9CbFsK0c0rULGsx2cVnKV4wK3quQikI2mSHLyooGLXuJI07YEUE
3dO7mJawVK5/9LENyOx95Y0XIvtACY5WNmnMG/p9lCqm9oAb+4mz1+y8nVLCoJOz
kfdEh81xZ5ATFNwHwz4GcFWMsTm2h78DTOemfMyX+Vbo36e8j9ju8Po0euyEUPTc
eXzI0Fn/rnqr0DeMYrhk+FB20s0jx0SQKG+gpKGcsdxWxfbosmUydnCupZRmsR50
5rPaGFeu7oZCNu1qja7wjkCyJR9te9b5yDmCPgvR3UL6xawzMwJni4nz/ShwW2CZ
YmstzweNsNLGbhcpTZlm1BCP6+J3JDc/YmqHtAbiulpOvTCY5ZN4sRLcDmhgocCD
OsFqVgVAqiEOf5S3S8U1AEhz03Cq6Lw74/UnFyVBVONTM3RviCdUddk7RaL0FxHS
mbeqB0uMpQ6pi0xnOEvXABlDGCDk+MizeyKixAnezQ8QINv27AZMKQbQKxShJEua
p8++Ngbyg1oF2mhpnSi5KMS+JynJuQvNzURbdeAyBjWZRxwWTSovHnMPNVhjcDQE
SMqMK3bhRdWIwzpfy1QyMtq3q1KMoVQVZeNe182fSxErav6Pjx91JYloMSmml/US
b/ApTyTrqy7yfbvzK5JRgwb0DGALXH6WSyAVOu4a2peK63Rp2sjZxopCT9T2Iyog
aEHV8Jki5jE49fYhi5fVkPIrDJUj6x9qpwFEUOLrhZkkdhSA5H0SZBd6GW6xpemj
bf63xrk4FmA2fAbzV2H9sHjOlMpXPThXfwSkrvYITJr9tOciSk2Q00Fd+EiYNZTW
MEJlbk3ezav7B3y8I2FR696YzShGoTe851vHuc6zx2yVEDXw+lK91L7qcvn4MCxe
qvpO8/IKevRZ8LM/hZx/6ylrLM4CG3ldgFsWGddlHkc3xCyupXcN6ntAzGKODI8Y
1Skob43RCvVlG/v1SOrf7AjPTSvl0ctKwWN+Lqs9+oloD0g9+2skTu8xtFsJ8aGO
N6FG+efUzz/G9rCFbBiwFQZIVGFojCtuNPCsgHjdYxjlxWOZ1ZWKEp2Hscd3UaZ+
0JgkgyZaX8mT9dVJb2vzN0ahk5ihi8xpESH6KrUJLo7hH50Hp9L4HnH+X9MXmpot
F75ULdoCZC7ylhy2BWWNrY3NnQWVwiQ4ShSYdijEowgRnkDJiOg5UI+LrvQvyO+H
VQhMsaNMl0QdhI9r6O3dadwDBbJ6TfoB6y2rcnQD0UjVQcZXhISlOLPi7lDSPwEx
dqgfGGX1nzWyBhOyxYWjeKXAxsyps2zOjZYxrkKUAaCBLdJFi+jc7ia6BIRevA/V
Djg01gR6oBYnmg+eJdAFY8sZBtWKeQ2thzvEZqp8nuI+ruO9pmB+P7iqAy4tokni
14WSChH2tFAJmbdiYsqLHMIULwU5W/bZu5/dX2Eufdn/WSnM19mKjm4CiRtEoyc9
xFGJ5dMs22+kOteEAgGVoWSWL4by6blVDn3ZaATIqzrDFAboL7P0nXIiEY2/z5A+
lO0l7s42I99bSFMb2teld077Cx2S5XTIFHRLGYoSnYZ0Zb/mDvXbiQs8wotcpLbu
yYOUfMItIJffasA/e/+H+V2feWTIP2ddHcFTMMp8IZ3DscPfdsX1fotsConJGPjk
acsWIHrks/tHuwe30NcnEke2WQ5uEuSFFQefjdookV+lwzKEq//qzeQ3Sz9D9CWO
l8wni7mSjyf85co+2tgppiTYf88CXcHZVvHRHkh1voyV2ixTd3/4Hr3hqly5Skol
AF4AyxPW168Lj+3jJTZPrUriPrawuZYWnVXKTExHLHS1d4dxHzYtkyNt36mQguwi
aPHS4UQmjZIZbkz3wunGynJwFWiP77JSxtEcIu8t5P6/fGQwpe3KQNVcqg7Qog+y
C9O7SVzuV2lCX8jQw9Mvv9WfJXBbp4JFP+h3FmxWJ6CEIEZIqBWe13OscllmEFiT
sFztbfrthgsGdRio1dYs/fNViqoVvyxieFNSw6Yj/x+4Sl/XgUfNIdETEk38af5h
YaJtk0modmYeEgj5mhEwdaKmXgcvYqrlMbAKmoOEgaMOgElwQDVWgZvOX++DN7Sw
m9ppooUYvOdbiieGJ/23MRWPG7Cn0Ii2lG5B6q1rPpQeEkYy2Z73wI6Ho8FE9UU8
5hpWjrHJZUf/rfFMOigeK3IRYr9bdSuhWwIzMboYiTDaFCAixsRown5S6KVE94vK
Up2PFz53dHOXADsj3le5Z6DGFrwBZuIqTSveON7rkJ+xCoNL6WPpZhAexAlWeGyZ
yJUJC+6p1kBkmclcytRY1tsv1/mlVWYxyRQLozL7aoVlnywPaols10B9IZQz4xi2
1If0mSLiSmLhwWA+qai1WtU+UixA1npeUz/CGUHDrz8XkE4fq3QICY7WQnUoN/rd
/B/aoXcd1KGruWwMQzacVwaBgpoJh4eohlIAciy4CusowHvGIJoy3R7lnCNbVNMZ
SmPfZe3KSlYbeYQ4srXx4W/JSOwatqYwhaKEylVjWR0cnOFwcfq/1gRDAjQtmu/2
RrgDlPFjOkuiLuYtg5spA4jpFBrdF2D2jsMNmShIFh+oNG3PQ+1s7WJVMr2CXt7p
aXfJ9ZzmOORWRe16XUT77TdNN3FFJpaROxRKvUFvDO2spgzpnh5Sclybrvef5DuG
BFONbMI6MUTxywmYED+/i7y6KUCH47D3co0ahIN1Z5ia/G9CyfHVW3MHAHtMqJmk
/en8+8xULIAkehOKUDUt5lnTQJ6+v7EG1Rz3VaTyFxy1svh/Ek9XB61bGUpAYNn6
hUKYabB0S31y54ZnVS0kRgeCOLyls1M/qUAaUcbkEd4kLZ8e9BtVm+ezUkGHVOrT
tirDfo1nzYDw76dEmoYfGJfMXDYz4DRLZnNh0kJAOuMQCas4ICOyfFysNn3ARWrZ
QaFN1FM9ctmTte35iANy1vD052kecmKEMYPc8+E+h3t1kDuYatPA+0kawxraTcsV
0j/NDM2m8LeVLndroIIX28CoEwbjgsl2TPTmnFqtAo8OaxKOi7JmuhFMoL9UDmMI
Jtqg0SYtDeOXRAnuVpLx7lF48Y2x9Y13Hlj0VlPrkTipc29M5osyt8HEH9JibEEC
NNVZvZeX4DjsypM1FI0nWlZ6WNFSBa+jkHnlNHbByF17ZOvKMvDqeON/wQSGzfzq
CMw054XC6RRmvrrB8+GbSp6/8OfUXI4Lhw3Fj2Ro0IQwC0JPHtM6LDx9ET+tOh0v
V4F2LtwogoA6LQmZzrB3q2R9LgRE0KLD6NDRP7+oVbm1zB/biNkI5G7+1MQZl/Bg
0hpF9kqxH1ZNnmYWJVieq+VzypiS+EbQ1syTqeKSp2vhUjQ/OU48hjvPQS6IP8qv
Zdqm0wLKsjqL4LVm55i6izj8FnwcpGfyNUT/K2nzPVAqz34qw2tyYguyPCikYV7Y
hfddn80/ZR9TXKTdPLFLuqD6IokLPrs09zXThS1IRMOCfnHLYk8Lr7qahm0i6KfH
EVEW4R8tB6y7x5cs7vz8tT8Uoi8eslf8xw6elApSTzblDg4DliHZM4113u44Wcg+
9zqcWBnirXBoNzRB5qYE7a1tnJCaOT17zFULdwpq4ba07uk9H23xYq5i/rbe2V5j
xRtGUyxrvKp6KbtaKsnR7j/6iRR5Mwm/c6WRLqL58x7eoIweUG50L8ilw/XPMQ9Q
HMsS0mf2AFEdpWPUCd4osuSRA/Qfs7eZCxAJrJeRMgMPUWZzfKOBARZO7bTPr29m
BAEeb2Nfg4O+6cUZ5v+3MK5OdIBUeYWe9KRFLyVB4/xvqoEJi02ypiA1XuueYtdG
yW0/a7fRf5i9eicKTIcgoEFA+gZNpFJPDhG/riS3gWgylSLgwzxiu5Y8qUyezh84
h3kREneac9Hj48nNhU4aObr6pQaeC/dFsXVKB55kpo9fDtfe8NpvXhNxb+ChP20d
pkSH0gegAxBv0GG/LWJWtoTnMqr/Zq06e9RK3yli40raq6T8lyJqBNLjobjBKpao
77wkfUkv3UYel8sTLHWKkFNaqVHnbqmomM5c41LmVBZmoNV6ZhklPeqeO49sbziP
u7z+U8d9ubLIUNIyr5dJZ7J4r/GAqCIKrVW5h8uPoEiHXQ6QeJ2FIrqTRApuju41
KCdEhj2+pWZsV/w883ZpOMzz+Foi3YieDmd7RLfGWEky/4/xkk90IG5R8KXoarDn
I7czWNDP9j9sqvsl3c5DC7sXaBmsXxzF3gvaVpPgUUgl7jcl5NbK4ePIjbxZ/plX
wbFrllwxoxRseV0WtRBfKzn8y/UYLeZRJnlVpSnMRqMclACP4Al8totesAxGV98c
9jdom0S1JyUUy7RZT0q1Tvl+gQEOtR74iix/7SNj5p9XOysylqmJ96Q/UuQZ2yq5
AsFZKMy4CNuoXFHbubQHR+jU8AVosgLqzOTXflQ/43uG2kywjO4BH1qWldTQ+Hee
cRG9GL7RptGijTWEd9RapaytRUK4+iC8YSfBsjVBbfsNLUx0Y0QeIOkTrm4Xqj+f
dzHUn41FnvkGfYCYR5LTEWD4+24iKNVyz5YKmusz4gHhW+DvFirZDEqQBFeyufW8
29E2NXtI/34hgj+h5r8X0Y+WBCeWlVE41oLmIe91JJNEGTOKz5gO1IirLm8KcCCJ
hf1y0NnL66DH+5Gz/c8jzfl18FXBeZek5QjkgfL5gmSqsz7Ke9DFmdFctR4knxPX
TwjMJhqj4Z7OkUknKTv5NvfC75AKcSAi7FHWaFOW7UBhbBJLJepVRqagWaOvFs8J
+K8fwIoUatHLTrzQJeT7VP2XX5kAXiLZUDhrJdqXZs55WZW9BM0NA/9y9w84h6II
rUP4BlrR6dvb2YRoCn56Zpm7ST7IrkNfdNRlutrgiYVs2lChiRaX7i4AamYd8XFz
G5cD/q13FhphvQADJto5eKjxqj+q7sqNTlsV7siUIrclUVdWtUKJ6Nkd982b6/Lt
s0c/x7wW2vHxIGlcQsQGqzJ4X4KDPC0TIQPIvNND/4AHxu3ecEBBDbGR00SWa8HC
gUBOSUjXMHLMbNfy2o0uOIQvcKIdYfnm09VSuUO3Lt6/qsTEzug8tCZ9nXXgUqbs
YYusB+FrVVxYig5vL+qS61NwbPJHVr+mwWRhzIaEVlysgPG/yda9aDl+cWqjxQr8
3hslAIZe9c/aHF2nKCDJn0rh6Blu5YLCgfGHyS9r18I99MP0l09bk7cXD17uiaAS
xAAz1mNDCNQZbfvoEG75DRbMmJJEtDlw/gkHFDm5OxtT8RYqLZjK7RVWCoKoYcR5
glBl+dQLr7iuDqGlqwSA2NnD7VSlke2J6mwNpYm64fz7Y9PDFE0sjOVVhrws+DHm
45//tJ60VRgo/+jsOUZYLWygrJIUXThh2oiIUGY14mi42WnphqUhIFl3HhKArbZR
D8OHNd5o7EoqbzUMdJ+vuClhvRSgDeBmFE9nXTrsDPJi+knkiqcnSrfDJNoYh53Q
i9jTsJ3KF8x5PF9nl+MCELXj6G+O4ouButpZ4Q/CO90AKgF9Au7cvmnXHST3FomE
nY9TKXBScNB+fnVDmGfTO3+56t37QtPTastZo8GabSe2WWsJEmCQeOb3zNq7mLlD
UFYs10dYjHh8rquDJB+4/B7tSR+K7F8UDnQlvVLe4ZwtWNjHqGokXESyoP+OOS37
LN/T3rpwlYp8V8XlpLABbYgTNKz1korQ5zXGRbuwu8trwYoh+jTtQ5h0bDyHt1iX
p9H+qQt+mdOozrijCio4qw5AArRxYdOGCAmqgv39TS00JIQa8ujcl+sNFwZWBYMN
OsbGVKmZvikUbKrhOV2yJjk61jEEp2XvuzkHmow3EsCWKOmsbGYnv9MREljjv0wa
1TZH8Le62ogjbUN3PdblVbCrbuaI4VHsJkmbaEjfzFapLOAAZNerdlXA58t8dPnx
ELQjB5Or9wVvBxlMOAG8ppk2eOUKwGZMCOjL8nD3/sVOtlCBQXcsIMTWjOsvRpJM
F3UbC0STq+5CN8bJdg58+7JmGf+JdatDGZ+GXZOMl3xvYpnzKpBayeFU8cerSAxm
VkllF0P1pQjmgY/yUKMw1sudn93L+3pvihBeTSOocEx6qfN/dTV43h+momD/x8G2
ZclRddsWZnNpxNWJyaEs8R4kknj2v7RBd/USpFYL0/KNIEjna3Q1i+kyNjU9o1Rm
Slr6ZHCb5a1dYeoEIgRRvbvQPilfm9laclQfW42JOcWa/mTXb1DBUcPTdE3dBWmZ
O/nhenOG7/+UnC4HBzgtE2A5B1mmyFCGuzrtpDnbz02H20wlYAnyvOUVebiBYW8v
bPPsEmul9Pjg72KteB+a394Ug0gUb7K8GEqXfFSbV2RbHycZ/57z2RwdI7wT+zqt
QtruIkozpfkGA9NJLwwpDR0jTRc9qc2vHxKApDi0xLPJe6mocGRT5BkKW0MFnW+H
VVuBQQp8LRH1yRJLyfM7fHQrw/HZDbyqtnl0ccR/+U4cL2K0nyng9AfUrCZYx0Pf
DS4OIoAL1u1XaswTMQvM6J94R+czMbNjlk4cUgIuCCRACCrHUr/fZbexF20P0MGE
zCLVRITtufjNdruHzAUOvXntU84V711EFSWRqnf0GDP/jj7YU7qSExXm8PZtHA7C
MB2EeR63H3ZHzV/x8YeG2r4Z+yhZiNylm7/FeWanpRX1M9aXXSatu+lXeptysDIR
xeecMRvbUBySZZZW76cjm/27fvPrnVBP+JYBSt1vpt+qVQO1wrNp09XHRM2tNsar
K1+PiQp4udMMyQac07nyIqVM0jTdililky7gn2O7Lrdnh6D3g2vjJBXwHzKn6BxA
sD87YnBVxeZ3J6OMtEtsRs8K7t7xIG2aAop3IKfyNQ0BEE/2ycmeWn7pbWqttwBN
vqKDY5a6Ra/g9EhmfDlgLWjH/j04YF8LWUHA/elbLfEQZW7vrcJRK7wuyh22enxw
S7S8GwRrKFU7niRft2LyauClNXeNFIHSFQjoxtLDbBTedCPUYTRBBQoX4SV7DhKs
hLlDc4lW8oYh2tp3JSK8JP1PMMLfFPiQ4WFdUT6WPFON9/VBwjtUQ15Jy8jB9OKw
WBBFr8/J4LSK5Mio9riJGB9AbaP5ANi0oFL5wB4rJK5mEGS9iJ6YgVPpmOw9C58E
kbUsYoYRgIpWTrUvNKCvqmI4n0SclrgOxB1bfWR7AEWcgfKd/RRh1o6kZeirhZdq
fu1eo8DeyuNSoS7LdT21RPq9bVQeQQsQayUwula4T5rTR3+YnKIYMZf9cfk34ITN
KMeFfwnqVMYnG7nAXLm3tPiCSt4Y9PaN49FMXn4ptns0ceMLK2bvcQNtjz290gr4
jwlNJOnFcIpDGaG74M+vTim7v6hctYEhZ8Yr1zFz8m/zB7d0eGtobETmYUNeLSIK
S9hoBzOB0RgLXU+0RzFKjeAw8the/vG2KxN2i6Jrr1SzVfCBQPmbtS5XD0LverNz
A+BZ6wKrxkMphG5eI+f7BOQEt/8JtgcJ0FpqaO1WtqvkpqWXzCJUSLq7onluZKIt
dj6W569WZt9+ydKAO2WN5GbAdjHbx0xFTxRVp+ebVctJDze6htRzdY0/uTWFwZJc
f+q3szTm09GjF2VwS/Ey/DkPwBcKFq+r5PK5oY8R1lxB2K4bA3SgRH0SzQ6vLJwm
PAsvjQgOT/m82Uvjg7aVtURqb3BgN0rOP1aViImdrNbdd7YOunz5UuJIEkw3fxYU
ei2/4QGT+YYXLfittvGrv9bMUHwN/R9nHtdourqc/SN/ot61dVLqPbh5Jw/NYuWB
WbPFX9XZcXEyAeVtsG9PHTFxE1pPMPgag4gAouVpOrkU37LE8gW1haTVSdrol6bG
uQMBlSf350QzDmM6iAIP9vDLJZ775ezHSMCdwLbYyenCeKp0oi3mkelBiFYfTE3v
uX3+KQcNIgoaMchdDf7nLo3pgLIbRMU05TQI3hGbb7Ze38FgfVh3srEZalvnp8P7
WZsy4akDip2ESIdwHxDgTEKwkvc6tYhmJMlE6oDmsMFlZlTKIyEQyA7VSUBmpenD
CIf3LglTsvF42f8oheRz9YWWLrLogkXb7AlUkhEaSOHbtDWJrCKBOamvqnn6U+Ca
iSqXwo4IrV1rV3u15odieo1D6qrDK3D2B5dS+rDeZ+lVDpOJsXT7mIGBKbBpZjMx
dRa35+iORsCDlJg7xfrzOXmsrC0FNmPSl0Wpukc4uXmW7mKoHFG+9yv+DUggt2G+
r9QB8FV3g/Fotykg+ZEjaJN1QfoYWX+90vWplVdDTVTm1ENURP3PpEPj3IzMyb/L
bOLBadTDV9+hPLM0GHwGoEJz6dW5fwBuN+bd77nvuihmNokujPHAc/7batRybUhB
h1OHqtKWzBsaq1s6YOB4IDMC/Y+XcPy+fNPxTD0QelUul56ytKnI/Jx/tZCgszQO
AbtVF+e46zBKcODhrH2Rtt2WhrcCWdYHJu3ZFwD8kASrLVXtnFIs35uZBYodKv5+
tPmLQCuk1a//E5v7taGkEDj4EQcImT2/QL+i/AMR8avjqmxDjpr5HVNMqY/aAY1n
AkikzIa5OL30WCVYqMu4I6rObV0DqDDLq7JqiRg5aA9K0tFaD/Styq/nqyM18QAj
sSpU3bgUUVIpfEX3Yn9V2fpY2jk4NoqyORj4NzZURO9s5Kr62aF/sajR+jNFiR7B
ACXq215F28XyHfKXMaPOxCMzipMI5j8aK+bpfGaKG/9N9kEk7OM2wQePSTbczWO3
T3MKj47ieGT3rcaKQnz2iVnKWOsOUQOE+CXRZhyFN9N3lBKcFsqvrrbud5fd1fMK
7waNTtd8T1bcfL6qp3CFp76JA/8JghfCay3X5LULxKbaDn08N7OGIOjlXEQU6usq
ER6jPcCXb1DBEIen7C/psh70TvbSAIzqTdPB3TspfvnzAoclifqTjxpCugSkHOAO
H2WcKexclfg4yq39UzJXxgtClEP6u3oO+Bylg6uhDdMG0lX7AQYUJNk22hxNhhSd
oLBvXrEUzOYRAJMXh+IOjQ+gafo3reyuD/uWngY4fuDb5e/HG4Pudv6yVlGDMbpj
aZ9J26kHjbhGzzGamtRjo5XDxuACLo2nOuZFMa5JraKctUgN8lL/rV8pAwxEnCLW
owGJumRff0azhWeaMmbSP50ogQVjkkCo8xviB9jE54llrBNQPmtkaDNwgg3MTISS
ULqXtJLywL8BVf1YE30hADNmAUhRgTsiqa73GabTLWq8qOfvg8Bne2ba5K7Cv7dU
LNrQdeJzNd644lRnz6g0s+nPkQq+xn9+PMFqVGcYewd6bdWEYEduY6f6CC5+HOKB
5G8iiBlDePrrJrMAa9R7D3k82xNjWd5Y111LMYf2EjI3Poyd4QIr53dbPTBN8NFA
JUsCtSsIX87FDO8VoxUXwl7f2K32N1Lg+jYI1ZNvSwvjlP4tdghrpf4OSqjW+Ffp
kd1IGkeYyfufkaK0YjHsIJW75ZQniZE10t0YH4WY6NTRgwDPE1HuECv3Znh4EQ/2
x3YtwIrVHlnRVAzrKuhsUDtSiW9W1Yj4LUtVsD+2pL2hH+PYXMp7rkc09V12Blxt
3WrcM1jBZ35+gFJBBsXflVVqxBCxt9FneES1BHj21mxOHgwvIo0e5e0w9rYhWEiK
ExCezvuo6vK0GUwQ5qmPBlHG+kmkbkHexkoOWJGD0yz5WHNFxTFmUGR3NmfaN/Qu
cBKcwyZ0OZQoWDR+0upg2dBHqYAII3QQAOUDEhKc0yZ/POFtXLxw1kTonYG+l2bN
IZniaS6pGh3SY3WGKzF3OFWf/PE/Kkb5h+ea2pAftH6cX7vm9KG9O3czZKG8GiHM
qe/o2kxYm7bdDdmmGET2jzjOrAmrnVgCpcTrEVpxq2LYMkx5wloOFR5C15uRK30o
4qN0+ZzM+Q1HwlaN3rhHgOki3R+zXoisaLN9aoOapnfQgvfnYPztApe7lu1/7EpZ
fE0gybb0fZcsf/TWJ8Ql/x3aD68BxL5MqvTYxrEmF+mjK4Pl2W5EYVqByvX94Ig6
JVV3g+Ep7qg+/swLPZE1GdKJJ46M6c8iR6hsTbgBJYc6Ha4xB+bPAgirHoTzVQAT
hqVYjnVuMiDI0QKjkAM5zqkurEE3RFZSfAsyeLUGhvUIHt1GQzGYMoN39SFIb0Wu
cADpd4yzuXhUvSbQumaZBIurlIK00V5Br+TtcmeP0t6EmmcnUuBh4yxif7Gd1ebs
X9GIhLaZrvUi/fiZJSkP5g/2ZDjUwSoCmBKhcAXhL/UCEDa9mSNek4lVIilDQPjR
OslXowDv5aSY+OTgNnVWjCiWRz7mZfUNb/cPU1xFcdtzcN24ScJ+pXRF9qFxuCen
eAm5r/TwodKiDPb6Jcyi8CCr4uhtJ4D9U0qLpXRc38ljDHQtNGUVmPJP3DtLBJTa
W/qrG24hEd7hNh21MU+ilzYeZPkJjTjw9XnSYXmr/orXmD428fhJDhnGTtjVh88X
o7ZM9iERt5e9o0y6cAhUX+UMp7gBObEaPYEbK4rCFOBtWL0F6jI3qmvsRUyZ1tVm
gElRlIoG5spn/m6/vdG4eWDcxVGx41QQXO8yOCumGqFuV3cPVvQhVJQC4IBUIokh
qPOzLl4RkKsx1lDLxrm6W/dz3qgGFM92N9sBpZWirR/sAC/q7CYTLI1hbwYOHKyU
TXfDoVmoSQIPzAiqK8j/iDDnv6TZ6uL4r55dpqYJ/k86YDRVayPU3GCKpjmscyuR
RqPHbrgrBIUDa9l3KpmAZhd/ioVQNT1o9gkDhUfzxQ/qc4nlfc7yRxTOn3OeIU0Q
o+rCpFyxlib1fZhmLsujJ1ZyRlmRXMi5QSsYZaxX7lSo6gLqBymSeIDZ9FOLSswS
8o+kkpZOd99cqdihjiCwkSLnEnCqajB0Vc/XhhXVi9b0v4ZxrBN8mxcCdve9L4Eb
sOoRL+opg632y1E9afSIz9oXivAZXzVmoQDd8htlqMDTfRrLir4vap70O1LCWL3F
UtLi/HK3wIhA/MJhU+Xl+Kg9NcRDwswNin2uKge4GdpgVSH38XgkxISnb/E3Ld8m
41xf+yBqygSoP5722VLDIDRs3aioM8L6PKWqnBT/MSiFDxzQQDHqwztAUVYCjK5J
babO5kjmVL052d+w6QF4L+tqSy+EVcPliU39r4SshU6W6d6XYeYDMs+4aEeFYHLr
GOEQtEZpD7ViyJnfvUqSvxEuh+VtGxpnMfiz5BJAU9NOng53w6EPUVXLDQKIoqnv
hRp00plpzucMmJZ7KiN2SB9l4cajYjXgpZK9gCrB/gf8XnHClRSjb+k90bCepm95
0Bz4KTM1+CHN2Zwj/R9RdUsqueLyL7Il8f9gICYPrQrF+1Pe3EheeV4ToEpO+Mgw
7DwUbXP2jXyv0hl30H+3yVDRApvbXFD9Jv9ZslzK5AJmfwENyF7mUWI/cYGd053a
ZzAj0znJ9s3CQBzzawYz8Zx/iLvgoWPwuh/7Q/jYhYE6e6ETwPnNPSai8fYv/R3d
dmLz/tuocTUzp4Jc95xNvoz0sYVKp9CA+T2WQMYGqRK7cJ3tQXAC2aDdPClT2NIl
gFFAfcUw+ah8z/VhFQdPr63tfSMzI3IH7mOfWS2e+huH8olJZwpWLdaA7/YiZAdT
6hdDzduXYYGHaDmxuQfnk9ToRLhQnCX6+pLXTBMHAgilNylR+jr6krEt4EupfqsM
Jnotbcl6Nw440j734t39r3VGWkA2Xf1Vhru1kqrYqOBq72kQZRtpDNl5gnxOy14T
FJDF7ZCPA6iTgO4Yja17zyPDCXOtF2scWl71tyLpKCc/X++kWKxoiH5zsbRDUgIk
/Gkza7Lfn0nFZpDfevMmdv6FNMaiEhQsPiUQ36fiUjm12LDgq/CNNDMwUJBGluP8
OzvYAhdOxI/K7e86DXdYl6JZAhylLAXqXmssni5LRG9oTpDxXAaVa6fb7k457A6Y
pSAdMxqPQvXGKE/VsxcoBkb8PRzaeJ1Pk/G1NuduiMYF7WCD5H1hcxf4hLoa2FZ+
vY2a30grSCbOdNshZ2gBoqEuGNrfrDBMwuP/bsGUBxOqbkxSN2mrHmj0cmH/VHzs
izAGJuwIyEbH45b/k+oScAwgaQREBQY7GPw/33j3Mk1nQtVMfXHgAW6wXZ6lVpc8
eGJjNseZH3OJO1YLVOHGTP0BJl+qSdEe6wsjl6l5g4+jh0x1YrlCdyZELVJPnShr
jDAOXeuO3v/MuLkjr5EFod+H/E8vD7Qpj3MKC3HjMvD0zoGxjXfzlfAcbRvn3iU3
mR7GeinievepyJeLaZX70lBda0vGtdqAHg5u9x81n3DOQ2YXOLQNX9S9pybq+7WH
GHt/F7LhqRzIDKTbPopkUPQbwttE5J36JByuFee06qiGFMRq/L6OFRWF/yXQ9nvJ
3P/QqHXVOedKMfl8mzJnQDSUHgKnVqfLjE+PL9Az2yZsrYSnIKuOjOXIrIbIc5qt
IoAbEGacwp0Lh+7K8euq0hmDkKGmcMHa2keV0gcwbZCQn9GncgciVaAqa0uQoQXi
yhf+Gdg2uu4uKiB1H0q9pPp8yRass4AAxcEhDkpFGcinxn/UgrnRxnGmOWUy3Wnz
WpG03QV8urbr5HvdBlIBgyiNlpQ7ZLAr2mwfePYAyhN3tE4P2Ic1DIABrpeTX0/U
Aqy7wVuZaPGblVpP9H34E1YQRZkSwQsKcpUVp3LgNq8mxNDbFEE+jP6Td+arnVPR
ourB+nfk/Q/284z6axhfIvE94nZMvFl6SfZ2kjoRFL95WrIEbqVxsngIitYPB0u3
xAO7ItlxHiY7xcAgVcIqt6j8SofyAUnUNrAzNrqYsII9KZnwT9u281502MNs0LJy
PgpLZmIfqiiVKUxF6vfH6G6e2+nGvdNZAA4yu2+QnaZaGSgG30CfL3o+88ZB95H6
tjZUjHgkHdp1k3UiyUrjVJg28P2D7cfpJd1ebIr/CEwHS+CyrMio5K47SXohGto5
GHOoWf3gpfbbcIWcVnUIwiG6dU6olUHB25vuRo7+CmdqLLQY/v7xwRxnTHoUOXtP
QYu0S3snOoRyOCYThumRhwqGsgrf9TBiU5KB1oR/MfRwPp6M3QuoxdSRX0HOER6k
w7KuBN08JVncnt1lwtMBw7OpFfXHG2X/sHx+CKuduiMmLlSYSo/VuuthT3Xg1I4h
gCR+hEwLAs1yk2t+QS24NkcFs1vbmiqzOH3oEQa2Df+TdDk6TUygyUKDCERHX2Ea
EoRgnPFPfSCC3sK8NWGbw6bJFniSNgzeH1pdRjzaIPCb/xglrvke2CjOVPeniN+p
Vw0WjB89JR35DmQ22Zoh7hH67WSET6K9vi/l40bDA+Gpyo7qAAiGEtsZiB4T6TlX
h2DIlAnZ9FtkGjZtEaRa1Ja0Il4GtATgjAl84SO8NnS7D/77aLSUuJhUuxRlLqL4
xwm9j2jqvVctEBPxqVChgr6eJ5IWm99IjV24YZ8m/AZcMj39rb4ermWKfvFRPiNR
aFPsfCvuIHuFWihH4wvvb4h/mTaIUIuEQoELu0FDkBmYgJgfZVQUeInxUf6Rn0Ay
v8xI8JULjGySFt2N57jxmUAeWlZlmvteYrRJ2+7s8tbquJc/XvxrrNKLnbvB/doD
OTDADiMzu+DUH3LXnZdqliJXrgoovMZf+WlC8GdbfjbYIZ82F5gcLL54+whFT+Vd
rNzfPExpF36CoT15IeIbvZEGwbqO6W2prw+waTjWMMjrKkYZJypJCI8DVXkmc2iQ
TkZScliBwiC+bMB5m53LnfEiTQ/h7scvgUA2ZOK3eLNWIOso5VC45n0pu59OSN7a
1VYdglZ87tINngdp7MYsMqapuE19/4SuFqZU3WDbhlBJ/CKwj3bC01/Rz92hEsNn
IotJY7WRJeFValLla6q6bISxKZ9yVEkLKkmZmr7zsEIBgaSG2bNAZGL/liuh9cWJ
ZvwP/ESSIscI/jkV2xKDTNODt1ZlFBxITvd8W1XFchTiGEiFb5OEf+U8F69w+w9p
RzQx2aRLlWwRvhhhXzHW+B9YMGXdN1evzWTTx3xhS8Dkjemm9Zg+NQxh0fNMxUS6
ye3OOOI+Tn6AvGclI7L8GOF3E5m15xMsGJaJhwWkScwfQ3KxyS7brRdqL+SN8RCp
SwAHwjJIYLl0d2uxM0/cxIxSioQgNtQIALCEsZxMA6WlDPyQVTWxCxbF5mkSlX1S
XmIqvGVeL7K1x1imwAW7aLqXnGBtbWwTxdAtKZFLZL/zdXf2F6xVDXUozQbn9t2L
HUmLJFxQx9A0xhnRJAhjitDGvCrbQtiW4EqaxrupJz4ttzaBZavOK/izQubhi14I
E5dXoVnURfaW7+ivFsw1OM+ML52a4oVy897AI0WRixLbu+EyWNyBo352jMG8zkyL
7vzg/huny+Lpmzu1aNtE4unPkv/15exOXEbAtguW8ZNdTjtjNz9aRyiTzY4F9S+y
ON52WKjh7kTu1OBcPipvrXI9pkHWMllTesCdMUt6akjq6B+ueVawH1upNv2hQgnq
qHTFL6dpmYWhB8vWceepgsVcExk1sUYmTM/uMGU8b5T0iq7aXqlVuFqdSd+i5sYq
OibrPtMfQHRUxLFaC2kFzedVhq9xZ3X0enz1lLTv84+ZGp7rD7I+2f1YD4V++0QQ
w4L5PwNWkxg+Yp9bdn3cKjVSNpm/narro5tovIwob4HKkzHNCXb4Ge55yAKEBN5n
piOG4iJxX1Hvmfu31xutPGnDz1d3tvqCo6tId3bFrLvJawWdP1neMKXrb2VmveA7
rnw7daacnB4GsiWqpRdcOCNxS5eoJNiwwD07Dy8IZIgy5SWBpLuP8p8GyIzcqcTV
GHyEfs57agfWFXwGhmZGVC/P6SV19LvbPjDIBVtqmBmeGAue3pqzsaH73fTXiqKU
Y1XpBuszSBVsqUstXnikAB9epO06n8zRHTvcm1WtEgHpEZuPrYvjdGX2VlZmmpdX
aYG+FBcRO6ghu0rZCMBycKFPW/xomTU+22QILDF59GT75oyrVSyNrkXtInwsWRyo
JfrB5faa0ScGdkxvO8uuw0u4Dl7EBhm8wevt1Awsh4KkBAr6oNFL6bZcWBxvDA62
LEiUzOR40zRKI7Z/VmCAX7ZPt6tgpOL4HK4qcLNIgMNi4clh+xqNnOlUdrdXo/DO
Q/1zBu+K1G+O9jqK1j4EaksWvEQMqYh4rvIrvU3M1DARJ4A1cmudha+8nGFoAARz
4NBxFw6wRePfMz0DslnmOBzVNjID0A6aTBtY1idEybceIPejjyQ3M9JEEO8IloYq
Jn0Pnh82KdTN+xZVE4Kilpy1dsRNNk5byAstLiDAfmNI9SOmkvzV+SkCAsB0fgLq
bWMkJ9hUa3/OFt4MrLSQTdpvWoivHxX+K1bHEGCbgPuhJ3czlXEAovAvNtVs+YoY
9B0Gx17+uMM7wcrrK2p+McibPIQU7UZ9YRfzR1EOaV8PwVxOA5SkGUfAcQ1RiYdb
tjPOXyNUdQEwlkHCs956DCPYkLHQZfTdE0UOG2iN4bhI4bakxinZeI6vT2QwyymZ
3a+TWQE73wVHfpOt79pu56grygfuUW1p/jDiATzVTEdmsU1Muo6epnY4t52Z+grp
GSPCbaAsRTj/e2eb253ImOYGtMS/6jBSZHudDgB/7t1tDR5l9XJlRz96nMAnsqbl
augfAhvkkTtTwmyH+Eis1KZzk5uZQyFTViuQlaP097h3h7S90jjCWarMH+SGhtKl
8xWV98SlqWKGMFxC09a2FG82+9Tzd0S2DkyHWO++7WtRmts1Y/utLexjPrWO48E6
5BIsbdftLEnyvbmkvPIFSlQrnKiH/fKYar9yYz9FldYfsNv3kts9Qwc+hN6TkdoC
wqElYA3bNLBPf5Ff9sQFjlnZV6a50Si7AfBvL+GQ+6KKot+9idRw1/uOFPDTlWCG
eq1fDLHc+YsU1zfEcLphEPmFy1HcgXPA1402IXNpcw+U7ZWUws/HWTAaWg4eGV0c
L7uG3Lt06sAe1ehMgGphsORQO/FUxqiNEInNICzWGv9tDPil/wuUdO611Kh3jCy9
ZoAEfbxSQsY9SIV68vVVwAnZVqvbe9WwYPywqo5H9CH9HJ/hJUz7flH89AXqJMcM
GiInObLEsI3eyfVdEs5Njnrg/ZSgCGqAGUFpfQhYcQWKkYaHFU1O3pHiXWg1gELM
U4cY7gbXJc+WaVap6SCtVxKyokFaaOI3N0iCQQ2ZM8aqCgYpn/7mFOdHJkrM2rFt
XRtg4n4OgW3YRYCShty79Kjp/1Jg2cKsvIIKbDIMR2dpAQFHnzZdvoJviGGSf6Vs
odfrRb/RMEnIHngNRuj2VpNpPNXCeQGXdruQTTWLAPzyQ+c3abQbZ6baiB+FoLnx
XRHS0jkLepuWltT+4ljQPRzCHac604ua/uLW8XDGAs/tA7CxF5FCPldD4ZZzcWHM
a8hW0FiBP2bsUvTMd3ON25VzV0J1yKk542U9ZMEL4AZCdyyc0o+1n01HrDRmA7ih
4MYESUZarGAFAb0tsc5uhnre4MHSEjQfgtyaRyDDcI/gsvXw5zrHhmxgwKpSlYZW
D8PuhQlLVzlpTAESoOw3i9ER6sTILHr6ltLajMpOhI0dQh7so2mWM5rdXjMFOoh3
KPodv8Xjkkp6+ICZQrZ+Ft4p2FFo/FqwRzbb+5w/PIhyysVDcU9naGwBafD0vykZ
EBayhVRhC9OE+ZaEfA1ohD/BLiT0UPSUxpBhQY/U/4P8hvwOmheT43RhR5ag+cjA
drh1kgnUFN0EB1GzW4+yyQaSCWTO2BHfyl1kgZhhKUOWKgdiwuThZK728G29d9IU
FkiKi8lvVb1NuX7EKe0Cbko731L0N/oKuVQvHUv5pQD/M2d35aNXxnY5Gh7lvPLb
Ib+On4uPwll9tGXmjM7eURZQ9CNs4QLUAgAEeI58T0L+vqIfWdpAuWB4WHdhzlj9
yCOBwe3GZ9CF2NqUk8XVKirgCU05fMplCkAF6smcDNGVZ0KTivYRIkG7XGPSLPHV
S8KGsiAvA4VAHoVKuFqUe+sA68HL4AHWUVr0bNuoYDuJ4/cmcBJ0fhCRbv2FBRVo
NoaocyErzVJn5D+GciwP6oscEhftxe7dzIY85fBfewTQqtCoPRBVl6VO9Wf6eZtW
mSpk62s7EsAU/BhvJpycPgsU5HsT2ZnHD/3xRDE3lxZCnACBjjZSlWMA5xRUv8sF
sH4y0x4NLNGwuWnBcqGmjEgcV6QzD96PdmUKU2oWpuEntjcZhFH2txqYPYLYZ2H3
1Q3A/N8b+dbAadFVqM9Nu4bj1POqIR3Gcn6VPxmvuiDYWoI1roa+CQ+PAk46PPKY
mJJoqbswsq5QLC7zviKb1fiHHesbF4iuic/df37TxVS8qKt4S3ZzUa0OaqiPkJEO
92pSGaLMw7UF6D33MX2D9nv/qNpvb9NmLIi6KchjqgcsiCC/RjW6XywFzxmNLORQ
BRhUYQ0nTKD+wdNhQY4DFy9c9Bu0Ez+gxmzlgF/qtjbexv/o5abJHBAfKsO/bhrR
9JGbbjbX4SC0odlpy0gKUWJZ4XgSzrvrjyM8BEHujVdr/OXUbZtgmU78/7VnffYg
OQPkHKIKinLlfIhRiOwC7S9HM35ELVkZq5nUj7SsKMjQfxhmbLDr+82K0P9SII64
91wpl0e7liDa7KhLyApr3PRfiXczkJelIZaIHJDQR3YiSH6Bc0FM7Tl3R5sPKffQ
4SKbOrRPW8YRvDG2jsGFai2N0EVH+fHbeh/ZWMPtUBVpkJLIM2L3Lxzwd5tD+7Lt
EXnV8Y+pAhIx6jQU+sjTfcxud+KvGlvwt3gvFLQ03XPGC17mPFPucOa6bB+Z77se
K81n7LwEBNhZl/2wuOiAiSa67f147BebWDQ+vloj090cmYxDqqQ5eQZofbQUaAxj
4xmbLT5xR/TkyrE0FOYhyl/NKCOYx97rv3ASMBbrjUabhnFlilVdU9ECpyV/YC2j
HH6lvolS2sn+PvpT9wJzywY9dQLFpIgUrstWR+hDApDHU//NHHiOiP9gS8uG5Ei4
eLlvb42STc+TW1MSrrvEPpQ57YNJ0rbVtZ49rYfZq+iF5xy49UkAccyM7wbu1+cl
vED8U7e9TmhEHgRPn0I8lvffsla8JRJI60meW6hpiPOQ43VdtCfrIUe9iVetzyk7
jGOqJGad8qIpapD15YAVMG3qGfxN1UVKse2mkfqNIe6uJfEU2ehtsdQuT4k3QqQ2
M84fKH1T7fzUJMgnG+o1YLoJTrb6jtfuR6jAUu9bxoxa2F/DkSi6Mpwkl2/Jdo3x
KKcmBVczoWpDBvFWnjY9VOLNO+aYZTFjjr6+FT+Ml42fIfF9L9BeUoI8JUB7mzBU
gKHGyLco4xMrLUpNsqzG8y330HMVE/Ve18LvTfMcTgcM8Y1wrMk9NTIx6H/9nThQ
paldwjMiR6HQNuBI3FPRG7bzaWQ3QEMnJ8cmZHMLS0Gh4HeLRraPin8sIlLELlAn
TT/670VLgUeXqNzknhLdU85TRuCyEQQ3Sx+1+aHovAFBfSwL1myXHEMCiQqjKftz
G9+t3Guoo9alX/xUYsMqSDk5b+Y6f7XRyHcRVz/8+Nb/XyHvrjur+szvBJOlR3fO
tEOIFBzk8AUgLSZVUUyDTz0VbEnfMlJ5KeI5pse4+TRnj7MWqNAYI6ju7L/GKq6t
obkyQ1wSIxntYD1+gl58oAXfLdeAR0U/sXcT/RNqAt7Lqv+C8itdDHb12QgvAZan
NaYhOTnc7kKHZvrQmVkZ2s/JjWJ4TZU06qY0rJ7itqLmwxehTkV73fccX/ry5ZFK
2D0Zk2ws5fPkOLRekFB8gw4kKhfxTj8YFT8AI7rbqwlcK8xDE4GYtMcAGNesGkfM
yHitjxxDbPsTzZn44pbzgn00UF7aV+khrGY0Cm/z2jJkn3xacdhBrRomgreP4cbY
mir/cY0DuD4UuClHhBqCsdsN7MOg+cMwqlJu5H5XQy+BMi6RZRbHqUrDWKxFAUjI
qncH3A7uh/RDguThbhelt/DP5L/ogSdIKH7ne9DMG54hSDev+k/WdZp56sYqJN7j
9ndr1L8W4jFEa00xY8ZfGWpaMO139unDByLFa5vERD+PDE6yjjq/70d3vPNE9nVK
JoEwWE5WZH7IS3w5vdSdc3TT5MkshSmG65tDBq/TDZN60nUEB730+T9HxPpZ+/C6
JeO9fqrY6HNYKtccK4cwP33K3LmwTbrC/XOogahFqHMmkuRrVfOdmLtPWGM/wpNO
J5tI/6UWIclHh5aGp7OCSBaIOxnJn4ElPgj+cdyXCTLMs/umIf75niRJsCiHuvV6
x3dkg40VatdVrByLZ1Bh3/x2X4Rul+mcHtI71DQHpXCt6rlooLyz8R1pYIQtibte
D9hqBGDnGTMLco1wY/jeDQ7KG2VDQYgZHP82JBlWKwC8muWFicfegujNwI/GjYNz
GfSokBzHF8SkQOFDc8w6+anLu20mn4Xk6rUhN9+iFLnVCvh12RUCznRHS2agJQVl
q0g8kzKtmwwcswKDtR0XyV6PQKfFl86CY5NgSI9LXvSIt3hnxGXOJuAqySssFW28
JnPDFneX32cWTlvlRA48pHcQLX0lFqtzjky05n+s4llIzomjeUH4z7A0ULbpFtO4
567Ah2C8EAUJ2c/pbKIro51YDR292fMrLqQg0/uafExb/TVijxoUBSJl8syP92uf
IKqHLq+DMQ0+m9OJA2NjfMmK5YFocNiiOkoiNTuNj36vhgTZuWjzJY695UQlxDSk
Kge1Nq3/tCRi+ZhlR+/thuhvpigT1LMJsWc6eKcbOY85V6D+TceUCGNeS0rGoqAs
ZPDHqLba9ZZiIINKa9XGJKlrI155jWUZkyoqb+01RSzKky4P4lYK49SEbDuWDaXs
MTBpY31ZMKddr46ykSix/WyUecYmF3lFLq5TlcEDn6nbGpzDg7l4uW1FQjWhSkR2
h1qiP49ySe+jLwCWsLtQ2SrK12nZbz+SyLxFG1htRjqVr8g6Z/lVtuZDsFA5GwtQ
B22D6rCV+8YO3PZyV5HFfE/cyKrYhmeNt6YiFJ7MP4trBwWzLvMITxr+4VMt1Z8s
+nEm8Rjz1Yr1Svl8Enpqr6CUdVS2eWrXcuvXnyIhsyG572AJBqCIQMz+grTP3KB0
lffgTIm4rCQuYtO/Wf8hYnVxopVHGtIgDl6PENiYCzAP7wMOCgfqRVxAeaGFjC/o
cC++MVPmU1TVYWEsPa3X6N4rLo2TqJKpkz8jkBa2UhuLkwUTBsaxsF7MZ8/8N7dY
P7HyKS4mHe5Q9NpKEKYdHdneR8Ca0ID38ntV2y8Jf6BoEyOBsEaQaS56l5CMMo9r
bsl2RWZh7wzh4i8FXml9H9KD5+eOwXE6rP2TjauZ6D4X+ECzG2P6007PEth56dfV
ozgjUFNnYrDPNxUHxnTw8MsxKrQzsG56LHddDFpr9qjSmGuIZh+lZ2IIN1nbn1Ua
BeXFRAxM/Qyt9aBFcQNY4ftPDGL4n+z+Xog4PJPs19kbXojGaxm7xH4ORnrpPgE5
M5eJCkv99ru/TTmloUtt/P0w+mFD7c6SbZnBQ6Z3VqibezgIGP+9vzUuQAYQSCVz
ceJE7xEgSUFJabbJHfnDLTa+2QlWjfsG974H0pOjAGCvLtQ8/pShxp4WKx8odYIv
LQ5R2roq4NAVQMGXghgnfGdHeSF1D3UeuyTJV5WZBgPTtmjNlufRTaMMAgavj8SM
qrY0OTldMhUeCFcZGfYGKKBeOvpP2L+gWVKrnnP4zJHeULzOLlUlTSJA3qfZufkU
q76SKYuOdM5KqehgOmz/3rLb6Mt30OGuWFEFTeW01xlaiF554tfz88ERMs8fL2Ea
Qavoo5xTTWogWnQfFj/dm+hbu/z+YWMM8TWi5Lr5ndkl22PLmV6GijIYU+iLi5Oq
KIC1AkR4YoE33FkG5TGHBKIKrOUtwlIaeGk41ZhyWO5XWhG5u4pYgcqfcUa6YJK/
rolZm4YOvNWIm4w59zHXCVzPf7zQyxCWpXF8ES0+NwJEkljCm7id22tox8xXATAe
gURkdZ/D6GE0UneP8RyQ8ErZsQ5nDjNlmr8k5p7hDQTHZIjtOujWT3bFIUm3opSr
+9AKxgAKD96LQ+sSQO+0jmYyfpEbQxY4OgHSkcVw4ATcrzs0PHPsSsWvhtmFmG3F
O8vmeu4PrPL6CGpO2exFfRB0VHa9Pg98qwy3G+hQQZmHGUOwCeReK0C0spAzR92Q
7YBNDApRk3peSrpe34ImaHv1GYuyS8Z1gv4L75GNuSQre89zON31VmlAI+d2/a/F
dgPE13RBx/cP366es6r4+9EzpgujAdRM1Q/+RhftxKNl/NMLONWhznfnHjJP7+nj
i+86ZIG3oCYQqC/FTVkwiKlWDdrERa1g06IKMXeJMlemnx0WuPRJLeeb1bRgqIRa
Fqb9JyCnJcwD/LEm3g4uEdX73ApW9XSUjRLSec6u+NXbcm96vpqewIXXHbY/wi1q
gW7eGBnjlXHakJ8nEmBdFukKXGTxXwopF2JjZTOs+GtbBmbtGgS2wDfFUzcTvbwn
0haRJTjOpF6no7fCKUE+smXDNYdpN8JgU90eaOdaRkwvBf0qFaxli9etRwWTY595
mE/YEEg41klYAW0gJs1rLbXZi30OCvGldqe5HPClH0AiNsu+uKK57Y2IsMX2awPm
otkCyL3INARh722c7/yej0uB6o5mbg7pxCX8nL9S3oZosTlsTiopZ/WaRxtJE/yO
ABY9RyUk9zmTDIwBQSs8tO3Zuz5b/U2x+rusr8c8gzdUjrFFelzUFxZEnGLQIZlk
2IS0Kjkp4QKuiDf8NP6I9wDeRpHd+aLdhhKexjUMDZZQ5wYQxgRGx1p/Q8cHvKPY
/3S1hNCpV86yqokwTca5olg5qKsKTtkoZk8fJUMU4VUBbFvVVJf2pX7rfHdgY2ac
z+aYxWfZbzNcIGPSSaRPjldJJ5n/laBkj1gcWKkOWSeau8k19bx2gu/tbu4JENzR
2Z9Fkq4XOpIR/K/8YJuZj1rtf/sddolnnx47k/afeJy/kA0Ow4+OzbWhoa4Ffjce
fpK30wfIAS8BSBXGuUrYWIp5znIkEtFnkkOeVhNOFvAWLRqF0aFgMIR8Dhpey3GS
lQbQEyREbHg1UaDK+0v7MEgKrT8mM7vQFdYyUOScs3prbo4cWR/kJEV/p+jWMKF6
lqxbQQEJ9htKjumFcmloaFKAMfMMZbsr9Ag7iFuXI8jUfMrIJZhVZFIMA+gIubEq
mXa4sNbR2G331+7DDb9OWDz6ZSu8kGfFaVVpjNdGh7kk8vKktSE5LhzRVqXpYgc/
8bicAYie7F8GcOlTJtJxsqJ+b1bXG0+QZ4eGMBv0ZYnx/PYnVsZp2Ys3At7YP5aK
BvIjQU2JQBDrGV+9i2iN0MkAFJMNrtNf+MlW1dZv8kRLrgYicxHnwIlj5QMqR6ol
TcLDfoPpgtQrWkcUihzBeMKJCsMQLEaEnHwrOU/GvrYzM/7BSVJ2ZyYbodBVvYh8
Lj0gruPTwYeHn8On3IEcZtEGn/x/u6ZszkcRzUE5s48TUseKzghiRnXryOOuHwrt
KD5g/BozzbNAUfxFH8g3HMzFJZvZUY8uLHGHAzhZGv9eHd8mEVJKD8eLdAtMktxd
c5xhXoqkSxVYwMJMQU10IN1sCFRs4nsLT0904zziT7Fxa808g6Iq9OB4CAdu80TU
GAQRQNbKHfIrOzpBcAj3U9v/ID3rN/mC2hmdsyiSPakN2goRjIxzglSUja6AJX+i
RiAx1Mof2fJywu4S5d35RKR5D/WX6hyt14nCGvI9NU0pF4R7mDoPkOQeDWuy5V0V
bN+vDsHV3/KNU0ZgZoz0eLIfBSMbdA8FOovl3KJoBgz2fbIT8gZ7UCNaLIrqqxCZ
6X7S+KZjw0wkvqwZFkDaWOfERZiu2+AFpYJU/ffU6S2oZOczirhMfJ58bsHVo3Tm
gQhdyAqyJL4PDpEHpiE3DfaBFv5pZoBsLdEg7DXj6KIxYa2zubH/wnHZXwoBFOcj
sUSPPp09Xsyrl6tj3xteQQ2nwFcvr6bOekBaf8Sv8Rkra02BVJrfBIuSaperXU9J
KNvUad0rx95/St9N4rvpgPEMOc12WnQEOvF4ns3phJan2eandJSRJz9WAVnGb0C9
eAa/OdU3Pus1kfpE9xeeGxju/Ygwz6UJf86mNKFNsri4mghaX+bH7i7KTDJVcu1F
SeRKFMNa24A47ra91yyjvLXVPgNnwEGr2q2Rmiw/0iPCh1+ridfwcTZeL6TVDWhF
rCRdAGpnI1O1vi99IYJjL8MA+apVBIBzASGv2AO3mhHWb6Q++5+2ZVKFp+XdGR8O
V/5xvFdmxXg3dQk9EJOAxL3wiO641hSZoUEG5U4rkgLIkr317ciue1oYZ+I/9T3V
+IXola3VCd1nFThthh+FPfNzbWK92Ha5RCn0OauhwaS3ivkqWhYlLKlscNX9FoIA
L1O5GV5h58uxN+2lZQXFmjAFfamZrEN+WMG3wjBj5XgQzaBhzczHdN0RQT4cTfpw
lJlTouM/U4UdRqklSPzMdXWFC9XDjpBp7qy2jyhyL/3pJcrbkebgQAc1+ov9SOJu
4lOhUQrYfH0yVZA+uwdkJGSIdUpRNrc8xfh15YELWXdOqQrkpk0pBkfvGjFWe1jw
cAp6rVRs966dEXjB3/ZzLQmyrEkHiV7E4m2yY8IQtTdDCAzA37wfTtNc8YyT/E16
x/NeA7qFdw0gI0maSM4F2oFUfjpvm+UojW3m9zkGfkVD3myNF87hgy1DzFYps8lp
OPtT+0WHEHyTkeZZXQmuYa0HSgMnvkQBDWWzuJ1BsP1WjLxPs1OC5fcd3Fhi/hLH
g5Vl9YFdmTj6fbelG3kBFxGYsT24+P45FwlJ/G2Hdw93Eo0VxJGGqhJ2NtT/ZIS+
hB7jdjLRngxH9xCSQmphxpU6dMqV1P6KIG77GjFBXjGxVyFYz2F/r4VtXlW2aJqQ
ayI9Y1Pb9UdCAIDj4koBzDrYVpJE8vwoKTp+dyZ/oMb1C/WMoQuQdWjHH8njDKJk
u6V8v3/R4E22UGPUVSCuK7H6AbL4fgmnd84q3/0RRDs/+Yr4ySkKnSJZ0aDYF5iU
cPW5a4c+BZlJ4aLQdL+JHONuXU0ACXB37fbgcoGU/s2vHyOB+PNZZpxZtVBJpwse
kRxXq7Vt82+BYB7kDiHP8fOS3aymEAc9xQIbXm+VyB25mwvG1zhEMO7M0OJv33GY
UklS6nfABNawuodkXRziOeCmMEFXFFZCh3iApmQHCOhrnp4FJCRZgAhgTKUbiudO
y8qJoABnLev8p172/9ImbyAYhccSsbNg12vmnkIgZcrMkt5gd4Sl/+Ad/szWTDt6
oO3yxX4j3Ru5lNg0TbqiXecWwAImUKxLEMcxyCxMlcKG/tEH0z7X3jIS+4/Gh6Ei
w809PDFybgHj/eQ1QCCIYoC0Wi+vWJTdx3u+ou29juF4oC8fUmCQTXUjHUezz50l
/gAm9dNS/1SIhHznEW6Q0+cww1ENxfCHsL9kTIfJXvXYiFcyEEFKd5gHVt0NtA7v
6Y/8I03jrp9XpI0SANsLBamqxm7KOIXTjXEq45Ycv3Ecp2fIKlb5zVIel6sBsrgE
KVrFCrYyLKDT1I7335Z9doBb4anXJe0o92uJ0Dnt/pHOBudJQENz6+LuyT2zUw9q
fyrN6nrR6DgJrxMIP2T+9A7UzgZ6PzQ8yDHi109sCoTI9dnI8hILPAHWIF5tLqXs
8WGt8A6elfrKjjT81vtJNcgBaB/R+CHA1cA9opnHWRj+bMroB8uS0R4lTyZmr7Dd
nfDBhqkmsXQZw1nBsujo6R/7Hx6E5y6ffw8Yixi3UXYrecpiyXvGvCfpIiM6SVba
T7yBoLuLHbjGl7V2AeL4rHtUH0GeQHO0rUxvqqkjbTEXGbuHGLm09eisNPFlVTkh
Hv3U7vXIHlBxQ/NNu1UeJ8z0BFYBgLaE0GWuMSeiN/aj98k/snq8PfHLelKyxw8W
0sKqXPYljbIvuzrAKU2+f8Y6T0nlhA3txeMjbIXzYCaO8L0T6pCV3aIAjYYwNDtb
O1NpC+XqQ84akhTfRqXngVs0EUEVid4iysBN8SF1bheKpqTuWnmLG96+ZCVYEO+L
+JqXtMbwzNWZ+bCfwBY1vbKgdcmShl6zamZd4Kux1q7bpT0dvlErOExieURiq6uT
wdOKfUNnDDoPTk/E7jmy99FFBLh7GMUYOudCWIbRcP8jQtjShTwQG365bij8zkG4
tA2RZQiZdyDfN7V0B51saD0O0LytxobL/M2L98IMNfEYIxsqTo+uodVxLphxYeXY
5FEPcJj/qUzKsu8nFpKHTzAHZHwjZAmIAVjLFu0s4+XJoqTcDsPlc0xoZL3s13m1
rMVk7Qs7g0L9XBy7TXJd0V9jHlCoET1Jepr5ayG5p8rLvdWh+UC4AcIlK/ftPmOY
vHOB4f6aAtlNZKDhcGLw9Ot20VY9visUIhn5w8FJb5A3Dsznhi3nBcoD6QkRQtDB
umnRGWkqZr49axODfgbxf7ixoQBNEk90/pqYpcXyOzjpsbzuAYJcvJQVqccBEEPJ
NgwVdRpGS5KOpfn2/YxdE6AsQz2v50BSqzRsFqWoyUo+oc+8am+Hv/OOvEEfBFjM
xkLqW9p9/QPP/Se6dcbXlay7TvuDi+vwQGEVjRRn0VP9fFlNXuwAj2Eol9kXsOUi
gyuTBA7xtVDk48viZOX281uh+X6TmVBfhhoVI/N2NcqHbMQ1l+DQvyIscEEfI/kr
Miz2kbMQrM0Vs0M6xVmx8KRsRQlBryH0KXokWWazCv3xgNvTtbHUXNJzuhiFxexI
CG3jbuibrPu3AVxHLTqiygqqqKtTRBCu4rkuq8gKSwJxxaLPIV1KJ+CjAdDVBaIm
TnQJ0WovmcIW0or/3Cwp3JPykEWqS3DagU8nwaaaymoZUYwNoYuqPFY5ncjY/pp/
AgnYvDO09/AosGx4FvBUbKENRedHDl6SBVcHlErJlHwlF+xwlU/KibxMlJ2Fo8b9
9xqpd5ni/l85raUJSFCe5zUXYPh+Wwgo+1ALPrm3P6xmlOMolph/k7ZLrQ52Cpq6
LcJCC0svy3kADdrRV4DsScw3bvAro5Ix6JPLErK1NnPPo6wfwKpWbsyaxaarNcJd
Y5LpcAMRP5svNJaim48e1hBfM3qEdnMHrl3XPIjklQ1rerPsTVY3u3QbdaMnv8aG
INSlNXijj4qKtfUuMqOPri3Z0T7pK6Gt60JJ+iTYu/ewC4Imo6cuOOMKz5+71uQx
hLW4Tt4U8Q1oKFNy0Qfl2kHOiKlVRlfGOCMzzhiLB3jW8cLzpNlCh4VGTirHWzoZ
1rIyeWWEWtT4ovDtClFxEleUY7A4Gty7/JG3FrjOfXvbVezj2vc0HXwgvAuDWJvX
g0ZXceSluYstQrjCjyRIr8tBOlZI0286vfeu17pPOgCpkgHhgnetVUGeCwvobVsC
Y1uMm1HVqNuCAL4o5NB8ad2OWTQdk5HPcsaJmn+f5O5OMV07w9SF0JWbz77G+ayX
qO31WccAIKpCyoB3URgJl0n6+i1/ktB/a1DQc/tCW4rBYfzEsptG6ypXxLxO9+gf
eThbm4UDOCs+OzUCLoMJx4PNVhpK2FcdAWa98IZH40H5bEHC4ukZCdgtML04In2R
fJlsBgIChR4TtfAR0+NkF8EhCoycSvqzsuqohxQpOHwrJNHtRvj6jXUVXsNUvuph
XJw/oI7I1GLDrZXb4LDaZxk+xEBcU+dCDWf8KKM+lDnp0lSc0Q3/v2ZjsQBVMnEu
F5CYCpzgi9pvqnhkABLBBl/tCvCE77MoLGO/2Hodw8wCENVxIgmAK4h5/7KGFfDK
a+isgEpNQT5e4hcbV9IoZXPq+RtFRFXhSiJwZRKoX1DoP+1IXIR1aybSWWvBu43b
G+YrE+ClSiYXJaFMdB0lDfz5obdMOCABrsxG9eTdjvi3WBUIhQllUPG0HFD61rvz
iQuhRJelIq9xNobyU4jPAMP9d/iInI1JdX7Nk7dAYnjnOUooTsm7LVYEE/OEUnEe
CuJhzTqF6eNsgPB5QVRaWl6L2nxgataKsZZ4uWD+nVJ01GU/uH7ek9ys4SFntBk1
zPuErOkerI/fKRyxQcR4AK2FdFLsM370ZtY9pRPswikCo0hfOiQ2aPQ8fKJAJfnZ
eqg/mVbAeac6/JA14U8Lp9UWNohiovMufzbQTS5p2LNk0Pu4GE/fNZNmM2MsgwKH
WnOmP5tKxTWFIxJcrME/XB+F4KOsAvnZJ+AjCEUmdvRcDCupcOcVd7s1IA9Ny6Hl
poq3U18LDYYzALXp4e2GfM47O9F5DJptKMaj8nEJVBDnVNgDJuUefeRiC/3C5ukW
izCpPvhGsfKacp0KCfvpMuOkfsIVIzy0P9BlxrSED+sZJYTYRAGg41gj4Fg62N+O
t2tZDdZ0oE/cbmMCq7tGI5ImrynoLA6ppZAjXCmebFK2O8Qvzkp+B8wcGq5wmzUr
5vWDJJ7NkuqsKyhuWvRuM2Z0WpUpDRV5J7oFQSwWZ3/lVwdTrpExxIPvyheq2xUo
kPLLWHsvF1m0t9GUik6jhPeOrCJe6Mtv5Ws1/wuFEAWQaiObqRvRcFlgFigHBlZA
H8pdt4K9tLt3Kqz+5B9s/W7MyvgjaZkq9cxrI9RbL0odglVRSm70/Wi/lQmaSRmF
crPCGCSG6YI25zyIufhGm99H/DeyFoPR6O+dF5yvqHXjkK37QJMOCf/5VEG9jZWV
XazxMS1o7r3VG5AKuXNLVyyZLKzhgbCfn43IIFPdKh50id2Gv97aE4T2ZFTE/Iax
CNTCyTu8b+AKx9QH0TmIUbHrCbyXmqqXa0QR/nqOxp6NuK9Awoy0Hf/qY4gM1SfC
92gm2Z5Sru+ALKYFUUy5fvQUoZMtEEa68IZYkmrnNYnrPSjIpZEP8GKJgQlHp8wO
qqVG+PVu3rGaTTakoFqnJTvMV+pPnsocooylMX/xa/Kx6rE8fK4Ps3hw0BmheI11
NmBvbNg9MCNH2uWaaOkrmY5e3YYCKx6xYY4Fixgz03Rk2hlGVtwWJU4If4QbS5xx
xra2gVAZg7QTyZ37ER9yb3zTmKa8kLngyFxxl+v1rqpush2k/Hh703QcpNMUPuzT
qAhhd+dk4nscKdGYcSS4pN9Xm9KJI089Zj2VYRqhfJ8XfRS35EHMu5IAhLPlc6g4
RjidwQ+WOSDDgJA+dF4VOMJMyUr8nppFkE6WJfcO479sNPbeq3dKcW/JEDi+HGKy
cmpdV+WpXhu76p293/qm20CH9rbty7CtB0mdYfogzZ62Jd8kmvkY4AyquzTxLpdz
nr4U1ot/Oro329VLgSwbrAgVfKPEQLfkp0IHieKjhSrhgUp98likg3KPlIt5jLEC
wo/vdDn2JAxqUvbr2kEYwYhdn9bv+TKtKC7AU4AcNJA5B3XGD5n793mSJAECIqdQ
jpCnvPMUhwrVHeUvvdKndVyjNIfulw+tQJNIuRTJ4a5OLHY8wfd2VU6V80ytFcld
lMybHLbE/tTKx39GTV8kssO5Iat/0k6UKOZu1OVzBWqPu44SECWP3xKGcvFqUKdk
+PRIRTBgwh2wEWbNBpvv9b62eA4NlEjGulKTupVOfKkvNd5lSu+mvH8veTuENVUU
kWbtDEdqYBZ/8YpV1KbIjh3LHWeWDPIR6yM7d0Uu/fsX9Xk+8tYGEWxkdnePuD0a
kJpH1nMz+1GWCzCnZXeuDxj9Xr5ofYcwwXx2woh9gTzOdACGMlbbT5HWcPHpbPzC
sE+4uamFlE2bRO2bgeoEleyDBRuaFFklRyYFwjUtdDeaIMsu4nygi0Qdji4X91vd
1PTwn80qV1rDWntah6RevbqHXA8oDO7OY/oQS3Pe6NZFaqFujdXG7yFwV5p7LPqY
2Od+J6EwjZMVrVDKIYDgl6XrSCrNLtTH+YdL9Usk/QjjBHbzEWK4ILTzaoEQwz4/
xMTxn5672qHpb7CJ6SS9ZgejryyO/I4vOipKO50XRLPJi/EmvQ0vX3Mh2117uDS2
6dnm506faTW2ocC+0Wg2huk9u28gEX4FoJWAkZE3hRWDP1shPat/wbmJpQb5nAFX
RGEHaYNCobxJ5/k2byiXp/11Bs3DEeu/ZQPuYbHWlphvAVZZ+/0rZx3z20iHrp4W
/d8eJWrWW3gRm9ez3ICkLUfwevl0pNNQzK3kQXlDELQrBgfBB8trYfLPta+riYmo
YxR3Hb0Fwp6Fz6e2REP7ocLqIMdRUy2JSKZS/DTTjq8FXGrn27VpIXv6chnmIItR
XpQdajX336FdK3ExrnyinO26JGChWUGxdePysYpRyAJp6XARJJz6vAqd/G6I8nf1
OO14o4gHD2TYq2gwgbB+zOolWdnFwRWdO+Ojdp1SeyEjVIRgcLOTcNAGCG6UieJp
H88aw1JlHUgDK8TUQ1Vgf3n5XGkK6hzHPcsHYJ8ymhIDctGb52widk64jRmuhjL4
ZfLo7iiRgHuubTFmxijr/q49zWU32gqyitd2mWB5ITsl/9oW2bPm0sPtBWBRVBQk
opPRtYiL4PClRw+mEYvq7PnLkEzauMtKrZre8NVXNS6kUM7GWrCGc2xE6gRHavaL
igh1FOgho/wsW2QTgL6UdQQ8VVzNHIO1GGiA8QVMIc0BpD3Z8lOYjkAL7WIs6nj7
l4duG0HxicXRAkQLmQY4i8tPEB+oj08o2WoFQlpxyLR63WmHn0ha5i3NIlPVVHnd
lfxKesdK5R/EWJZpdUg73lsSr9l8UZUZNw9DRQpkTs2ljooHbn3I4HD4wNt9ymp+
ZZZfswp7JVzIcHsNW61PTR16NA9Nniu/o64yJn7MrNLr8tWmPsFfFTWPOcWWemTi
iOHPFggcRCIcWWvsRe0T2henlfu/nj2qckMSZHfzFKSUKqolWWevj/Qlczkto7JE
TnHVp0gDc8BI9P7NgN4kU3ZUsxGhBPW6pKvWXmihnxBD8rH3iHWLhqXtgnHL14zN
Mn1kRCGID4ihpBpBePYMhQ7C4/avKeNXdkPxC4VbNPfjqFOJQOIPE+XYfZIJO7D9
+OCphq6Xzw3k3MAi76XvzKWPrlMgnNhqryglHHlzjoTulHoA8lcA5ACIJFg94VPH
XJ07LCT86HUA7qvLySOgA8NL8MhadkyXFGGKjb5z+O4EIH2Mt+sksj3t0/a+I35F
Iya+1lNSb4Yg07zkZnjAxHiXv/uSRbOCe/Z0CBXfwpy4vXXeMfK8Oty96Z70VleL
GxJz+0cRN3YhL1eGsRUyzZerMhzPF1aAMm4s/rORfpsF7OXXEMr/ISIVEZc4s7/u
xH3eI3pkqf0YZFvwLTBfQnbhqr++aiw1nYNxsltXFdvBWAwDXSrRN4tqJB2wtPdF
9oSilbKJ2HO8e20oHQEqrsDsWXFMnRHe/MAxz0FuudccD6OBWiuiZ+XiaTTXsBSz
XMIDTJSiYfQX8QAVwA6RDf1++5aoEXH8JR7GGiz2udUEGLx4UOCJnuZQMDoeNJlK
gCW25ha+A/rGFyL7g1SyftQ+BHlraM1rf+U43worMLZmmp0T02hi+K1T8/58Dm0z
WlRH/T9iGbSP424OO1cyITLmQw6VT2UXFQUkp244Nw4em2ffbQ8u3OM3MxagL6/A
3Keo+4j7DKSx9rPJZEIbTWWbazf5b4bRR6oe3jiLouJGhBzPoAjfC8ltWjcKdvY7
7xHj9HSwTWos5rIMEICEpRNA2QUBJH/vKztYy7Lr82B4f0rGuakOdagsarO9vKQI
tZwkACvF1khhrWjLPQ+PM5wvUTtxEFtWgyshBRXwgKUpouADcL5ZNmXKwTYgPTqJ
9j/V8/3uA83Nk42fv8SpemYl4RN8QIgFrMNQhtXOil/f9FTcav56Cg/zpuuBd1Eu
2o4I7ljKAZVdMFJgPRNX7PKb6k/3TOv5JfXO8TzIuXHsZxC1PObFmfM4UpV3z3/k
N6BwgGau6M2PyTkBsCOMATTy0fCi4QH6ysu22KZcy78RBybiBgPpsYU0Si9aJDFY
DMntAOHQuOR9RhYbXl6CXE7GP9iden8PX3afFAGfkO9VF380qHhfm9UZJ5nJ0iIK
ICL1wBDkqGzlAIAhPod3cN8YfgfFBZlzhEq+JmHV+jjjZVZzW3DT3YCpeygB9roK
Ns43GqA65AVoPduTgAz8sZl11yOIt23g+p/Hh4d6iXlkHomT03OzEr19pmQSJZY2
yTqNu+8BGlySugDy56L+FqUQ250MX4IfYWiqL18VovGZIzPBxNCIdftWHn4vojfQ
8/TvGEBXJqu8gTo2UCpPSG8Tk4+qlMKTWoBdTNYa4OMLrMPW75OIDGE9tlqUwN7N
iHYQ6m8WhibN5aWZVPuM4xgBBOAUlLqOtYHfPC+sxfH7qEp9eIRiECNrVp6cXEoC
SFBsFGSSWddT36+euH0AbUnDMwLAHr0B3PzAjVeBc/Qiqvw9dRTbtmS3f3+dx9uF
4dWkDEYVdvhDYTKxN2c4mEvBo1vEXvYTKPrUXMcG4j/1uq2xW+rMcPIDP6WQ8Lzw
N/YMVD0YrPs7holVC7QR9jL/JUhTj0WWhtNzfJPEUN40HGuh0FYRi+wvodba9BE6
aW5qsekMJt007mEg0zxeM3T+JaHqAmXk8mwj7B6aShTeCn4EDWGSNgJysJMjry8X
U/nEGHrTMZ9zs/eAdM0sNg3io/G9rcjXhFhvPpG2ir6arbHcBwujnzcRE9i7XJVq
DCeaDotPoPmOYGyElgeDlk0TDJUp7Q/1pW7PYz/cy8jY+ZA0kv9A4Iuu/Ub/AZ49
bYUe/ExInsPeEBduVSCsmrkWdRw9VXhvTBAH9ye0mqptU4+7cYIvPcUfMLUEVX3N
50arXiDdun73jkXsVf+KT1ZSiLru2kjbQK1kG4IYaBPqIFxDnWs0BTObSI0ZNOXp
JkIxa3KgI1f9jjb14rZy0ts+/H0jNEU62JAeE73uyAHhaUAt/P0r5YsTGrGfUhWw
R6nGXO/eIE1B1h0Uc71j3z1KumaD+0su9zCCqi52zietQX2/Na9825liyLqPwbeZ
76z8ElvwGjFmKiS4VqVneU9rJdfVQavb+cJGM/eCSy2mrGbYorRssumzVLSODjiY
Tx3u7/J6MZawvI160fiGIzZplSxzpanJGIjkuL2NqgdAONzAXZwC0UOXIEBVPCRT
cYWsXsMq85jfrSCKnugICRcsh7UGaSv6W1icuImuiTcxu0XnFYYulV10jYtyJ927
wWM/9t+Wl5ApTDlac9fvazvMXbA8PV4AZ6N7BzFsSIRplx5pmeVTOSqwCR+Wngiw
aLpl0izpYuEaYD45aTeJ7Cwf8ZnKxL87JQzDFPMNyGfZMk+o/8O3rpT8GXsI5iVb
NCmRY9/nCb7zduQ4wGhntsqw2dVgyQ7RIS+3jUzpRHcIYCaHZY7WQ4r46gZVqqPx
wO5t81h/l0CRz4gHawILQS7/vpALYWifUM5fVfocpsC4FkVWWE4i+VokV76Jd4uf
P28XV7cieo3bdMvR3kEbyl2m8mdgS0q7gZ3g3KnpafGizkidx91NWsAqLt1rb/SO
7e5NW4RvAffwG6B7Hkdfgw9XKMXRuBbVdVzjunEgADWVA4d1KUDkiiomHRxLLGnM
bcyVSf7eUe1W76h/6ROiBGf7JM5tkqBPhfmzDSHt5iyzhD9G2cetA87li+SUEBg4
8NqnAUBoUXfRxFhbzpZg7DVB3NZ4N+4eB77/6xgc2tKfY6GfQdRaVdVhi/KAwuxr
ofaUd95xr6NkBgPKO5bWF+/dNKnBl0b5CuAqhnfYg//6+pBGRiHMLTB4Ddk3hdQa
8ZFQo1deasFpsnUkEPkl4c/kqQaxL70TL7yXYPk0R7Hn3nkE9NpQhhjXf4/0GZ4s
hY6DPS9GSfNVdKcMA56Ci5TqD3KZjyF8ioA/Bx0CuIguJaTHpwl8SbXSQnM7pg8i
OavyDXtMDZ6vH6vNkir2U9oMgg4cKzORx3gfPLk0Nzn1vYh9Vg2v5npfEHKWKTSm
qRGW/A8+hGXXFHRjsTNKSO9111dF2GMJ2Vckg9NrVyrD7G9lNC/hZdPtOD4gz8OD
d9GmyQ2pBagKsB1iyIEnOK7NEfPcIudnHZpI0KZoFslW4eHHUuXJQn1GTpk6moZm
eYhPwAgErUSje3MEPGBGfbBEm9csi0ELGunKKkYgKPLourV4q60Y0NVmWIf/EWc3
1Fm5BzU/r8NEH2eehp6Gq7nt9wOg4qCpRRJsXzysBFyTlzt/2uOcUdkf6NMyWMyj
Ljn4BXHyX5ViQdfExBXGxD8cQ3Re5t46g8DHIVi3OAGLsan8NA6yjApZjuHGflPM
y678+DVXrC4QpTu+PjJoDO8a0sDvkEVpS5d5EVpAHqcaUyzlGcZTpD5pVxIsSFXn
JR514kOOyJubSJ2q1YqdLd+6FBVvt+rPZofMfDc7rXm8Jh2DEYfxE6veRr/CEyTc
Bwd3+sUIUn6TrlB7WENapZluRliviXDWQg769u2++b9UbnTQeBHPgN+WjXjNiiCa
3XG3bc2p98nIwyjgUTOtSUQmFJYG/vaXuVn8RYdAqXE2O+nMDuCm0fLE4Aoj1c3t
/cgq92Nzcnz/6ic6AhdnVsAAaW6Oa3f+l1du6ZIvfp0pTW80NOKap3RhX+VGyhJy
g9MQ27E3ZP7HY34VT3FI2qWifVl9ciaAXiYdRGhU7ktozMhQi3R0VsvCVLF6aihA
P+2cMxgvqrI3koi+eBtIRLdYlqrb9xjXp/By0Cg+lPipu8fRUd8YnXL1b1M9wCRP
cIPxXOpJxcdfn++XuKpRAd7nHCe8gh30lRPnDm63i+uuKTewx6pvuBHFybbGzxIv
SvJHVnhfqF2mtUV2DUl7XolQmr3tsaj1QaKvT3X6H9tvIAxsFtqDn3V2ZFwJ68NI
f/H0TaNitFoYSDBs17J62qxHFi9bhjyUq/Ve4XT2vxcyeUp9DBn6kW+em0rWY4Fe
KuJjZvqaIWTvYQw4+SsGej04IZfPQWVGq9ynznypZJcErc3d2D+EgZJPNHG7qzgJ
5j4Az4tFand8SRLdGS/pNCj2CUOXrE5NIFhEBXN9UHu6l4HUv+M5PqxbEfqrU9dL
eQtWhsMTo32dfGJGMAD52DCZ56ea8bEgW/pSlODnd67mGzYbp3IpsPRZc2CvMFT+
D4nzT67tQit4B8CWIBZkynBVDh3lS060CmkC8rsph/O8BlSU4wxIXxzRxAf/OP/9
RwItiSJRSOtF0Cd3GUkBIAd+w22oKgc0VnXffXHMUCYqsqxX9mLsZ6QVuRDPK52h
FQdOW2eFEGwrqXWEHIE/0NiVp7hHaksbzDeRIu7bZr8BQxaQoj7RheQlOdAUlWGS
JGKUiDaZtpWM+6Je01Q4K+OZh3e7m8jmVrpnz59ao77Se2Id1Lj6igL13FRA7Aoo
fwe4a7J/0s8H5FL60uxknPiWfqgxpgoLRu3dTGn53ldA5Iz9RUQQIsRQ+YiWIsTV
PAE0kfsQBmQ37kIw4Xg6Jl0/EZq3Whi7UZ1OBhcIc/X411i2IwTUF/ILTJsXBqtH
94H+dXwGdYVKqIKAOGYuA9LbDjEEimtaBCv++9lExc+l9+oo5x0sAQC30pbJALCd
oq7w1F3Tt3/8KgzTBB7VGr77Zd5n1lPXp9N+NwoyAl1otIt46HKFWLLo6iAxFo6V
4bxskxAFEFngxt6Vvr85UP0l0q6lbt3QWviBczkb93eaJ2mYoYncLtbaCHYQ8Qit
5IVli15D8KO84BippVpQAw3SPQLi1qS7gDlaCWVFuW+R1eyjIBZPpnYVXJ/HAQ0L
pHfpXXNSjBIAdVCcTKPTGIZp0QPT/L3Ql0BfkdUTHRqGITDEE8Q9Dhdt6+cCeUrW
fY5wEFGnVGSOgJ2+IHnkm64DNMIGgz2b5bXpYN/Bdhseqmj3o5Q1pjanw66b8Pad
Ome4H2krQKSGIlL1pXIU3QOw5N4tuliFi7QVhEqzf36XODit98VK+JYPyDlV/eTo
3r6UGck/Xn7DgTGrtOJY6X1590x+6tJx4yz+t7X92qMMJx+xvrKDEenvj+trSIDM
4x6wrlT+c+Lc0VwG9IACGN5XUV3gCIaCbexXLQRHdwOE6A7g0yzV98vOJrPVEA2m
UZTAtTLYrXAlMqUikHRMzCf/nkR1mlGS6ZuTKCR6cjfHF0FIr0pULbkhODCpzuWx
6rE/Od2urw1qtYijYimM39OTMWUYwJ9YX1V/sfmp0ugJBmFHIpmhiXi7YoM9kVEE
cl56+sts88KIPebSkIUW4g8FiXHmuBMcrY0b83P8nSpvYdO6cD1bdSSgPjSFwAqL
i+lBYFcO0ia5G5VpW67g4YtNDfrwYW3IoF7lqRrKA5VnIZV2CODnqUQcxc9sFkfv
G57oqs5ycfZ0FtEbuSUzazduwt3bxK76Rx20WFhFgM7fvLER7fbb6a29xLDE/nlu
8TLRImVDNmkMgQviFGbqLOe6GfJo43RScSoNRDH/8dXA7bbRPPzQwJ4lXQD9iNoS
OWsNhGuIJMrR0/EEMGZ4XDtnvCwZyjnw3/2lLxI6iTKk22izooe5XMfWqsbc7Msf
`pragma protect end_protected
