// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L3Sjl97ZZQaOxBGF0xX99aWPJKssB5qnYjj3bJhed8j/N96olIEaQW0z+qhK8NT6
RfsFKfdE+1lfD0Mb5Epk6RlWGxwlh4Vaa922JwnGQ2LbNzpGJdboa4pEc5fxQY6R
eaVlx/Fu5kERXYkfyTutBQTeJfnFcBnYWXv4BCSs/CI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12000)
eL2uZEAxDnJa8zgGS9fRn/xdAyFscLUIJRR6msiiVDuO2dvg9s38xbGGyapbss8A
WcHbk1S6g00/YmwFCEIpW2A0uN052Jl5gy0L7TLOcbiueva40GiPpEfACvZ4Piuj
9+jITZmwGE+kRf/iB0SC+hoXmbG3gmWYcD2mBZjnKLMhPW5RuYDNakSNXReYF/+N
tLIkGo4f5YTMNeePDD9eSG5Pf3LB6cfWwqOWVqQp/dUj0YBcpx9ra0/969j5kuGM
ze53GfDsjh8AfmMEpgA4NjphYPCHvJhmXdy7zeHjJL+V9eOg2hK9z5ik/sETqycX
Z4aXAxy6H/yeB2PO5stwxZhlEraC+6ibJ2sjM4LLhJ46jxOeNmi4sjBk55rW92pp
vSGXS59NmCgTvSlqVJAG+h3vawTHYbJ5klYVTKZFOKzvfqdkoCwrI0kb6YJXCx7e
Xjz0gi72moLaHfUHsTJ2Xhx7ixmi11GH8fRT/QjL3bpc21CaO4r0ryi6mW5IEe+U
YypdhXQ1tHXq+n9GOveYKx20uWdHap7XlYDlK40juowsl5LJx6erQAtrcO3tmqfy
+5ivMQfwHVzKlN/aTOX+4uDkO29UbCLq31FfhqAKmrP2KtCW9gb2Ztcjsom9MpUB
Oj4yyaf/iF8AVXpbIRfbZMXCLHlyDjuGPN5mxDOcFOhuAw8BNqs00OopBmvS+dgD
VAsPviaO+hbDGpbdk0PPIIg94adpNKcSvFPsQat6MDutXUbYTGMeAuAcLomo25nw
3HeY/SLt/5lvDSM1sBxlkRGF2lqvh0500QTrzVsmW1EiVYu+ciH4CchGG7qDl74O
3EuomEr11ZR9mDuW5MsmOCqGZb20uuoEJNnlaJJeEjbofqmYyQVU29ku8KDGc3HS
UdZtPAIUgtv7t2hRz6VHiOJwyj5PL0knoTWO2cdUDNtVF6hkNAupV7uNe1PTwntP
i8knnLrSwPc4Gowrv9uuPRinht0Kh+koheqmtW/bjjnbgYjRthmIru1q2rijjZiv
YaUSD9wOA0PdkPqDSQKHYfsCYSrsF567ZIy1vlXuFCq8vGVEhTIcRSUfLNQxhbfE
B5ohNTtPACLIPoNmlL+QAEoMTXY1woFDEjjJlI7lmTVDrSGX5sIdc+JiFOvHjDAT
6mEIYCAmNg0ioKSmyaFO+ZlLlYXBPz5ZdT7ZWxTp8KJQ8pKxfCkXubRkt6Qfq21c
49pIZ1tx309d+4n39qBjcEK2ph2o6WQiuXUJwiUJmstJJmenPfRr6fGBMTFpG/Nw
mUOAQshWZUdW5Lga2EaZmL9XGWn+oE62mLoF185iJSoyi2E3IyL6P01+FbjURHPf
kGWh3u/+P/q7GatoUi8ULere/o53QE/9lV2lwQ4Dc81nU201lu7Tj+SiBNkX7uM0
oTwM8rgqNJn6eK61yInHNH2bk8yM9s8nxJ/YpmxAVrrAECJGO7+8GVM1KFOtpejw
sz/ovDgLwJq+u5vZZKrkeKtMvbAGSUL1Tf4jpKI+dI7C1kcdfxg2jfbcm0AbRgiR
pOlnVu8PxyXKC+yTYR/dhAMHeGT3PrjaswT2Q/cARxYRO0gjz1jmh2ieQ0lTR5cg
xd7bmdcV0IdJYJ+zkbGQBWfcEbl9QSsIbyzA7s3qiursxs2IDNyalpGRHiKS5PJc
Tp5CoeKZZtNZj0RY7Fz+I2hdoz7bdfRm6vqKm9klMHPVYDUGCpc74JFY8jjzPehn
+23gtI8k2+NaPzIGkJ1PblI0BIwrW3POAc3py3Ffn9zVayvtjko+berETGLrooW3
V0NspbEL6LfdTNQ6YDGk5Vv3xYBgK59iQsQptEp3JqLI8HUCJZsasESSWhxEl6cQ
AuvB0eRKsTpXGLtnew5lwsjSKCaUCYuSK1u8W93pJ50McZO1bFBbeRruvLdp/6Cy
inyUOYMf6PLe9eC5Xu46DwdA+SPJRlYvTqP36lF17oyghpbi88H4R5XfIFSmU4Jk
wJqemnXcE/RrofRkbW+p0FV6VSbvnuZmx6PB2p7nY56nDG4N9WU9H9wjA5SXTDHH
cxQ62xlKca9aq5IOa5IqsQkyFa7fmk/LfKQiIRdb4Z7LqA9SkYjAy9fvjsLeDJ3Y
ysaM10RdfbmetpNcCzwRG6hd6CxhBkNsmaps9N86wcPO8jfz2V7WIDxLhhySi5Eo
qf7tZ+HxRGnkOtLkV6xNLUyknqm2UaSHMNqMNXqUP63FtOeY94VwhGpS6+OOo1Tv
D2/MjLVI6zifU7oER3u98mGyyeKW9s8sq1PLULBEN6prlVJ9skiaaxJt/qZ4KXWT
iuVwtTw0XvUnpWCdV25XO2bCxclQlM3ymWL4o9HEjZt/vEg/uof4YeNQEzcNNi/o
R62vKZV+B5wosOg0Nx0SOJQ2TFZIARUw1wUQyMc3ZJqfSA6XQ5eRql31aWKlupjD
LKv8X3pueJHXWpbxPAWU2oVYXBlSyiz7km0hqP2ejEh8NOZok0M2M7CsIC7LgRxH
PY3gnfEbEvtH0G5hFs8VOlitnpmYvx1VnUfxsmzm5jMnFKtENJi/E3WLUJCPoOpK
Kl96OAM/jpaBUGfNlw1uFZsStBDNs4polGrFTgIkCCUsPclY4DPY1CkSqInRqStQ
4boUqM/snUDU1BCWRP29JvaEQvulY8ENLIeNJWJUTeiAhKyn/cGIx0NNQJsSMkUq
XXpZ6HAtUzYd1aw2337GInSIIBJgY5PlkeKeo5vtRhPQA31IzBVZOIByXcG+JcWH
dzkRs3ZwOUc8s7kM8E3HIUFyp5OBIzoDTfUnepon7cy6rpDhNrp8QqUdwqzFNoAN
6wGzsa8Avthq3nlNH8YVYAfikiN/ll2zTQDWtTxy8gTVqa/TNOn5OEk+YAaNGKcJ
RJUD92GPzR48OFbppIgeUlqg6gnqI28n8GeXRl9Fd1nOSfZa75xp6mKMETQgAFLW
LUiGTlW+/OqlrWy1brdQSG5Jv3jv7omkfjoZdVHBN8KPwC3c1RpYyQCSZIAIKaLF
LcaoMPZDJpO808zw3ihRB4blkGgbdGC7Tz+BjwhsNSbbcdx4jHmYBVz/I5MQ5NE0
PWzA2pmsBuC62unAj25Th3QP60PivWHIOKTzkI8hbUbURfhrxMDat6iqs8ok7kaf
onXTvWm3asCvTLEShU58QYi3QjvldOaGKeorYIfCcXAbFqpi+9U5fKjn7MviOI5p
YrRtDNPWysgLiLhaeUBXge/PIr7jCiZQ5zIvldB8UI1NlCsww3kLZY9d/IMSyczm
Z+ykSiu055NGd9DhdA6ZVnIZ1FR3QJHnm0+0LVgnvY51u+xDNPbY+oDaS5lfMAqj
/Ox2w7TIHeyj3ekfP69dRRzsixUtcxHTA/cfU4Aw4yOeuJj3H3QnTGSle0pbpaOi
Kl7qwNBso/krL08cd0Op3jjvM7TwAXB28ESIg6jSQHg6I6+DyDEr9oyy12e8e9BG
6LeqCYy3lHQYW6s3pZgwyIYOjKlSVnjwA2lgz9bS03DdSRW3UDK6EyHKm4aR3T2d
3LVSVtPwlzYS9Tf0SeeM3/vrB+FXzSdSGiyO4gd6Dua9SFnSjMV7ZFz/smF/fiEG
LxSgdS08MaOWZbTaGpM+L2WJID/vTqm2X5VfDDkLK3xvwaekRaCSFaCJHM9dq24c
XTl4FMZzb8gV0yjRCVl+GyEwHTH3Qvy7WB8CRfz/o6Thi0fewcpuBJhDHSrrMO8O
HQl5NOCoHtqnlsN+shf4I7aHsKimaDsUAghXGFSTvp4vOelQ4zwXoSR5EizHNuVQ
XV/PG3234n7b/vy7FhWv8dYVsE/9zp8GhoNLbDotol+8p6k9aykT9LqvrsQnGpCj
v68To0M/HCoLwC0VSdGYVK2kSdvv47PT8Mge6ZZOZG3L6KvnaiDNQ0B9ZgY48ftq
vV7HvY3V0K24cC2whXqyFij/kJv/RudjL2rnHQea8lmOsqNaXhLUEvxy+vlspOLy
/TVP8WDOzF3J8ZeO+aWSQgzCuOPjOxzK7FC3agcrpS5JpfKTIuzw5hEh8Saz4J25
3Jf4zZ4vRXonbIKJBc2g42gVOqSEj4yvwsDjC0PUZAUKjrISRO4nxIQknCCJx8sa
PbE549THgwX4kL5vh0Oz6n2Q/XbNYF7mZrJq0zBpuO6gKpf36Ao52RHKw+TVLHcD
skQOyt7QskC7srRdKo8ufnKXj4IymR/9QdVqxOD9dO2Rr8BTx7OsxBgZEuH+GxNj
aULEm3AulHPn8bjbL2svjIiwnnkMMeKxIyhh0O0dU+zHPTkN11RMEv8lKWXqbLEj
nXOqLeymFQWJrObYd9cL+UM+Y4YTVYlBmdPsHSlyzycyCcfUpdIpVmheTYHj7U2e
8uWlWJSvEYDJOlphhxH/mjy7ZJdCV4Fg5buYorl2vqasTcC0fnludUOzotj7IF3B
EJ3HPr4uvIzdyBKXvuunhsMFBK/qAtATF3C+Zqv2wrC+LXne5GxJ/qwrjnJhjvpG
qmYENDWGznhwW1zlw6QWDy6RE+mLyNHDSWUj0OeoxTgZSA73/gQDwbSaSazYNbMR
2/YsiqXAzlqMUGnwWLjhll8aQPfLwMjQhewVeIypHpQV9zljvrw1mQXKpHbxtohT
okNfLBk1nB07zGmBeoKAMBtYWV5lnprT/sDDFFN1WPaRWP6Asiyd4qD10nqxAvfD
nra+p3vrsusl2WyeOIzlQLt80w60AzlcrANdY3MlD8wCgePizali7w2AfH/lX97o
zIcRbr4JUUukSKuDAcwCe1mWi18b/lmP5agCIvH8WvG0tvsSDmEnyfq2j+etTV8u
zAL0hS9+H6vWND3hf0gOkQLhs4Uf/TZuyLoDnOK/Y1UEzPC8+eVQiZLheVEHhz1/
GA/HQgUqXjEEQdfM6ZfN9+uQWt8FSkia5kzk5DGAoFW5iFqKDW5eoEuoxxTOEvI5
ZTn227AQsbSEW+4xrolO+pWJDb4SoQwh6Gtv9twTPb6TpUeKtNGCSrK5ob6QYpNv
j767caENbiKMExaWjT1jHicsvNSVxWCBcXirlKsYpdlxnNoEKlXj7Yi/ff/PbEsp
G3YMAV0Obv71IniaFaioy35gzpn+5qOPy4ea01JuB4KqSLfYVOd+DbP01DssGKoe
hs1lT6N4TG+dC7HXxtBYCtjOer9yrn2o8niZlPUarvU2tMLS89Lw1OUCBSI+iEde
Y6tiJ94Sse+ygL3UAhFtXh9rFCuZDExXzykarf9wog7MwQEeGGJqLlLlGF58hZQH
FGvKpxIFPtOheHo47SMO633CLPsv2WOod6GqtjavdvkGAQK9HaRfNhQQXFvqzSKl
cRtCDFKmiOiJ3HoQMANQ4zO33DhT0OHfH8loWIwB7YP/0xoWahTTKjmLYcTiN2EI
ijwRWZUYIZI2nlQ5rxDvIsiosit6GqU8V3XIV4Si/MO5yMhBRlw87PTeeAhi20up
lTeKaCML8rlbT6IFPrYxoUiTRMyG3oWOzYUwmKEnht0t4+rPMlqaG6/FGhCJRNrH
n5CymhhaYNmlaj8eDZdtVdoUrK3lT6WKZZn4qs9IlOc/6PuUDSXT689ST2t0yw7A
1Lumx2Bx5ZqmSCZbRIZ3Ld4xzl+AvnrUpCo+fxZR5klxJxH8cgK4xks6SiqTeXbK
DTkDOk/1q5JzCxVr0VKcMxJSdRd5TlNS4deZt5nC7PyqnLZgORuM/Cw9zDAHDwgN
JjZZMwrq7zKKJWqpTGwcGmaD/rGeRnh7i9rNuaRzndV/XeMCO4FphdP4tgzAc7AA
Zl8ZPqycosZ6bA3YyfG1KQtJxekATdox0rwQf3QqHfoOWLjFhAc0nS24DDguwZXw
JGMLP524zGFbHV2qIH6+iOwNTHrfSoiSiJrB3qaFbpT4UxCGbSErnTWysRBoepci
Izzb88FVjePkuJMClnNCCSfljAYpvJeAwDYSFIluXIy1LJF3mYX2U6XOujUhEOvs
FoVUt9xoN+GF9fZES9RaqRrRADNblf77tbJiiSukvULwHFDG6p/Yz/fBIxbNrFoU
m1TkdyjXWLKy6kr9Rbk+ux0qs7VUCAh3Kw5tppasEyviv8KigLBgfaZ329q3kSVg
vXyF9broZS6zPGc63Uw0jzWH8X9jhFvuzgkIb60ragaqCMv1ERmEFMA9ncG/zS7K
oNF0AD8DnnaASNNeaHf1yx08oCbepbj5thtUpfDm+mDoTJVPiO/9BnwaH0Qku6l2
B4Nb8P9k7y5G5cOsz4JX6QbvGS7myn4tT9i4QdA0gpObogCOl8xZu+MCu6IhaHkM
fl0ekLi2V71t94rfDVmjglRluO03nkWm1et/u6REkOjOWuHB8YmN6KS5O2W78fXJ
JE46YqsixwEgZrCfS/I1D2zXWNGW4DNdkZ0ebjkEXX7R4IzUszqQ0YiAPFCgvfqE
IzuxHz+H/lAStBax951WxY8E0EmHu+xJrYGOFDu9WBSUPPkDsuPkAdymWgltzHEG
7fMuwvf9Le5kcq3alwigcVyGm4vCMshFKdDtSWnxFiNtL8VpNmaBsBXDA836DoO0
Mb3tF0rMAT8VOBtNaLGQrO+UIpssXtCV11J5R0KRqMzILn9pGopv4yU+ovTwbXNN
5A2rnyoNSE+xGwG4a4BqWAejFjwLhb//PMLKqzN5TTZsa0TcR5eJogLyqKT9hyRS
faH/Mjt2byz3BwZlo4GDXErqmL3+myp+VacYZamIWoBI7+kF6EmurIl9SndDzpPN
+aGX99AO2QnWZZuj/4piZT/eGfXx9mrZsEpy9Xeq+9afnbBqjsTeqERXhSEaETCt
vTvrkKvMyzurz1sShHDWVzQzXkNonSHi1ewWLemwHRdqCJYNAY8IUQcc/4OiRxrv
z/ixKIM5wLUSohTB4R5H8t3yexD0q58uGHtXOMuHK/6MpqxQNUbiazHRQaWHrTLh
6eMNsfIbAjHehor1kGle+ZtJswkDNZjFXFpt8G3nIOQXzEpbzoR/GicZ1ZG1dqRS
IDbxfR5HCgqIKz5skvXL35dNYXOWKDOI8z+Ch225uhucny8EELc+wRj9WHIqeCCC
aeRNQR/PLdBwtDFy+hKts+OWTgSOwe147DnPgHVFQPjcRPyioYBkJDIYYeLNjTju
wc0IYDaxov/XZX5BpTEQ7oE9bIybOXYSAC2F66MnII79HV3H5rnNwyPRsZAvMZIH
GxiOnKKoSWzminClPCOsezRB3RXvZZoU1OOcqxYNugmeQzH9rdtMrAr9PCk5SE0u
BDwQxbI0RRaFzJzuDBgp74JPiTY42WN06HpYbtjlgz80X/VIBakxplMhLd+PaWSR
HFBJyD5bTzZO/w/P+nDbgzPxmItTeu4sdytRkPv4+NlZTrA8Sj8wXiE1i1NH9IHF
miZFWJiDW6C6xFrjRt/wbWbiBoS4Kj+g6ySLZaoGszYfHidI8ZnAdHeA6VwcrBwC
vIzcABgVcnxsuWNJ+x+Yp390Yboq8C53niqW0HqrWdFAEvmSEjvq7PCkpojb24eJ
EToWOCRvdN9mm2gmENPomu22tKU+a49wPZd5Yg6DXQsY1eHspaewFsRJNMdxwag8
Rd+MYI9aMI1qYmLemg5cNHAEeSmXnzei8PdKPfK2883dRBdIvsqsKlCb+ax61+ow
LWn0qAg5qjgPWFdjnF32m1V6aOlUT9BxFYRFnPBreEKN0Cyh0tty5x2gMfoWvkAN
7aDnMuYIWlhX5hlHruwO0AyhWQjq2njGNMO8dqDaEoW3d5reBFk2EGyI+SAcM6Nu
m2US0tNsSiWalYsJD7cNxs/XOHEwpjqq2tP/pSoqdkXsB+G4z5XGZL+7/2v04y06
WbwLlscarMeLPuQc40hGpO40HqCfXNhIXPrpbgqAmwR3WUyrB1+N5tXryWDLwgn+
cBiitv0M6/2Ezbnbr3+NIPKaHGmiPqPC1AvXCdxVtvk0TkUqVvToKs75c0ExdaqK
+HQE+XB9FaRdn47ZLHVP9BP1PEnEApZc1Ev39kIjM374nKJCAGTENFlUwlBsmT9B
tK8doAxSOwOHkZtumUu3mDiM+/YIv3zWhimiBhvUXnBzlPFzw7R/JgoKXVwGymKC
3myKqAVYqTJtJ7ZSh+MO30jKc3QK8V6ltjlraZb9R6A/mje4K78FU7b92kNdrmdq
2sz5J77cnvpZTANVmVBmj8Nu4y44m0RU21F9SH1AAY425NR7qtjcg5LL5XGDUyxW
J2xsYP/kWuf2awyyyzmviu5n1W7vrP/u7Oseez+du8/UNhffO64I/y2rf13r3u/v
7FPozRcD6Mclq57buqaOnT8oOGvIFm+yfIbKgcLG0/5j9Vi/TL5zNBVIgh3xVfTS
jRxjxijzyyVxVVT56mq5Fbj9L/cVNvhF6LU3vF5PnSxL4Fjd+kX4u9yLd3zlSZVk
yAoaAfhIbYsRQY3oklfzfETBtKnVf+6clnI7BQrwBwwYxrNt4oy1CeHsTHDUpOkc
hocYr2jTP7tEyUFSze7VHpce7b7NdyWuOGNd8Gc82KdIlKQSBCfLZrlucd5epzEi
rhJpIrymBNt3uNp33obj7IUzXq0LSwrwZJhKv9ddW+SX5YHKRTL7r/Uvc+06+dEP
h0hViZIU/ulnoTY2jI0d/k8IIXMrZSx8YVY2LGvE83y6g/b25nmKmgpukvrRJHfH
8Z49Q2a1LazRIyI5p9GFh2W7O0y37nCto77VZ4aTl6wVXwprS9LmTVIeP5Wdb6f+
DLM9ld1Qsi0vSdXYbk7zgrCEiZ9BaHykKGKLJxfDl6vKOuTFgfaIxsrRxH6BphGt
xWFGgXd3sUh2S/Kw5BrYaE0YZ+5rW5mO4uXWKyAlrpgkRPSxRApb+UEpSL7EuVux
+6B3dobaNyyREYxDDtUFHt16k6RXpEgDzNaN5+Zyl4Umzz7ZA45um5fdnWC4NfK/
EMCEpEGhWKzJp3k47f7QQigmYsBlP823xSU93SJG5Nx+6gqEOi2qVq3RWNXx6YMh
9jFc6h5rtjzPfz0pEioMtaoTweaiylBcatrENr1/OTceon5Win6qq7x2b0j/bhO+
WutlCkulnurF50qS78u0le63dpDDwFMwBQGKGxQaHKdF75Le4WmiYpLdCieSlOOr
8CJIfaK9hb4doInTbj+K07ul0ZR/hUfdcFBAMKBiToYidk+Vp15ZqtltfrZGxudj
6zzhOMJ8WTx3LLw5bAVz5xNUnwJfUsNZo/U1aQzOgrGLB7ivqRXohHkvGXaL/sac
U0RZ8Wu6wklSL+MciFMN2VuJahSUMIR7V8zUn63e0nkFFKOHuZwOFMlzmKixD/yG
P5iiDx3QxISdXvVFvMPBQ/f6TArUc10A4Aq5QeLK8xzqBF5nydTjx+pcOOl+4RWN
x6nGWfUoVWN3ba1gNjCkbV3E3jHfcVbXzGHP1XLsL4zMlV0M0vwj3UssjWbcZaT6
1U8JrrHqbAmZeZY8LAbkerONN6e5+9r9846+Ahf7x+Ek63Qw+SauXIkTND5Ng1/X
81odz12IIRy2AwtzQ08PY8LPSgxaXuv+6QbrDi2VOhz4CxTvJhBBt/JMhBLl1LhF
vvy3yvUMMHL5R3FRMLe1t/JNSAQCHnIEJeGov/BxEJUsMrLDpA1GRDte95SBGywk
I9Q2LoOc2416+VUytQgMGTDNShQmLoZt6DSsCkA96xWqfx/YQJq+26mdVPHp92Po
+hATQ62yrV+0Yyfk9zuBdcpr79MZB8nL4uP39RGm5O3RRmfuaCieC4X/DshHG6op
EgTLpkw5xK6aN276hKDsZCP+Rq1wLJnopqsARbcpnrjqZTH63aAeJM7pZbNp7gZM
X+TPeHfoPMOtpCmVDM7hSHYfB3N81On1W6Od4A5iNbMp/zvAtZc7UPFd4wNKIWs2
Bv1Xe+fFG/XaIK5htuNtz9PSbxLYJ0bmrVA8EAOITNHUxVVSPD/WT9gMQG6UGufW
SFR7h8nia541nA5tC/6VptfuC53Q5Pzjt2Gs5o/Yqu3qvjQjmtL35sqI8HbwyM+1
xlp1h72j6vakZf3j/9knlRFvPgM/X3TzqozsIyPOL3bTAbZAiZrNcyhPWho97LXe
r+Skd9co/L/uyVzQtYcLH8MC0bMcRNwq+wu19AmhrVoTECFxREXfSduIELtoZMX/
/cDgIyCjgMLjV+p02dINGzyR+e50nqS3yvnFsMNyZ9rN9g2+SWwKo3R3bjKRuL1Y
5W4OuXk6fZNjtSF+LwssQz2r9sK/KzrCjiE6u+HTkykjPh8w/Da5PDt7wjFG0xJl
ta2fw0Fl6waeQj5cyyiuPh+rELy2wGix8KcK0VCQEgOgS5rft5Axr1bFTZS75MwG
nfjHgand9Wc9bo/D0fy9bhcUPa+k+8L5tgqveIS5y78ml/iqj03KVvflwZW80P6V
25VNCiHfiHCoOGe4Jj1ne4N12vqygDiDCygn98+D7o6pWPO43w61zMflYSC8KzLU
YhX1ZDjIuHpA7G00DYEMEjSjLNH4llL1BNk1N4dHRYLyycvjZLi0eoe0D4zpOZhi
e++BLccId2op+ltCUferIOfG11SgFYsjQONHOKin2dk3SrIGyhLrc/6DfGJM8sfz
eBfNBIkEnspqbAWqDqllBLjf9icOZmpc6QMQ0NQWwscd10OnVuZAwpNB8IK6Fkm5
IWwouEQQHJc1UtXXeSxb7OlPaC0UUOCnjOHyYlLVJPDZkpvnG/URQS2pilu8vJJO
JmZJ/5GPCdlQGuEMN3NZj4qmKU5CCbh/A5EB8Z5P9aDygVT4T/a6UighgfDxRsz9
xJpXNEUi6GmJkabaAIswb34pm7e+Mmgi/dfBu+EUSUQyJauI9BeYbPCJYIMDd/fZ
/jmR4Nv6kcNKHiFcvYJvIBA9COt0YjObUO6nRaFNqA+l65N9ACmzAtxjbi4Noix0
EwOyyVUr4c/XWw+t1vnsMljbyTidUDnL5EFNMJtnreZyjQ3Wa2RkE5oOuYPa8bww
wnnQ5R9W2xq9PkmSGiOkdZ90rff2aVe5iMueP73yulROuXh2VcBH7QPV3UkYhfWf
aDIGqsl4zE85aEx/AjQbt/39sVjjLPxr5iCUHCvqjq1VbR38jKFP3RjBbb8tX9xE
/PNomA0i4llBzAAZlREGKs72ctlqm64jOo9a7cMJQraxzPLSEqGasTZVNNMOEvPF
KEM+P8vp4+mtas9E/5DJQOoo8cGzhkW1G+lf893YQJRaufJslFl/0pUqwNssv/BU
nnf1MvADdlwftJhZt7Y6ENgJbpMQ+7v5vuAT4XgjzBNtl7J0DIYrvtGGrlOnvd4M
jc/Dfw6OoFYvOGPLqgKpoCUxAbXjuwH+P8I6P48TDV3LMlgggkF0NtqC5O8ceDgu
JF2GTGxU5XK3HS8dAoh5NGgupaB2vSEGFb0dYpCxNX41INCjwFXMpds+4+W4cNbZ
7e/2FWBebgWlzWd4Bnj+C3G/Nrr001xNEyhNp5jxdeDT/3ZATAFj5Rlkwsof41H3
M2dwcPHnpoRKb1wt3FhKGF6yX1JkVdEyHgL1TazHLL8MbYZE53LhuzFcEO9ygjTA
daK1GOhBptG+iY+ksLL8Rum8kBJ5K0XSqfKerXhF7v9fpj+rsQDwEH60uOwvmtDk
74CpxMqJRZv2yy3EVjhKzu54CjbAEgb3naRn0O1sIB0myKaFxxL2dTSrDWXqeMNl
UyB3jVhS4iI2sc9v2aCU7NsaK/VbJxUbyGSqX5NqYfGkV4szDMiWElKXSLOXnTua
6FhxRWhOLDoISpR7lMTtz0tMZ7cmHnaXfnibY7ByBTpEDbNkDNLHO+z/rS7xpgzM
7DSzE7p2Xe9/4cuyITb9giCrYhpRrkBmOm8CbJMvvYDepcEOi6M8sCG0OONs8/nG
96p7C+7auQH/vyKSSkXEdkh4NWeStcv/aFa5DXge4+0dPmOu9O+5gH42hnLZXIye
owyEeiIHa3lbwTygL4Cc2CtKiMN0QLnj7YhElBxr05jLB+8UROL7siWmLHwNsgWD
hbPKnffxMqzFN3qAC2WeVE9jZtR5iwItS3DBRpFBLu0tksScGTn7ayR4cSLQBRYj
uwpYZ6RPofMImiBSbvlvIhLVggPI3AJW8VqEmJSyufmyRoi8AANeElkTXaXPJu1m
lHrfRK55yCArQbJRiSiUTk0Ptamrud537DHNVBR7voZkT9gzU7cs81AaaWYoaTll
E6xoJrO6wjtFcez6A85+wHkHK/7KJ2DhSris5InsgTEb0CvWXOY/Oy63B2+xmRxQ
NGZJ1dbT0PiV1BmsssnK1V7a2nL6X13Pg/UBWXFRFXN1qS4wNm6NPNvUY3iCyAVF
31FuCjueAKW7Nz6mQ9cPpA7TioKgGEdL44hkRMxxHcg/Ylm8U9kZ6jhGxls5MoeW
rhc7MlfQYYtYwO6/e4fOsWbejGASb0ghrjChB8BxkiSfe4xN1SYiDEUyVRnddTbQ
K7bsvwcbXR2s1jBmKjuj3rL6seemqeBAiXFCEr2OVQ6ivnh5RtPwAvBPvsgKWpAm
a8WzE+/yl9QvTlg5KQXkzx2J2xSIUXFvEpLlX3jcMtJjCnKj6FHMPwfF6pqvzPcs
ZCoZh8rLCNdkdQiTxmjdMUa+b1eK+25dnO1PODdLzGZocfoE6FUviS41dSU/9HiN
WSSTkMHVQlLhEVTgqFdVuWUyDxZ6h+SNBwU6s9ty1R74sPL/jBvsMxhq7UiCRb6S
OSNAM8dIH+8YAVjCY93Sqh5AWgU+2i8Kwi/m3oYb4mzhyx4VFiq9KYoOYS9nw6cE
mA0xDI1oU/CTpJl/g7stSpKrL8hopFn03cyARA57KqFMF1BP9IxY0cfM8dwtG0+L
A14jEk/HO4Q5LQf7jS5vY8smJuNiHTagr7Xr746s3pO/5tg5ZTGuAJicos2dBYhX
LXltOZkenH/D/pfUHcAMF1vssw1Ookyhgar/4vzab4uCfK7Gubx3MFMP6xXdx/X8
pZ00cPnx4utt2iO0Q1UH2T2/2dK2MhBSge5hitYG/ygBx/TJ+iLxBVRNnySL22zr
YEPREhsxb9aCoFAXJsDXPKfswmqPSIHZ8WQaeL750k6N8K9ZFAXiqZrA0Xz3xAO1
htx1mqVP4rgpWj5UnOSiKnnBDZOVIaVMqimvrCnIpc6XhAQpTmSlyyOu+da+645W
jQTBuZ9bTtu/8F+ZQ2t49wDfG0K6HNGF4KArvnpXf/0fnMVZxS5mYX275VwNHyq/
SwWro1MIcyOElH8ahqlcOKGqm7BRqP4tCCPxxvl36bvnV0izlPsO3aMZsI1n7aZf
zqwh/9FC8Yj8FaohqroOJzHOMr1r7NgpXIHKNfrVhZ8gwt6sd9MVcLn9NQ3cuCcd
kV2xa60ROUICvwYTnjuz4NDEH8HrPjn8W8vNWlY5PyOaQww2HeO3Qjy0Y5HKhRVe
eGwWDFfapcZmOeftnopn2s+h8J212VTkpfen9jfg9Qu7TtTVVNaS4vB6ulhFwprS
G3qVfe4CbtZqc4EkUUJXwueilJy1EahjsAkMnZkZ1UawWRYCIDkyZWg7I1McgPs4
gZDbzZS4S5GIqGmKI+JZoOoY0xCWM7SmUxvbNBfXbm6XiFtPHNhVYjNpDm7+8xm8
0QT8q+CA3tk//teDVjUm2zU9QWFsaofPvuOigAUr5IPk1PMRpMhwAPmUgvs1CSib
PPRJYy+Q2jF1akr05DxpWTFvzi/nnGIlynQzk/7iBMBw2JvwKpuz4EEBhH4lt8ha
7CVGGfOc90PyB9VyPO/8o3dcITvM8aM3OwnokUZsCoMo8GqVUZMpKndN1DlCbFrf
yEEwchb19bavMk97Eq9N0iZiznSfCL0RGd85eBiDTLG6+Hw6y7Hi0jGHRF6WQlX6
fICNoF1qRt7IF7xTN//KVa7X9oBC+I6jHHns1Oa4rFOqUM55A/eBLQsCrWUWPnGq
5tSFrDLEtLMjLxDtCpHXbywLJ1n0MBw/y5JJIHVQ2w4Y/f73zZao5B0nKK5E+oSC
Pf5J8bSomqEfES6r28MnLHSdEOD3/M8/2Vm/Lgw9+D7IduZyqp7AmSL+PQ7x7VDu
LkcdcH0wQRHaCEirOypJ6BACaoYZrDTYJUvMvxSSnbxwh0o+kd7E7Ht67fO9VjNW
z+Qyk1uIIwLQ0iSmmgFi6ZTYtK6hwyWKsWRe/pK4LRSRtl6bzG7eJ+/Rk3C8NKlx
ZALPZpoJqwC2Rq7HEOcblM8qqSHHi9yEtp9Ms3DoGQSq3VV0qD2N1yXwwrLrPjwY
xBNzdHZoKIK9tEsiUPmlcEtIOcrIBECU3OriKwO2gLiLgGH8UZO2OW1F4aej+1br
zBRXsVSQHlgPRHMe1obD2P2xPTxY8U3GhuAAFTuIxMiY3tv3ywRWdM2j58IAJ/9q
DeYMqejB+jRhUtS4F9kcFWN/SXA1LF9Zjx/AV59iMcHXKZyOrqTVUT2+n+ZGMaE9
nUHF1zXKon5o2Vsms5SO1jtQBbTsi4qwGrQEDBUFQ7xo7fvBJ4aYcbMGmszhNQij
FsKGjqCoGfxUVG4T45f7qTGxbtw3+gE5WFANo4kWH9gnHxaiflR/jojrsx7B18h6
Fa7dbslRC49hWayaClZvnphjj4U6BdqVsGJGHCrmt3skoUwDiSlP29XWd3eaFhSv
2QCs8Eudg5hdARvd/94yqwU2iHlQa8jWVY9riN5RZwhUztz04WR/BK0pdRhuLITR
abasF7J25hkHdCge9PV0BdfhS6kHGoCDuupjHdqTMDJgDE/Gb4Zq/uBKJkitBvFT
Hi/xIdf1TUdT7wrcpDHTNwuOr4ZRudkNZSUt8PbWLCqxBEHf1Yt4+q8GqVngEIi2
opK5r9xkvLevGEzKE8DpzUJSNOSHvjmMwwKl6vInQiZdNPcBVVRgMoVilG+u0irX
94RYWsFr77kFBhN8yPoW5pYq2QxgB7II4YP35+LHf5fN1+Zw+uj6VBPOCf4SU0qH
M1UNEdYCwkaH1+lqaNfVazlVrJxTT5prDmSKR9ln6eAjVKVN4m4xHUN0BZQ85U0M
cL6ulHl5MFN2rpyZk9fs91r6pUXPMih7Ij6l1E7L0dP4wHpJoiVP/RTxwSNCRd8O
Q5/SCux+13vc2dYan7zkm7cjFGW65qg4IGJvRHnVhEQ/B/6kaBTwTCfpUFWg05Yp
dLxsqqFgxs76DANooit2gUbKKPZShjwIZxsh/U/o6pqxIcm0CPPkyZdWMkFbtV+G
+4/n7ts2M08mS8SzuGZr8dVGvFNTTB6Y8YEhdg/hbD3EggXBe39KoQ+HUxSqiP14
mbf8GzAaac74EROxlWKYSmP/uaZEVNXzZMCoH1yoleJqHnHJtoBlzd6D/jhI6BSO
5HBPhowPOJEpHz85D6beqAJZFbMvFpSMOMitRPsRzDkdD3as70CVpXlGgvDQEsBT
CqX7/dQ3IR64/29udxTrEBct6l6Gse6u6eAtGjObbP+6bvjpPRVlBfIbSbzKDkyU
6aRal2Swz4uwjt2sa8MTcRxKQMZPZadGr50UyH2+zFzJAvfKSmtvMyeKBCQMDVrY
xYAuuvOMpKqSydK/u0b2ZxbUuQQaNt2H8Y6lm4xZkDPfHXDy1ehKxPUqSVTXeuGW
hBBQ3Pz9taiJBXlhPKqikZtYmUhA8GlW+sCkF0cZE/U6rTy0TAAXctRckkv0mTzy
aar/0Da3jKBSdfd44DYsnvsFGj9zE0VHbdwFg4gZd+Pkh3JXNI7fBwhO+kMLBv5j
WPduUPOVNe8STbkA90oraOP2q87qZ4V/+cbeY2j8gP2ktOxdFSRBUg9f1f1szoSo
GvjUbUl9ljaAxRvRjj5uA7BBRSKVRm9B7K4IawKtC/ieT0FZGUuoNtkjD5/LdlLJ
cLUq2OkBhExCKsVmIv6UcinUxdRfRztidZ68opbJ4ZhY6PilUg28cpvSMUzb72Ts
bu9cdWAAysSGfDLdy5iIvSPdlEX7H/wcXleUTK6qMokBzzUw8RqxngxM+OdqTe4z
NHHjjJ/Qg/zqLMGZbzRcOYS0nNe+8nVAm8aVhcqqavaTIHi+4OzPOAFf0jul9dQ/
`pragma protect end_protected
