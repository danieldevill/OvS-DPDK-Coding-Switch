// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A+44Q4quCr2dqx1EKbXBqgNTeWOSEJYwVCJShpJskWMYdJ9F7YCqJ/iq+AFVzmgQ
IGyVpow4pg23K8lsaqfrdS5YpATQ3SebIueB1CDlOfoQ4uFwEFviuaHEWiJ9SiLF
e2wAIhPM9YlP6hmEv70rsY+NTtn1uzrBDNmd+7cyh+g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2224)
53BKE4jV1o3aTx0dUsz1xsKwfjfn+99Jf2Sq+8bq8j8kwvNTgf19QCYV2VdPbcnA
N9Q+gTEeUPYEfp+wNvL41sQy3weUmC424SQWiPZ0LK+YvfAgGp+d+wZWHfIiAg8Q
GZfNYQLHUnCvuQBn/ytCUz6x2pn7q8hBaxqqhz7sFbA+mQFfc1alrySG6FLSRXxr
R406R5azvUROIQzbC/ObaegS+uPHIpkh7ggdsvVXMUF7OL9eI0BfNsVBbfXCbzL2
4LwFJnKxNer1ybA98uvVZ1b6jBlS9JNY6ZxUY8926CYOwVNQv6Gah5EDLSpZOAfc
E4I+L0QHvcvV3LQEzm33dSS8N7/UNmHXKfgcvACz1N3w1IrJdclMR0JNAyq6M33D
QoLC0Hq2U5Nqg/qPfDJ6/cBBcJni7aK+SL7kZOrE3tFDB0OB3bKBlu/6OIZMMMrc
NVNrcKRZJDdIyv5u+7dGBwm4fB+STBIe0M9JAUxgMem9zjSO0hbfID4h/y5OYgM5
qaI+XI5nrDnpZRPVBLpi9Pt0wmxTNLNtfgQw9bSykh+PLKv11dISW8k/e9s+NgXf
ImsJrcUhzWpXo0hLAxEQDy2/aBLj8ww+g8ghuHqjbYvMZNz4e1vzqI0knaC7TGCJ
KajSLPUxKG5CfJevy7/GkmxpMyBwdKWppLL78HvnegppFw9fQAIGb/a49mP/IF/Z
6mh3Eysb6QMzQQGFaEallNxcTfmRwgyGyUwtT0NP6Rk4sy+qqnqLZMsfndTVWi63
XAhD8Wzx/PIpNYytBnOrL1CEDjj3GjqpCRcoZ4nlTv4Am0dmDBx359qmBhhX8YR5
Kinl3+DMaPb3oxOWeCcMQBVYMtcr8CHLwUOK+2qqdIFc/6jywOn9kAH4gS3VpGBS
WpW+ztAUXAsbJT+wdRjhSgElSwJLguioXHrw8P1h9vCyq+N6ZNcppg8A9hQR6Mo/
ORthCiPkXNC/87IpObW8ygNrhSwrVwoARfs0eBNYpxIBeRyWq85ewr5tVwhmxqSq
/yYAaJ7/ovdsHYJA3qtdV7lsnHdXwDYieWej71FknHnA5ACu5ETnfMxC7WjI1w5N
y+gMqzakRPuNBVBYCa9ryOuEWAijAluK/AmNS/jyFAoUV1BpyrdlkTclqqyAHwbd
MKgDlZ09khaQQeexCzWXf/NJFuVyypvbWHKWoBjxjll0+PjlcJrz3nUom8QImUem
eMVKO6OVrK8/71tEBG/wz1wjYrUtkwXZjx6W5eschugz/dcZLigGTXxTySy9FWUO
2RaU3c8espij5XhpIDL27wGM2ntQMvL+N5+MU31WZFbTnIWkCymb+TkzroUbHQNT
Uv0cOFnfExIcvL3ahHcbln9VVcHXyUICtKCogoMpYQEC66MZ+BqK5352AXhS+V7r
oaQ3yEENi0paneq5hV7wkkDFe8HAJ2f8wFZad7i/bd1GPch/MslJIRPRZF7phY4t
LFQB/U30FWED3xKiQasiPxlX3cSPMWh30vVGYrA8lX4tDSsynddOvQwHc6HAdUBn
LnMRALbuIUiLlk/BkTasR5aZ14oXqSS9eCNP6NATdzp9mNjTPbqiJv6EVUhNo8pn
L+HrpSj86zGnDqu+7VItcKeMJ9Shf8p0kuth5pPwYD0d/VvVZy8TAZsl+sDJ5p1Z
jEKm7//0HZLu82OEG06xT3Wvr4hfVbaNj4+s3Z8PEjQRQJfhZC9uOVOJ0G03822M
zO6aWlv1B69DV487fZVF0B0Y2sszuokP0pOqh2qqJ0ynF5DVsYbM1GkY/XlcDe3O
Xb4V1IWhvym9jKOTnf3/rPOEdwMeQu9yfaY2brZ0j1cSNMDQHI3PFBIplXR5I2Ef
o+OZAulBmmIxByKGOtBpYrr+tOyY7OLfXpz73U8Kj1LUBnVpmXvvTW1lF0ix2QU6
KLdo0/0ebzPvPZE+9mbE57J/h5hh1GH488g4Xj4VD4KAKj0/bDdRol8AR8rqUDJs
HNCwxUdkuyS/nOpTyOBy8U7SIxF0SDE08DjQIs195rllEA80vv9EHnBH9BYnmEeL
k/F49jVUej4hkn99h9f5j29qjbyz8+nZGfCEIzCQPzTbZTj/XA2FWkwymQx4OtSZ
fTI/YJmRaO/BwIDAbwAxhmdUajx/LR/3+FUBcjPJhTeaUgZyLfaQhj22j7+0UhHb
hoIClIqzKoTrD/2Rg3Qf1Cmc551qhdoYg6GYDdMmHMV+cOpgagenQi8NI/R0CNwZ
jSSZ93t8jvV5PemuEIHQ5EqoTKXy2LFq8FgtRLyBlL/eJug40aEttR5ghHOaR3jj
hzvMJpDLf3S7BiwVKxgIz8Lq4AyjoXqrLMgSyYf8RKdxAYBZAqNRgCuKIM6tj8j3
a26OH04sNu3630ZdZx5EJmCpl5NnHATKkmfKlYNF02AgUz1LIOvBgZjKikRrYu75
j+sNIp7izZPeCU1nACvhp8bW6xJ9BzrVtagyCiU9zeNwqt+jdSfM105nvhVHZ2FU
4OHqZ0PqWVAKAHEv+PsxGBnxad/SCNfZtnrWP8IeWj3c9mQz24rLwzHu7YcsegaM
4GOPmbVZQDlKwqJKl4OlVlMXJJAD6xE9r0UWjNH9RCVSMAYdBz1Ow/uovoZ1K8cN
qpcimoqO4aeA1+d1+QZSPeTsoxkIJRmi3yHspo2IXR1XozQFNQcf2oh08kNAtpUE
A7HF8l14JFYCYwPhVfjxY04ujqsorqhIDu1AvfJhA1DAOCJJsfZFfjNVoBo8MII/
gUniMhsadFA/PmfdwtZbDVNmyhilC+h+lpOPqihGbqw3MeHWXy0e45B8F/Q6f2Q6
OhrrftvJLqMjTkHlbMVc9jwy/yw84tS200zWV6t6haSJQRRqMsMppigp4f4EMuGK
bHca7KJrxowOR36kiKRCfOOvMsouH/MxfYnmgRFsRhaRESn4ps1lkYxHZsu1IOEg
5s3vHvDB6+84BIWv3tPzOw==
`pragma protect end_protected
