// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pe1wnFHbgDploc9IS1a4ufAFHC43S6mWlrIF8oReWFJrZAePt8QHPozrfDk+wLX7
1VibDo5ip1GjUh83qI7cxfOO5KAUlnSyOtS5a4qxF51HMlgySgR1IFoMUgV39qVe
eBH5cyl/ZfjTdEa7YL2Royls4KoZfYOqR4ufaaqVWxw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34464)
k5sXHu7LK48//syKUQ7NAvd8EGLod5EjO5d+ql/8KuK+T3kOLWW1IM9wx0Mh7zY3
xkfNwBRbHIVH12oITnSFx7dTASc5nQ/jSBtPmc8PbCTL+khQFirsnHJuXb99DsRA
PqUa848BnS5vHDP7CRpDY10ixQ/gMfU2iG7CGc65YXRTb29IxCl+5cFyjIVSE+Vb
+NQUuKHfoia+brI6hbEXpHpdDSdHzEqbtwugdMyOkMD0/5TGbhU55EMsfPofCcli
r9XTksHp3Y3MSDObuGQKFhIVi2icoJxSP0RuV25iPn3CKiFhbUXH5opIIouKYTCz
66x5xYsCANh8rwJ1sZogYFSFWXdqgW/trOZAcvdOG4V9S7sEzLsmxro/0HlOR4X6
KsCfp+9sQxaz4GZZStuaFl3k3FE8sWLFbm6XQcGtqCMe6AmVC89QpatKI+R61rWe
U5WAfIZiRkw1b+cHZ62/rz/8ZX0KrJRVBIeStLo4gOEQje2NycD4aOtjxW6+Tct0
oolo/xqdoyaHfNangzzZcR+hEy+U0u1HkNIZlaH/ErUMYCg5AOP2pnfd9vtrOvPy
7Smmu1wTKfPDCE77Oy1CjfCi7z6j+FCt9ZpJ216Ey4KTDPKB83FLLPiT1EMfaQm/
h7/36SCHpuqYGF0vOFHEpXBhVGlKrMQj1/k3zZZLTRMkcAiDhK5HGITLL3bggoev
cGFLD9rI5FqG2wsmQgmtb9Y3E0pquD7xbt2llT2PcXC6OXrTAdDepBcaFgdzACz1
NWK4q+J/bFCMYWZSLTQY82SVHmuGzCq5CID0pAK2pwZXD1MwkAbQ45NX7mAitx1H
U4NA2tW3j7TV94e7vKgjDNurBgyJR0M9gC4fxn9k4oclNixsUoGUo0d/xLn2XjJ5
6rsipwTs+iv9IcykdrpFROtBVotEaHyIBMD7AY23aRKUi+MxoagvN9UyawlXvHlk
ZQOjohBExy4Uqbg+UiWCU7wLEurgV22Y9xdH7PX/99i0fk8lqhRA+jMj3yhHggaR
FXgOLDHh3eE3uF5CUFsqILU78gB+2RR2Y87ZRIhfDq2XkKxMea+JRKAQki7XVeSs
9lfsgGTiLYJ3ieGEEk7uefWO/8/BNZ87yo1g7o+b/q0g2/l6nEEYDcLqYSLULQhM
aNVweXKus9jkNbC2kXUfraGRmjNZz78dooqA0cMNjrQOKIRraux11FaH+LFMPJQ9
h8ulR6FtWAyzR+xfDzGWnym5/CIJqP2aeMpSPPgDX/hnffj4xzC4SBzNrofMbuC8
C4jomR+Ft2i4ee7LWkxPvsrKa18m2koSexUMIhPEaVAVL/mxu40nscetgg9nhG5W
egO3E4KHYWke0SLGk6i+ne2ISkKfgE5A75HXeqU4Islghg3ySntBqLiY0XApNLIR
y0ZK3XsInInirgXs32CtTnkLFUcmgTyndqkLJQGoiUATrGtxGOwGdQcGymVpk3tS
CNQlkzkgjWnn1tmjMmSGuUgoekou+bZDRUnsUsPPJ9jxM+TQgIYKfFUd6HDUdZ8U
rtrKpoeq2jalQSg15XPLqz32mTVrNGY3o7qNN2wpeEBQp3Q7qJxdY4uxfdUHLzOY
6HaC6qDc8X8qIjeWJQaol/18OUOlRelETnb0W46Qftd+wJmDepnx6ZccmjxG/MP4
99gU/l5jyA5l5re0dtWiLbhvGPaVrIkhDoYwwTJNYe7M9RN02IN1A++uqUnwyMve
de90ibFYdS+HPUnKgezSOuBgvaIe8644cvENxHFvmAFZZCmu38baUoWq6S1JGxan
ZOnate+Sm13BeZgRRYtKnQfUUtnuziEuId0bekhad5VdZQs0HbXapkAgzAkNSFZv
n/gN+SSFnTBqhfUE3+mm1nnL+NAMk6DXmIK0OEPp2j1cGqhoHGENFQBc8J6wZdJc
qaDicQcdLloNm0JhzNapU4EV9I2nuzKDKzTngCpyqLgUopxDI9gCTtH01jHadNd2
so8k6s2RyKJmEXwYdKs2f/tBjRSNN85eFG+w1LmhFJjy0tHh9HN2Iy+jG5cIo4XT
+TMpMeyJ/40CTix8EMR/E4StLin05rSEBE5FHcf+Dd1FLWehrOAajP7Al7QdLkY1
z9l3dG9cu2WiVAacA9GaifelvIrYbb3d8Xp3Wl0eJWwVaUBlInoIZOT+ywakpuf0
cCOPvPmB4ilL26k9Ati7Ld5TP6mDW7xIE3P9cJnUUrT4FtN1BFX/GPRXRaLtyYvG
STroHLOu9b+d35INYrAuC9FiuODXMganpVa+HKouLcg+dBtCE/28G//Q/RQBTJso
mmlRiuYUJ/dJjXVuTcaCGsS9i5aixAmTxmw3u7Klnq4jZAFPAOR+KEHJAVbQHgD2
zh81f0n3bHtU93PFtKNTaRIMs7buWrE6aPvfuXRAZ+H/HmCjK7/OgSqRL+mqKcQw
3WYjceAwm6/vjTJKKFk0bMsS//IoqQWNAm8pr0HmFnCuaBuTgom4i3lJtMQQFrai
Nhnqhg5SAIVTkx4X79cjH5u6H9B5BO29n/ZtPLg0MoWHWUbZB/9Xwk/v/lRVZYe6
+PCzGxEFbPuWz08Scx0B2RvEejDUile/dMPRDmOKq5bDtR0mcfUeuwZTPYqnVuaE
7b8KRvNH+3PfArGn02Y/oPjjqe3JkA1QdGdP+CgRtcuyzB3BNR6OIn4KnA/tCkCC
O+bf8xDw4immR8Tsd5uFgF55xkfnMaat9N674f8yxsex9Zhl3X7MGBFFe++JZuHe
cNg/cjTwdutscd0ECxgOIgKUWANJztBwJOIcCMiQeEgkc7/aYVXY+uoTUGQTm8as
07rr9Vg1lDNWxeqzXKabFR5U3JDtXcNESrKdUcNAyBmAhRineYGqLuD+whXEy9Du
Hckw45YUhVkhUat+30Lx0F4Ozd4C//8DPN2U9w/TuKsZE1wANAK4lQiGx8qOorpW
uRgQ07mz9Zdavc6lQzh53fPAf58bfInvXNemaxPDsntFI/SHKXwCVVrJx+FuG7RV
2zAOIpcF0w521vuKq8dEemS6HBzDAN06JVp1FTSS+dqYU8gz3Qm9XIBg4fMYsOFY
U2Gy9v51GLkcl8UTgvEN+ooBjInkmc5LvmgdB7Va+A2J2Kkz9obOxD9dLp2uxu7L
Bs2SICNfFpbZyuXfROQyuDnvMiiyf3ckoEYtxltCLQkF15wY+xWeAFt+8HMKgWt7
vpjiDFMgYFLH3I8f6zcsUd1M6REW3dEzyUZkPnvwJUIXikTlWAgHXghuyngJsvlq
rHCH4DYeI/AwkYVXZcGZlJBPjXjLfQRNGqQJoKDZ9bMpTLL/HUcZOGsNF3oiOtjo
gfTxsIHZDXvCR181Uu+27SXNNh/VaM+MUG2A4mUg3wGmboUZYAL//xtCLoOLQjGF
0FEagVMyUeAv2Ade/CZFJvE+B5stVWjp7X5zc9QujzCZC79lCc6x2coxJJ2vmDsC
Fg0P1FEmvd2GNMf4aYeLBDH+EQ5d7p7WH/qD14FgwKHYPKtXvIiZ9BCOpLLl/tl0
tcGQfh4aR8f8/tpWujFujN3r4SIeAz7mGTcgi9uWhiqOgZ33u050zFo2ZROtr/oa
Qwq5ZfPHaLaEioj5CuXx+PGuoGd2yyNn3jxcNQe50tKh+JwVR1DctJGsSzDYjubF
fdIXf6thxVQ/tFnMte8qShk4rblCDmVd7gQda4KOAl7nWIziPDp5kPifQ2uVByPt
XSfOFmtYPKqS+x/HzlhFhwsbjC2dZM24lRkn1xFglRb1r52c2DcwjjlaiBIC4V53
teXWB8FO9biH1xfMOCRs1t6+U6OL9v0esfTgc7bD6Ce+JFIZHrQT4MtLnrRnINmB
NX0AJ9OHRpgacPz72ZLR6hJ+1QJG78qcEB0ml041G59RiC1TuUSx4nfJ4/0Bi0YQ
EmymWZi2h07nwswt3hCdx1TlWrA9CYoizBlBa+8V206nyph4bdEFUXm1S9SOJmGM
ZpFOYcFGC1/TYcWWHapWPSk8lF2vEzOiJYKsWJf4CSUvAIpeQI12U3aKFLdMMszj
/SwC/kfqQhRP80BmLav3Z+AhsOYSicb/+wc3VFlfeY8Ef66sR78V4uNr9TeCXl1E
bc4alpfLH0jhFlviqAg847LGMS5y7W3xPy0QpSeVvlyczh/saLrrPrzlAOuJS7m0
0SMCDb2wmW6elp6sggv2xMI5ExA1k3bcMicZLxBrLc+OalAUKGpOHnBPrA9IK7Ic
owLMz4tFqjdBQma3PI+qBiXT6Sa0559MejgzOdov616tIq7JETdOwsFBiMacOTBp
wIgBRVGZR0LSYun/eG3OWh7t9jhoTk6uNlMEjXTUt1ULmYX9NEylWYZqDtJgOy6h
z1fWbxItwcA+/OQE3hJ0CHkHeDWZLUeJVjhksn12WJxN5DlLJtX1adhO6OnJt8p4
5obnE84OJfl08igLsyhSt9xdZzD/9TaXfbV2Nsd//2inptFapPlw25J+6/XTCrcl
CnyNy9LXKG39cXcwmhNQRbPUhmbiKC3+qTDfTUz6W7qxLqxcg+bBzoVk/zigo000
LBfIqyd6FieqRy8kFxC9Cp3PpIZmuwI/W6tw+mRwhs/pERKcozLJbS3RZtXL9S1+
VRy0JI4sEPO3cVS41YW3Yhphqu5GnabETvV7PyisBtzkXp5wWQHKoocFd/dE36N/
i+PYGv/yP6VlVFnvEP4/In1Jun3xhO85sQC7cpEfX1v7yRws3IEckB09OlrovDEG
1OEMi/QmckYFPwBOWirM1NoRh0id4pclsGYqeNR9tOCdKCZq1TX2Mnota0fW8+9X
WMeB5iJ2vAW9Fy5qnzWzi9jySGRXTiSERNgM2bLDcB0feBzZb7MZxMI5MkUhB08X
qTiFQcBFMSagO+iP+osaeBjUqvB3p7b3VlMW7gM5Qv48oXJpv9EGj5T2z2mQ43S5
3M1EaFqEX8o81uOA2d7ufxkBv2uiifBhq9/bdqqD7it9k4sSjdfSJHpgP5B5yq1Z
8DTf79ApRBwCLYzLys9sJmIeeBQI5dPn7Cs2Y4lpHygCTbxvz1/02ShzYV4nkiXy
qzY7BGqLmmyJ6epFZvbEsxA/qcWf9or/2BIXIASL9+/LGeHlf2CvM9acmAtysRBV
G8Oiso1Rl3ND5G1Zjs041DiZfo2gyg4qbqpqaFXq7qORP2Xl80ACdhghk26XvdwU
5RMcqOf1jnbUvK1QtxUxJGAtMLW8ipCI7SL5QZAFsQW5up+gBCgDLyLr5NvSNegJ
CHUpasdWD5qXXFof6PbEAFhHfBDkX8MWLuN1tsw0edFIT6eXZ/FnyorOkslutgf7
VfoOkaelqAbAVMELpfYH/rKMgns7s85mUKqpS4rJY8ZCRMkLSFDrUSQhrl+kROqJ
JrTwRLu7kH9qRxQOaUAodiBYI0rjitxHjnr6yAy/affuJv2tXZy+rOBAjEX0ikXV
/RuLuCv8LMs9JiwPr3oRhilfe2sL3QldvkJz1XbrRq5fyoUvDtbJxsKw21DpeTyO
zi/TAbGC7Z+3DXk6Aj+FWTCXUgQDRjo2NHY1YOT1HYv8H2MTi+OSVUoG/8paD1DF
QJdX1AUZGjQlobiP165ujzDGOb8Hv63Hw4dA0lt89+sF9NDc/6RPTPxvDvwf52OM
NnJPZ3UnZ7HyEGE4H7+TqWk/zi2vEffMWgWw+73yaTCQOhZRztAr0NbouDm5PkHO
oGes/m3egSzF3hX4ahvlEXzRmM1qRiwnVVgXorXccRtADU/iBr3+xZdWMun1X/5W
UkZAv+74gGcGw1m70S7tLtegjW1GkbJJfHgOM5K51RzQmhPxVV0l5fWwyL6l8WzS
1GtiRXq0TuWVebqBnheRt98D9didngdkynYe+hdrfzLROSfLWQ77uAwtGoZ+wJ/e
9DiVFn4kaKnW0EqvimLK6yDL+YWu3UALiEyfNAwxFCvuvpxiiAupP4Why+74R9YB
uR0bvWsE0HxNMNF8+nPWyu383VWUZp0mSPrn885P2HiqaOa3vTM3AtakfE+fOHHW
0qt5T+cSvVNSRzGi18295K8+lL4GE19TGzd9QA6SEs9txgRta2Ylf3xyWt+rILpk
YtjtHoyFVKahQsbImsQSOh1nperpfX6mE7K+ZcjNmLJ55kJ455KOHCQ3l/6143UC
efgyQ/QhJnUqS/Co7quzzvMYzQ5iNIXq5AjFJsxMbXniBL/vm+oWh9Z9wStsCxyw
KZgIDChl+kPcwYQdf2nGN4zMcR4nUYf5on2IuLsImhs9W0epCOhrkp80QiM+63bv
vcS5zZS2oXqcPD+Kj5I2MOOJwown6SGZyuPsJ4MPU3+HqKLV+uZlSLQXMYopgFQS
JFcwfQugNTtpsbcMNwtIGL4uAitzYE93x7mxRYHLO2IflZfKyoagjtPesThqM3pH
iK1IimQSHFTGNvjwHAsgNS0ujNZjb2AFabMaf0n/ZkB0kED+978rGM0c9UhhPO55
2DMQ6WShKFL3hERnJL2B1+axzrtr2L7wYYtlPKPVbjrPN06KhS6vVDYh4bATootS
0ipm/EwSKhBP0E9wgxbBWbuHrRFtckGYYYi8fkeQiSkBCk91czT9lKQks+DW2XB2
J0RR4AgmbKPtRwXCKPkeUEzA19oQROGOUnsPaLQs7JQUuOGiDHgW3IjR+ZRzcUGi
1Oz939ABErYPi8qWSp1FNmBJH5FTyY/G3nOKnlcl3IgasY2gibXrskqm3dv/ZtER
CJQIjt8BNk7jyMBYOkxJPzZfriVCYjOPJfeIt21cG2jyupx1kmEh30A+V8Bkfaqn
IUntnzL3x5Zzdg/I24v9GT73DLMpiteWYF8gdaH2x4GhxW1IKiff7On11Xvfa7tT
EJ+ajysIlZAAHj9fk+HkZ1xSRGMYSj7CTNWf0BGoq9XhaFf3gNiYlAwK15sjPC2Q
buqoBC1lYKr9a7raoRrhWiro/bBr55Xaz47CDs8FBBhUykvyINdGcUqEE62PSTAt
w5poimG0M9YBDHTjQFc72j+nR+GwY0lV8jqTohk+lTybkLPgggolT9cWYIPuYEHu
/4XEh2BswIK6Ylq3UwNS1qVsnvPDvoKLJYVgzOqjyYVfehRNklpXsE2GjBGO+fW2
4ni4i4aX/9nqVt9xdPXMuRH+cX4W8tBWQjTv5IHEa4Bv+0xhBy7Oug36OjIQV3mu
6Yq35WcRL/ObRAbHaDoWE8O6cCfEJQ812rXn/pgFY6vPDt4O+Qke4JksAYCNLgwt
cLJJwJG3r4vxJhzVn6ZKk8VNDDMqWWfI7uBsmRq9KteGPZH+C9aewzJZiw15CJEe
Wj7FrYtAKPqBqslN2jLmftFMzu/YNS+E5g+knbTHzCrqrqOabn6aVzj++6iGVv7I
JCAA3+o+4c39AB1/fbobGyG+YKdkioo1djZ3cYaNSsiud37Igc83ZeL7SCUNNJtH
ZZ7iIdwNAzt6MtchSA0qG+ngxzbzMSSrGgcQQTIP4lu2okT5Ejnq/okaisb39WA3
u6QkJhgghAG33wL5UXuCoKTb9D4eeSDm1xqF/rPKw9J2NUXQdtQXsm7/GAoKAOUk
ECGPoc6s6+c9No7Ivl3z+qkc3UOeONtvwGcHUQ8JdBiwierpu3NKkZtOSqzolxQq
c+yhhYmHW9RofjvPyTO/7pOBSsvLMGJVtnnpyaW9I5tpAvHogZEz2PLFTSocRtTY
bcOEBpafFCyMAX63chPFlpUmbn1DjIofpT6bBxVMERzzvtettQ5ess/bxkAQLMfG
H1CVGdWnnivVA2DhN/7cw4s06UU2/3fQMs/Z6pTRO9g0OwTFHoNDfLo69yWOxC7u
UOuraHPdvEHxoSShj4T9P+v+JYe6QSZ2B2foO6OXECy+OUYNFaCU9QVlUJXOo8jT
zjgCHPdqJtxbTHdgPKef3yd2OKeq8pBSBzj53D2vtBOvUS0anZF6Eoar4sxTRhzs
0vuMJaG+NNNne1YOqmo0uOHW3RewjD6tMPTQzGJViBr5IzTDiXwBRO9pFaokBj8A
cbtVSawFZ1l2WHVLbDAIc4EsPhTD64JNJhVDxv3rXh4F4e+nxhhiSp0skQASgzE2
uVlnFnvn950sQuSuinVypx86QTdqpJ11TT0YzWABDz7S8GoP2Kl8FfKFuoz7H2Eg
zzcFeBzqiK7pUUET7XdtkqY0GBfyafr2k96TjFFVADGYtewA7Jg1z+Zi5M/XszHo
LcXpfy9Qz9XC2yNI2aoUlXw+DIM99UB5M0VC+GLQ5KLaPHx8OBIAc7s6Pl1bu3qt
6Ul/UCEmXbJDJq64RZviW3nhwk1fDOEJkWMIJZKq2HA/lSF3BhgNoAV/X/mOPfp9
FLs1ABrwMp7gZN+PWAVkvL1CUvhbP2jrTGI2I6XjUC+urinwG64oF0jJ88DW4Fgd
u/4JGKfSpSv/xrnN8tTk4UAYP5/LlMQLg21r9TetoitBq7lhym+FqKYwjng23Ca/
x/GwzDkv7d5pooDRZB7mGKcC9d+2nQcmpykAnwWmCak/ZOpUROpgAPRf8L2+j6lP
vXSiqam5Lh/PxIIW6tz3UuZ0mDadt01CWYzar6n+he7jIq4HtfGnOgHzgh+QtW5e
1M53bvXez/h9UlZcMlahJ1vr1dZmAPGVswsiVu2ZeNki2YdNjGUqRK/CEqglkkO5
o2Y/+v2iTdxEiZYIPRqHYC/yzwwMPE2WJQbKDymbO3UfJegEr5kP5OMUSXDuJp4y
GvhziL4pWFE1GWb/SPtpIBVgbhPpHlvgMDyscLDnueMq53ki/ceOEHJVudbQ+rgI
9DICDbZuV2X0hoVxwVyScHHT8txSmL+gB9UBllQT5qDYZJM/JP7mrEEEkZ8yjotM
IYsfPyVM9OkumYmxoiBDlYPfYFUvKRQx3LVKRB2Xm1b1tRfJLGXN0bpudxuLKF65
xhWxNKvSDK/L1LEmvexQZVcvkhSc6c4IzkhoH6NCF3om0kXwO4YdrpgeUdjyc85u
pK1DKwqJxxMitlHqP3WR8/TCqCVfSH6ukx/goi4Lp/mbcTACOExa5JTjFek3O427
7SU037hO/zlwST3EJ/mOtUAgMGwkE+qe+UwKQNddisybcpAEnHurOU9+OONsmJcy
kZlgSWt/Hyj0kTW78NwGNJu+cLFEUn40ScJtFsB9676Y0zgKII9hCHLDxI4nmDiF
cL0fN3uuJl8Px70YK5uCZYIC87GNQzwFuShObmbtM0YI9mnXpPSTCnkLqjpdARc2
H+KszK47tL1FjnsaYFIqlk1z6yyX492VwAfzwlbEnJH/Av+QGS4c/Dwrh+Ta96O+
vRTbLUEH5qSB5zacuiwTygS3KWuc5Lj34pFO6iIVF6APVamv3GxQo9XqOeGTyJWA
Osc78MNqYfP0pq7hPKcJur3aHw/GJ4LD8MZqkZKe2dUDaQzvYD1ah5/rBn8cNfXS
CB+B/WQs7EDeCxUxBIfAHGuQLOMECVjIWL3Ci4KrsavP3EIksX23niQSxdbiebos
xt7W+C6Tk+vO3ZOX6aPlZaXhZaFrVZspe5AuluRBeVFoqznq+zkc3FVV3cQYdw5e
+HLGkdNQIDqCb2nFa9aF/T7mX/RJcq2cLpLCANuVuZAFCc3XQP0yJRpJpHw/64f/
IH0xV6Q6XEwdUyRY6JqCJfGNhrNmBYiKnaJBzBeF8lNz2HqpAtSxIyJTHXrh9Nxm
zwa+J4QFIBUA+JFIwd8WLPVstH2m+s65JlHDwUSy5pAugrkUt+QeclWbWbYfuj1s
XuC9Fc/5iE7dzhf0qv440TRTUSf4NdWkTSUjeMO9oFX92I6a3fRkE61CLnvOgOcV
sTI8Jsnyn1Zm0nqhu5E2bqPCcCPfnIq59xH5+WAuzA7M9/kWWjdPB/j3br/X0hak
Ks6xoGwB6HGdi/ze7CPXbFYRkmx7RtJ17fGtTWLqMTi96hasM/A1KVTBaIJFl8vn
Mqnnk/JNOtpotL/ym8M+NXczzZjE73isI80z8o+qRbOeQtFjm/SKe9lBnqf5hh4p
EDOYelIzlt8r+qahIquOUjAbNQlt8EHekQxc4yGzRW80OSC+yqRYhTz17xx+Zo7W
yOqfPtNNGHPuYip7XwSaEDHt3gulhGaa21tc/MlbReqkI9qOZZuCSPmdlhMxKn8k
1RJMkV+qm1RJwO4KVMI7bTzbUcTB2UzPDha7P5A/QgTEeXtTOYswP8xLbvhkPX4M
JYuT8C9L4c/9nQvSO2La3AQSnW2qEZcqTbZSdurGOmvAoLFfAmKUQLU6wbYCmKw6
dJnCvcZ2LTP8jEbG/lx/dXqJ/YJlGtvDf19/xjsjPBK0zub6RPjZka2YRHMc/X/y
apk2gQ9Yp45/iWIxtFWD4YCoz4oRMeb92OGhppJr/m7TbgWWk8bFACKaiZ3DvJDH
JsmnkkwKxknWST1QQ90QxV6PNeE5s5d91OUoKJuibDu+5AFqNHv/i/FD7GtCjTXO
8y7sFcBzX+0V17HeEjgJCUpB+7uFjplPyXxJHDmUXWErCutDa4jmT76sqOsuLaRV
1mCygfEluDD4iV9Dij3l+VkOKClcyCy5zuMTooM7NJOoUuQwfmZOPRY4dqd0/6Az
aaG58VxNTEsARRY4s3DlIMUNPx1ywGRbwRSSIjXf2Cypif4H0Uv4WpjvuWBecD4M
AVbvifsQA+28yufUFBEdVe9ILDu60JUlD6w+Z1LmCWsZZdQss/2ESYRsSEMyHwJ9
aZzbayQWpekQ1vgs8LZAJq7b2pIUKTjInehkhGbRv7gfNF7gbI6myXN9XFzxJEnA
43LXsvifh9X1qzz8QvgIWT6yUzFbjI27Bmdc9upqiexYk1Xw3u5tLPYuWEkE1bGy
9BrKR8QAvoc8zPYYFGbu7lHevHrELNRDw9PwEGtD4SCYmEH511LNzXssw9uLs1Hv
GCITqC9qNRvbeGOOtP90ip+5ZiKwga/KKHK4a0G7i48aL8lPEARdwQDsVBGTy/JN
RYAfgfD/7rmqpz4Khng4fah8RhSSasjhISrrfVIPyWT59QAN8/acygEcnyIGwciP
UqF2QZzjSpBKdlThgaYqk3CEkRZjcZVUVabiGWJgUA4xUeV30W+kFLWXKYwVjf5z
vkspYFi6pws6fAGjtWtFpTVHNhZjpg035javDgrGreEgWZws4lCSfDj2pZydTHLD
HwUa2ZqBpUArwaeOxGxO9xTsMxWzwMZVzsTgruGOZzO0jkBG4pRiG4CJDwKO6vjO
7TDvO+aVvFIVzfpTkVKrQQs2GYunoMbCHuiMR733Aq652qkGqO2HiS3Q9cYyJV++
F9d9uxCfilomiusTpaea0U0XkBdRAnbg7HAzTgVGHUi8g8BY9ICJJT9ViVPzmPes
9yS+DnfHU6hAX2zzsMdybMghNlliXhgWw4aBosFwDeLVykN/MJtXF+ege08e72cS
o2Xn5s1RVjIvFzwOAkZMW7RCnwDKGWfkEGyCg8Mn2YAKyPdvhCwEAIax+4KJDmxe
BVyOUQexO3fL9wK28ilYI9vSiD/hRL/a9fx9Xu42YsedxpARuTwNYpImUmJLAEj/
oaHn9lqAZP9n6/3ta5fFtJdlu3kB/aKoUonQfFN1hDMU6MvVgw/4ZQFF57zFxiAu
5rdH3AQPCQXnlZXnTKk92mGJqvE2QS75EPPrN0MKIYnaULwJVX4JQdyuQYMgxkks
wX4HgiIOKJOCee3R94WVRWL606zOQmN6IUaKpQFdOJMMi4a+X/4aupNf/LZasQV5
Bu/3jQW2G/KW6DKLsLTOv36vWDpQ+iZ2GSpSkZlwBDkyPO76WbIzKyIMyx25cvA9
MieBfX/drXwJ2OqnkgkFYgnIx9efwEpF4WgSOJzyFM5q4TLsSR1F9AFiwrvPGLi0
CKYui3RKbHXvBImNQFW8qXIBgQFWEU46S3MCZh1w9kAeT60Ppy6RMxECW+McOUv+
Un/xGovooqTlNgE9G4Wkr2alUMH/sLeL8PsIFNgcU8oWdA771NnVnwC19p4AmB7v
SreLNiW6AfrHUhNT4iSVOUQpR3yfDhhnbtE2TF52XMUm52juAJvFKWO3nVUzCzXs
XnngQ+PZxOk450H9+hnqIjFuYZVWrUjMYvglc10bkxG8NjESZO8BLUkcwOoDw76N
eyw/XrwMaWzXCo0OVgDnFQ2/+GU5wfUsZccnk3m4mfpo62eLFKSreRQVq1jOrmw4
fZz+s5HyrwC2hldhkRwfkTilSsfoPxXNlboge9NBXCMvSasmP25dzvEZV5m+Db83
i3NbsyX5K1hk5PQdbTdcPmUZccnQaSr4U7UuAhMclmQA4R3FgJAct8vJFFOmEZ9f
x9DSk2EbhoF1ispmaR+B6xyS6IgDHy429E5YTPHp8W7ueQUIZhEizdGMYfIfyZr9
IM95nfidmr6p7mnzYzTKPn8fS1UPxdwzYz1HBcnqq2ToZnHRh0nyUfIcg2Fl5H7R
zzGdzFxO+ehkcy0wouM5gQ1FFjE58pjOFfVS0ZniX5AWJGapvvvFLKabUHMPtFPB
so5fiQxhY4yKiUUemFAyRK66UwaxvxekXPUCkhDDM9MALaHTfYZ00HhsF+mMP8g5
onxmIGPlESO9AMy2D5oaXAFCZgiXHBqxJqKhu72teuAOyGKtoq2qZKhT8MHB1lCM
ag+jk8c0ML111WRGKiVPk5ivTXtKA4IdaK2LrohATQHHDIcvVxQK34GJxW8oKJW2
TkWwrxyzK8QcQ8FtxxqfUrZUSECs5gIWrU9QL2C7j564hx+QTMVdc8+63jdM5ovo
dD4ViOMTmlmONdxj2Uazv1MB9GcTpsYKrq023A7qRSM87zL8CF9rmOJfQYEuI9LU
+AmncxIQLBZqWfGRQb3GulhPaeTG7qsykKcZaBARoFeeX/bfJgmltB/k/7jngskU
Kd08rHHfhSyIGYmdkLoQfUmQkJ4LBAJY7wSyHRHoAH3m6tBA6Xl2NBUKL6LGlbhX
/BHD0hM0/frxCQQN2hs59rxESKQCaJ/g2/OGSoIuzn/12zrXdRT8lNu51V6aN/23
n7pY6cVh+Nj5lvCdEFybzVPS5dtdpChvzJEuybTDnzALxu5HqEC0McMP0ujMM+Bn
LITaG87mcW7GZPHwaSp7WlY2gWPUt01HUg/NO5OP6R3BtOff4YaI2gR7TzJTGWJf
/5zSlLhnVCmMaBNpgn9Qc9ca8oO1pfMqS69ozbYK8nmiqJJTWYDwSMtY85vG06yr
mQbalRR3XBdIXSRVlxSZxnJpdlHFylP7pr9QOqaWy2izRrzb0ZUi4w5eC89l5bG0
iZPQbjRufudRvgIpTWXM/09Q42pzmo0t0Ehh0bqFrDVaQ0Ja+U8UNDHkyit7WafA
HzyJBH4ybSnmtrw+Ulb3kgDlMSTguetrdmtBqPT0fJb0m/NboLri9mMMyZeibAWr
djYHhGgmRThTalOMpetgleIZGb968R15YjVpoKp/RxG2E+5cho917V4bAjnO1khd
xSJM4XBg7egMIwIwrgwcnClvybU/T51QsI9avtNRDyKe5GH0mf1LwzEqK+tL1ZMa
do/Vwwy6/7Ibx0hIXJQkA6ZCmAzN5De9rxvjbxKMJMuXNnhgmtAsmUVdfN96zhh2
USl3cEzkM9Gy+F1K2AFUEnrvoZD/6jof9svYiEkhvSZyN7ZmQ012djU7Y+AdRHPk
cABova3SaCwCZcks8+Tf0lN9hqCuaC6DfW6avfs5FcQrI7DsLMNeKTzZLh0KEba+
qz7Hwy28LXtMjNWToJdMM+Azf+kvKY/GDkVZs82lzSNb+YcVHLSBp7EzPXyZAdWe
o2fwkjkBXwikRctbzrx1C2ryepb77eEXWVbV+qawA62JpyEJCB401DRubzVEkCkf
swJC+KANE02/kROPuefAwlg29HVm7uvHkfWvmVTQWbfgq1uI4AcZmFKbpugOULrl
9Kn7LAtsU6jN/4GJz4byFG78LtpjNwUXV17AXK6koaWjDCwurUyUWXu79oWMBQ4w
QuBV87AR08D9UlJ1CJKztc+3BWVHcA24aTbUTSgNTl4OUCOohZw9WNTH38ENYLiQ
WtQoLx3vjR/UckhPsSPprzR58jwjWRBbrzfboTNk011xfXr5gN+oRmx9oovH10hA
HvZsSrYYHQPuT7EmvjmdoX2lZsQKx2CoQDdx6BOYtFxCiIELcjW0NiIZtYopM24C
S6IKW4161frkPutXGhmDaz1o7W9VccywkI/7FafUIFfxGvBKlr5JL+fa+7Y6vLBa
zH98ekKDKaBgFvmKhtTSE0oVUjchDaXahA9ebPnhfNh4FoX3qGh0CbnIYQyi0h8k
zbipaFmhITPAfnpGBd0qs3HCsHBcYFQYQ5YcJRuZDuHGfy8m5AZqNxGNwV61FaOd
fywwvDlRBRQTbxAb5WSSQZq7AVNwp5YmOLmYZMpsLZ2GDflPOz62pRycpDst8nqT
C+K8GnIOwq+9lm8idFiXnwR9YIzg1zt+Urt6AjxTL4np0AQgcs/Zu+cu7pi57CWl
QCHniQTxCKRSyN6oXaiNgtoku6ioKcOrhLlEIfzJ1Aywky1HO2IhdvPKHhDkc/5W
Gkw51KUBlYC+wQriGG5k9Mi9oD5PUvTdlbMlCMmrpGTg4m19i+hPKVZgJVzMjV0i
0HDZcgx0/jnK+9nsufOtxU7gO+bLfLul7o3mGGa6q/Jw8W06Gb0q7dkI43olqJPA
fOp4wkylCyP3g8m/rqCQN4tJjxoC474QU4slRg6qAeGhRZChqqwo1JV+D6DjYDxF
I32wgL9CD1zHgDfxVffxYa/hx1jkErWYF7B417l67C51lZNL9JHU6FHftXkFhiq0
E8FX5icOCbmP1C0Np97N14DqMLfOpB41YeHIijbEnPoq4zF5dgFpSrQyRNHXHtUs
3ZhqqrwGoHrabvNdzYEzi7wwFmPJu5v8cB73QLm4DhPj+5jlTKCP1OT81pTbm8tG
LquSZO0KfEKPjGflo3EkrP6mVHsT0MAtLyxi6H3RTFI7/1sVTIWk90YDj0ooC3CA
iu4sfWIdSamc68F0JQtq3SRbhT1fq2aushzMPmqrWDtMrWRN51Rao846hP6PgacM
st+qyoA1fIV4ZthhhdW76ZI2m+1RisUSbAnbRu2tppPkWsO+eeSl4SDJ2p09sCTl
KzACeOF8mqjvnCFN/D029+KiUTAfErc6PCHI+eek+nyKOiEmTbQ73NT/FMVgB37p
Oo46TUPYNn9mmF6aeDhNOmPJ07SoBzoVYrE+hdunkqlhEEF4s8ryqZhHZ0DaTrDF
JthOcUbWQGIK5QqpYnmMSGnw3QM42pIZMZpxNW36TDVU6rDM1KctQoxAn95/p9Jj
MsHJU78x7cZI8NoiGBpcFmDw2EaEU5J7uAfF4dfYpELMv40NL3Jcmwq1O1TeinwP
985+KFpTg3Kna2siQ4NhAm4qDUu4Koi411o/Xr2KBoG4B7z1akh6oRZnECwKN+nJ
dDGkJ/y33u9k7k7WnKGR0QkJBuADzdsUfzIdfvh3f9cOIzQ1XUUxcpvhTsGIYWe4
NehCT8jwBFAAOURLf7qg1GpQy3P3G66vK3nymdIe0AccgPSR5KWPgNN9eeq4ij5Q
e1Kdz7v3xLNS7L565yKGvTEM0iC557w/mtbhjqX/yWeSgcjyuxxUKrET1qKXs5qP
i/EmhvSlwzbCnTNTo+cNO7Q6tSd4RWPkJXIO74q2r+p6Dhy1R7CgLVVz2vikJjai
U8amx5m7i4ZXceM6Ay+0EtxL1EimDx8m5cu20ItBzVJNfeNzaWub+ILiM4tESxR9
erR/x8wlu4W6QGj9NoYENblWNaw6dgGpMXnxWa8UDItThEMolOkIEv18m7D8hriK
/Z3tfdDYquKKoaprT4Xq7MXH5v3nOHUglblrHZpG7Z7KaVoCLuXgS3Ox8YN759Vf
qPRipPVuSHku68J7o1Qj5LW2A8l6MKVK5f3fV2RHmawNrKKdfrKpmTvw4h7dfiAy
MxAeLQ4A1hPko1YwMHu89NN2Vsb0/BOwHCwNQzgg17lN+X6qfEEJGm8Jt8uXOFbu
Tn1Ikge8aFW2yy+x7QizPLla7znhaRbSMeqBiZ3tztmX3XqR0ByMC4+LJaTpkkVh
99AftwEZEuVigY//sgw/MTBA92XgPffxCyuf6Zn57vbyOXHtq559JcCqDcB6QO56
CrUSwiAdnMvpan9ljd8NmtrCcFWwDEfOYNN+hmw4JmGzpjW1xlcME/MKH3KD0+OO
WT02uwYHxb5u8ak6PEKddUqjsPdzxSBeHdvRwfDYC3XjVhZw2vo2Txby8Q/Qy2nd
sWdts5lkVUhTx+FEmBOgTtbR9ZJDxVdyTwgoKG55jTxe/Vik9gxTvqtv7N3nZAUW
DyVGLBsMwskgJ4ixweM/DQzUjJGFeP5c0qIK/D/niX7bbJvZBQMXKY5QupIwMTWU
cFOQZ6WvMY/8O/pca0BO+i6acgUmFcne97kOXQXTPOmuBUmAYxhL4U6BPVM3J7dt
gwl9hmXjcddzLwhMlnp9AYBT4FvaWZlOZFYzuYnvZ9GXr+Hum7SqjNiZYAjJ8aMf
fOeEH/yfnk019Livp4/xADIrDAokWmvtFQzzLSP6DrmDVHce/dvqbWX4Ttub3PH/
IEickzMoVe/qS81k4XCuk9Qm5UTKMXZeiTL54+EzpVCOQoOySQdeK34vhkdF5B13
geD+ltrIKohmPSiLi4p/DKaMtaP5zeep3DiQVCzml8UpR39PNP00360I9yITcAJ9
HCiOfPnYWbURhDuQvvcpFVDL4Ig1c7Rujn+pwleGFPe/U4gi2YvR4wpff9BfpG6Y
t/Xf8/dAQneA8yvEtzpFqK8uMaaurVqa4JeIQnxPO40oPto7mWeRfi2YkavJgbmF
thqBuDXHWiIFBFWUCChaBRGGa5s3dO3ayI4BjSDno5Wbfssyl91hQ1i9V2aapztv
KQseYgdXN9sbtIpJIVkQVepiR3C871PRoN20e+BFIvvGDW4635cLwyX6VCtbh1lk
erbCEJ2hwv6Ze9Z4WrNWHtgVV9P3yI292QWGVFNDZcHCgFlt0QCLTW7yixJY5Rvh
HTKqaqw7LDuq1ToquPBNcv2ZPypCpDJkzD0kjt+lVwKLa82dbVWLlMSWgOKbXh74
oD3pnNRaXL74wSnDN4CRrpR/8tftwABobNhmuFo/NEIhBKCR1PQVc9KJ0It3E0NY
UTSWgGrZsZOxTY7qrYBB+KF5wfoNtzZ56gkpEN4YFHXo2E4lCPNCl9e7nWTFLv7h
FgUOsa7m9Jk57VoSVg1o69yqDqy15XUe7FWngLBsEcWAn7ceO0GllpyueBNdd2ej
HOCUEOUnH5wjsGMKyzxv27Z35rtnZetYb3ZKtBkofSxjiq8JkZEowZUw69XbVkSD
DMxTReIW9Tfen1Nig5ECqOZ1fZ8BsYkbm9kOmUoBWOrVVX2YmtP1put6BSe/JuCq
LNuMN9eonGs7Vbr191eUVKoKcrrwfC1FsAcswgGP5VCKOWB0CGkGncNG+yZHRjZD
ReVn0Pscnp2BlTD+7uoCC57xsM2whiae5NSTP8kJwxWLC1N3b6L7KkEyOSy78VTd
qtCd8tFE/5TOjIGsge8FcqGepCz1jl2sf8pmXkkucxCGe2QVX3X4khbmgpnYcu2t
t/UVp7trkI/4YaamhcMO+RXf9sSl0wGE4rp3LaDWyelVD1rPge3lczGVuwlL35ov
a3wgifHpCcCHT3H+zZxrkj37RAVL8xsAchdrdQ4I57OsPYBsXPCdsmoaFM1DODLB
nqH7qWmgkMAVehlaPyBLoKPoBEnUMBrbC9tt5hyVLtNumBjAWs4tdNAwN8G8Xdfr
MxkjH1mpFIeMWTCFhhL2txFe2OiX/BU6/I2etIsq3SnZhWLfl9Q88b1C9cG4AKef
ns33K3jJTzayks3/qQCDv+10WVg3hHxUD0WyZWLspc4KAhBJa1rAUqbiBU5/CuG8
9jgajPk+DW0L/dhKmDEUNosFIJImpOYM3jT6CocWhfn9UWu8V3IJTcUK+UtCc0lo
g2cApmCaVzF4zZeApMfS7Kj5rThTaMPeQFT3BgxGJ2l0BJaX2Gygxqpgc3ai8ef3
urKM6E8Nkef2Nrl7EeTxq04tWilGFmlsPwVwTrkhvR2pMuBd/AhjlB194pu3zLao
MTwfP4lNXJEsExhtBRQB7xxHLnN/I1oFPyEluHlH90wBz79um9kD5IiLYRaOtREj
/pf/T00cub2DhpflHPv/CitIWKDLXpNM8+kK3EMpliEmTrQ0ygwVJsMa3a7UUo+G
SEprae6Ep8q7zDzpMSrKNV80ZXUj29r+GsXJXw3vPTI28rQMXUFW94YuOhX6sLZm
hshYovsaRr2xQmef2mUNJojQDzbW/Vw645qy9+eV2riuApC1h3qSBkT/QdysRpiR
4rV4Q4jxeGA0qpRkUDErotQKqzYhxQn8fmLeEbEweon3lQenJyDnE4+lHnWL8FyM
yU14UM6EbWZ4sqVZx+Xfcy9xWq/6SzB4Egdy1b9s+sN0P6/5gfQr+9G5BC9QAFot
4iomWGqe+z3qSvCMWVCpz2Zq+KmAaTnb2BIpP0ISxOddTDIzsgNt0sEH/7GQxx3B
V/1nvtBCEZVQ1haZuOwpu49Fx0JH/y+l0YHxd/Fb/whRJX1jP2CtHlMyECK097uk
XqcJaHnOLShNFKkHu0ESLdG3LIjGy9pPubUUi4urj0rlL6FOOWL2kgzzo7L7U8WM
uCgGENfAAeV8dKu2Ym7Dq2FT0RjZLxw1MH3Vq1kMrBmBdWDPF1o4q2m/4XFkkCYY
SS1xnUhnVP3LmdFfFogQUYQTDySCsEKFuqOaAYsmLVNJFsRGtaJzBU9wNSS2O4ta
IiiM4lMV6ACMVvVp7PHuu2SlP3f3Zjf6f5Sn5TnJQ03KO81FCodzMzZkGYqW3jOk
cm97WsyW1fiCMA3L8QqcOG8n43dGpVOVn4LJRNfrDy/h08kVWKplQnBGmkMgeJ5F
Aq+G/12+xkIaVJeRqzVULhb9Zj4xAGr6N6qpQ0ZFlgKIOEyi8jSpbJD6b6YZy/Nx
gx5LCO0ulDLPNFcDPJnZ7eDlapy51d5Jcrf03dr8vZAgIh11AJqk95GbHGFGhE0s
9OgL5G7+a1BkkRFVVQbw6CnxAFjP4jHDDXcuRx9uuS3+jvNFDJV2vOstwwaKFGA2
dzZ6Pj3plsc2oxUtd6Syk9n4A1w838e7W61ZBnWRz820A2+MDMPqbOAfZpBx1NIi
eQRRZbqX9C5teP5pD83BKcN0WB7bPv3ps9Xicj9KF+zYrQS+FPAv2D55jm96hMK1
DQ0kWiB0PhOODCRP7QUUlkPnCP2qCfbw7gEdUzhLimkoab0HVzFxcfvYEj1+Ki1i
eBWq39I/XnYuX3hYoSdzy0u+xrwcjrf9I0pVvw6P1smr/WPLBdFxVygoeVOcZJrJ
y0epuBrMat33CG9s9f+DlbhERthmhA41n+YgUOULqgMtyRKpCuHcWMqPZJ+hha2l
nhbBF5/7MFGo4PXLHszCwig+7+3TQxcylfILNzR0tc3vNI3PHVoSseCPN1ZqxJ7u
5bjcC12VS5Ne1m8SWl96s0YeSf+b6rHVxcvK/kH/PsAqMZTZ0zJThx60x4Kgr0ji
EG3QqnVxhHSZbAgwLsdImEh0cwfpr8myio5FtF9BJ0TRQT8Xo4at5YFfF1CvG0I3
ZmSL0rVBlewxoS/dmfpCDG6ICenSy7FeG2+E1ON22fk6IqQoaQcttb5y0hoHdcB5
Z/CWwStK5qu/idUDiT6mQpmXEsK330wcD/IFw/Ks80iN/mjw5FCmY5O1ouaJVkZD
SNUaDlFDrBS4DDLq0KGXdDj6wsfPlWWlS04HyHYD9xkFUs8YKxgbKPxdEE55g69U
l5Xb0EtxirhB2hnUO9g+x0zGS1NZigYoe2J3iTjqFqKEnOxsmKXbWJxohl3ZjfHh
YWWeF907S6A3boIONoeUmQA8eH8qkC7/BL5UZjZRI3l7s6ggJBl/V0OCP3NJvSEm
MJIbQiVaiAxVlmkJDucCMJj/48q3wKmRnczjUNakIgqIA1p8ASz0kuzJ+YQPAsvR
4ue9YHprqbz6u0nBWXk4P2qBsD28B4xK9/919gxpCGcB0Da/sxrhVm76rWZUo6Ao
vi+0KyB5ptu7OXyLY4MU+lqaZzw1PNIDEnVkYUl/xExkrLIV/5adAP53tuL5876c
SoduO7fupqeSF3xq/yFXHuqBQhvQI2RckOpBUmpF3kASeAOmnMR1f/QuXtK19Ree
K3d6OaQ3rQKbJ0ZyUoPDkWKA4gSdUewHaUWoFx4a1SLpYRa+6049ZLY38OTe7vk0
HmEC2Y2KdIdhrpMezyQHDZizK8sajVMeLhvHDwQ7dqefH+gs8oKH0BhJ/qGl2ftV
PFTsAzr1Cd/aAdYFVdzTb1DT5zr/hmgEFL6ZRIFW1AdrdiROrZ8pp2vEAUogSpPT
qWO6nfl3v5O1KhFTbc1oEfCPI1j2ai0odwKvuginQySVufqAUZhDU6IWdVD92Gw9
GpGcRmfFObbWewHSzxgM42y7QowPrwU6TTJwoKJm5TuZrQGEm0107X8Qgv0+YZDp
VdzoJK77qOseFzt4Z/2VCFRpbDOKFIS2sc/tZ5xtipWg0MYtqKkeJiSnRxGXjSMz
dXO5YBP0zOh+5bMeqHlBdzxykPCUrCcgmpspwS22vwh7ubm5O98szGnsEfXXTC0I
3SCOhxEkq1xxujA53P00qEGs/Bg/aDlSeAUhmGpw+7GhxZiH1PSMZ+hxrd5qB7WL
pn/vWSaqoYf8faOhwP3tLpYaNS7SnCkV1UBUv894FcUuMkbmOno2NQON+jbyFSyg
H+kHlCFYE1oaFaJTDUSOR8uSfhT5BOUrkaAU8v+5Xsx+eRJGkqMsppC01N3ORiOt
8v1sn2LvU5BgtwiMvrEFtguQSRcZDN3KgLwC6IFxHE0lvF9KLbcRUEwh1ICdUFFy
R9wEq8dqUoQjvJmHLAPknXhesch1oRSQHGL2yBmM6ppgB0dlQOyMjkqWBDY+SYRu
UMmb2+bc59votLpYhC3ouRG7YMiX8AwtUUUt2fyce/882wzdhkdpkI0CYvqxkQwI
cjLWUH4HxxBWc/PfokbaWU3sD5je9a2kp/rZ4vDC/wbEsaI8Oomrv1bP6j2bqSP+
v/yNLwmueZ4NMKFe2BBwM5HIbJO04YgRmgIoOar2YLZmMS8UAh7NWAP8MvAn3Wp8
TIQezpaLrrjE+RpqGiwnej9ictDgN6wNwoCMiD/j1FKaUEYqoAUu5/Pc0coZEWJ2
bzUSkqjKiJZiZw07zfDDJ7up7Ey2XOdYuuGuMGYUTAksfUUAo+RrUBbhYmhs6Hly
7C+h8UW8bbRmNVPhsTm0wsKFfLLPgp0I7b/lhgwHw3HJ0nPgJfsJGZksmd9omtHX
sngPoqvklAig/EKWT7ppgmKLanuxIHsx39gFV0DQ3IXGbKagL1IdnOLAR/wixjdk
tToWX+YDTHschryxiQetCr9nbSmV1+9qTCgacFJhXQVhsBQK7Eg598tNr90S8Q9a
woEF01wE1gkvvNh6aa3bIfD9yqpXaIpPosJygi2HW7BBoEURQkgiQsDg4C/clILY
qeGd2E4ztkmjzp09I4Bu2ebOCj/Kso3jF+Me3iREn2VAmW+Xaj/ZXvQ8t74zWVen
aIla+wlGnIRsngNvfE7/2Q4G/3C70RttBXbbhJdhgChuuMvr+blHs8DY2TQ4Z87w
z6UnN0cI6VIIwvipjtm7zlSZdXbWXN12vfkA3DYwXu6pmMhFc2WCfgoUC5Q8eyPa
2WGhT65W6x9Gd3KCq3V/s4g3ML5vjbPWnkKpqUWZKiMMD+jQPAYZd2ZuJRqgg2+S
i1J3QJM9/3B+M1pdNFzqXEAXQbYyGyF7Pn4VOb+x5tc8PGyySwP6uMaJfV3CooCa
xr7BDozcRf6ZLSjqR0Sh9cNe0s9Gr8BAz7FaGPIboigLbiToxGApox+9x7akHLMt
CMVlbG1cu6c3DNlfabzuFOoUEOrdk8friug2so5QiPjAqcTROPl0VFyvEKOr7E//
1R8DMDGnQC9kcOmjbDH0rkp6+MBlkUMyevBlog+FFZETXvjEyO/NxMbhOY4yKGXq
UhSXHruIm/gV+MV/Mv1fksG1X9kD6xITV1/cZztOA1DYoxvn3w1RGP5UeWHb8yCl
YSj+TSyJyRg3VjFFYkJLAneWQhW6UuWCf9rdlQqEKFLUFMSUqwNZILy2JDoWfB2q
roJQMhWUNBAU85lo8+fk7DQIKblKWtddn523SZeXgU/NlU7WLNRqdA6qdFbOvwtu
1qDz5u8ocQAjq30Ab0W9y1RjPU6DA8eVNbGqRtYC4k/huxnqZTSgXG4Y/Lf5yrLN
VptYw8XabS/5HGXOIAbutGuzDV24ufZ2KWAGqc0LCxXNX2Okk7dZfy5O7Nj17Wjo
iIAMTViMsb6jZhg9hBR/tfacFfNbl+97Yoi0iy5rn857IYPKR8pyrkXd1gzd0QGM
hJD5Siy7J1uhxuI6NtubnnmZJ5WleW2IHGbQv1qB+1NcK6BuYUsHrR1SzF5q/Jdu
isZUmle6BE2ymIsAt4BlG2xnuuCRyoWFpaAbjX4ZRJ8+JJs9ndJHLS/qk8nv3GCN
Hd78SP+DowfKdnrx83eqlKwxXL3Uw1/g7tOYEWQr1KE7Co1J/d+7e6y/GmdgsY6Z
2BQYmhr1T0bq7W3CI//LBo36ZyTPVa5iKQ+iXg1GtDn1RynHdkpG4KsNJ8rKnEB6
otIsoFFz4ZSv+mqtTxSM5vHQZiSS4CbkT0ozUSdpMg1R6mNLY3F7mChzFCQk9DND
tsZ+FXRDoc3cNoSWvjqnUMh0iLGnjAlobXvv6aNPDnu2KWQZQtjSTpLwWzAgMuph
uyeDvmnBc3tCIzH9sDb8hf/sfns9utvyRSVZ4mJh93wu7dOZa0TXAc0gfn56VUTT
4SKKflmj225lTc9ICQLOicJdnMlPmESz8vYYoQTUjUDlIDlGF0ljZnAio00meFMq
8C3GTCtXGzrwXYQytzmLZzKoeUGNcOt1pDPXa1Ri5bVIRgET/z41s25quxcgnBxR
51laZsJu6AWFGk7ojlBU5QDET3/AyWojjCYUkgvvM48h6f9rethbA3zeelrrFY7L
7LPYHInqbpm+5rQYdQKMtCVJtjT0fb3vf2nyVXzEhC6mM/rtZVsdFXXdEKqIGBjD
DEaHQ9Amm3aFdwu3/H3sf0H8hB76tWVS3I2P22uSY2YGCKuyKtwPEapHjXN9PIfW
62DiR2Xlq18qy/D7BllPxG7sx4tQR2EdGuguqjb7/LxH6r/4Sgr7o9oHoonqexjT
3FQ1RnkWw0hN1NKbqbyzodTUNxYRe3KdGrcmMZ0X5BERWDeQ1Ao2jyb/kmds/v9e
FymRyRrl+gCaRBqy36O9Y1B4b1iI4xJB544ea1iCXoLzU8b6N2rAqea5e9CmRY3C
BwQGpYySAh8VNpp+l7HtYDi36qS0kzbOa9JWDjCnQBAz4/JmtGmjOJGYZYU34RMX
AqHIacr6krKfiBVi5uJPR1+itNnFxgGvT+SI+6VgD3c34WjHj4OoWhVkjEfi8BqQ
vF/MCI6Xsdd986KqoV9WQV/hCFulLSeKbGAK7gdU9wfE/xOCjq5FP93rzTjEEMm/
dYSglT7wqVwcrp7y8Vdw+YBT8GmSZCPSahOXMUVUkPqIALJ+/gfrDCC89RXfQjSL
6MhiJVcPJK4EedzZit0F91kef+V1nclUyEs7gCnV4EJb2AAlcLqvc6e0uNRjwsAB
35k1/5vbhGBy24PZb71Jk5A2Bedrr0bzmFOyks5+D5mn1P1Ia6dYDeHzw/ctehrT
Uqm3rTfTkF2JqI0ilK5dlP+H2nduHzrhnPZFfFnBn+q9xRTcTG7Nlg71Yvr9gnsz
HKeA25NzXMENrCXtm8Q9it6od+XBpOEN3a+QFb/JIi8TXh1/9tqV9ToEmHTlnnFH
DjoPXhcZhxZ07Mk+dW8HoFsWcZctoh+YA1SS0Yk43hrMQ5zRNmz3rV+yUYHyipjM
qDJu2TL6l2b42J5+0JRCiYFg78sA8hdkOKVEAh6wGIqzQdKYqG5Pg7Ha0jknHjeF
3lyqvClX+dKFvQyUJdvq3On/wd9S3nAes+fuK3fr/oFzsf2o4hDGJtREG7QWlxcQ
9QmIc9U3xY8fwjQQ6cKfGhnIBncL4zd+ffFWKhyDRk5OdtuexF6NtbFidFoT4N1G
Ca06M7BFMQdmqd6vb7J8oMnDM/Tg7K3W7SXhbbsQoJuixTb1fGMcB2aVtslU5q0x
TTybsStanppXRlQWqd7K2y81+zWlDA6HNNMOOoI59+9bN+5ELWbGUZIiT18/Nu5i
1kK5CHUO7N5dxVdKJP5fXkSoXU2CPynSE0aLPwpzJp4pN2vd+NOKU0gWk+3YiYSJ
rjHeLXzbzw9kuXpCEodmqmpmKM3D2YHGWnqIDGlAlLCvhWoHZYX6ArD9Qc9qvafC
bP1FpSCLZgS7NbOwzK/sIfmhnRIh6Mh174RVvga7bAsCr4ivjKjlLQbOP1D/ATST
l0VTQV8L6SkS/X3L+uO6Kiwi5noblb6iQvseui3zGLgoMD/IeQWW/AxAPYh2lYlE
CVv5tOpgW0p+tVfZwiwjMHGbDL9FgZCXA0a7uIfH2X/xP/rizMoHhhE1B5cIjb1u
dG3uFCn978FBgxUtcomdWhEGJVcHY2I/uAWhvnCBECSi2JNVZoi9yk04yvn1X7E3
i2qoma6AQd0LFTHLv09BgSy7CDV4p8yBVY2eC4b+z9VjHU/1HkUmlLhpOERFi7LJ
0I3qgb/wkIIMY7GP0pSRhcGRfT8GHO9ZwEW83ZWMZanYP06X9IAhV+4u+HRviGMs
aVWGSVJmiQiGUUMimUoR23j66q4W6qfNPBMAUY5waqGEJL3ck9G1Qm3VYHkcmxqo
r3MSwjCqTXQ+A2sIHCbvZQ/L95lgApeGtaUpBRvtP+O+aUGfskbqDa9JOjmjcsWR
UjEzdHCy5M4O7tmlkGKDv2nIwBzq6Ezzz+tsX1FQsq6hX4SSBKRkfj4CMFEYEBpU
xUu7tSYRGmf9MSUTAj/Y8j6dMo2EYgkG5i4UmejgkfaKM/wVESn8g1N16409qHEm
I2k42VmFitOutPDxYzrXzmwDbljZVm3+0/GKvaFzoA86+KbgD0ebu4L6GrPnu9hA
ES3l77H8Ea/IjqNW93aBn7EP0NHGD2yMK2a0LruEsBuif3jOdl5Xgu3UQ/T/7zvJ
3Q6qsaQavHKn4Jyu30eugVx1Go+CvgNSxhbUOAv1bVctXSAQ/pZqMuRD3cj5/Ler
xDz2LO+X8zRWrfF8RVMuqgc6oYFr9b1O6th80+kZ4Jm09zcMlrSy03vg5bR6TWe/
61qdrLSoxiWQh2nkMTLrQPFs666AD6fGs5LzDvu6mDf7VYI6wqAgEIPPX7lwFc+7
5lsk9/jWlCcLbYcPzkuc8AZJa0okF29/wn7qoqiv7+Hoz+g/G1f6uC/5SC43Ki5o
VS9krOaYhmb1X3hZeAhLckfD3cDYUtXwuHYwpQzG3GyHZCMWMOS1y4q+FIlX+6y9
763kfZBrMfSPMK/S8t5mvBEBRpwa1hLI+7jl8uIoMOaePBZcvZqVmSAOvAV1KEHd
F+TkJ07h/zp1EC1AsRFHE+lP6ppB/6GTClRusK0DN52sC7vDEpATiNnSGOilKWRY
9gYqIbPeQHct3BJVmCibG+4y0Y+2KbqQjCg7hT7+bCdfVZ8nmJg1Gcz24z4Sw+pv
IoLyV3RNe1HorkUg609xWTsEJEWNCF/q9jgy5Xn/5H33vinddqCpJeYMQ6hZVKlH
cV+/PIVppCTRv1XKGWogzbbn6uAObdaq38aPfta36zMh5tLxH+vtX6JgLnvTHE9L
vCc0D12RgjUhQq37QpDVXTj/CXBx1AsSqPHSJ01HY1yzjZh3AWK2JjqCmufrvtT7
f3yL/wn7ip4XfyVowVVxTC6+BXCc8hrdq5FMUAVvLeGAUO/isPfeLxqO2gnp55cV
vBHyhuqRrVcFhQAqa/jykL1ScIxBzseIRxLhU0TcFJlliM8QrSDTgA2ISE1KD6eu
vOUZWisAjNSNiE6hixn1BPe4irNfnIGJOAKgHGvPqFcVLN+eaoOHbPxfcIz4A7hI
/TcvwA32/vZVOYfWxvZUTaAytwyRk4bElKMpLhHI7OXJCjkK9SJxlna30QXMU/Yh
HPk4Bl4swbFPSS9jyAK0x8rsOQuxB66XXLe5DS49WAN9AOiCqbwDgnfBVlhN6vyF
opHEt7+LAkJMa7B0nO9k/5W6vwQTILwd7LP6wyWYQibXumAf4A3dmAp+7WBMJyc1
innxYi6kGYxajWmreu6gXj+BUaJbFgQEGQp4keBd7kvJAx5yK7VjcTjxqTE/7Zn/
/KP7ScC+YYa9rAWkp0Ms8ulOa1atoTjnLpM5Cfj+Y25KWGVzFjXvcWrTZjM9a9Rs
HutpFYZzEthgEM8D2Gn7kRGzYGlMnYrKujf/fusGFvB7ZT9dM2IxfO9sq9HOzkEA
crORdg67cpSaXfVNAce40YL9MAwW390uyC5Pcm+cGBdeDedTM5aFDlAyedMp5RsR
FuW7sIM89IoxbCTzn/WZvvDuYkHnRJSdozJLrW4oaLUOwwzdStLCIObm5Ln+X5ZV
eCGXez66SDt8MV9wPr081Yhr9hFIiiWZ7VN04SSa1F8UO4vvrxBqs8a/1SmOWVin
7BFwl1YpGjomSsyIioJa0Gw88n8rIznS3+N4yBqbbirNTXlQrsZiXswNkeKABLbP
EZySpvD88e7yQlc3OtONvippiBWv2WemmnN383tAl0Jo3CidperONDCRvMr9AdKM
PfxV0UbQQyJaycdMHBJgE9Zj1H4tNRv63PoyK1rYRJURV/Yobw7M0h/Cx4S4pX5l
EERHiBGbg3NZ3ffg5nEN7hRNPCVJjggRbvg1yZ4lr/Hy2XSlGtDHnlJ4Qfj2LmxV
WOlBEZTG/ky1ovvloOysVQnEvueCFlYMzS3VlxGOiAuXf+YzYYKKvUe9bRAIlclc
8RSr+FybWlQUKfMFhTqSNnjPCXKoeVYiQ3NZEVKjWBvexCbC2lafxD4SlpmLtNE/
TadXNJNeEMSpc133LrkoWN61s5wD3oFVGaIvMl6qqErXiv8VuITi/eX4PMm1H+lH
5JXgEb8mxtbOuG1A9R08u2liFEQgtX1wLq+Kfj5F4LdNqB91QYYBX50kaS8iOICI
c4foOGyLJJzFZe2ffStDJLl8UbJEYW2V5FUHT1Qf8Yujf0PqW8YngzqZ+nlodSbd
JRb1oY0i4uBYQz/A+6KsMGXJ/4qAaaA6dYXw7Z4PKySRyxY8t+jfUqJQ0pYENdnG
CnihrzUzMNdOOfzf7Gn7dFDE9cE9bfJAiyvJ8JPEAbsxq3bseZYpvbBRBsPtcHKg
WMCp/ySB1bYtpvxOtbVzdu9c5iDIUuB+X0Pcxb8aOz90xcI1z1YGDv2bDVCo5Fso
B7R94awhbQ9uHGGO7CAWgnS1oD2k/ujuKfTiOQShrNfor5xpdBHiyGz+X/KcVQBp
Ja7n+nUJQu+NRgqqAy9+SvlunYbDrDMMMhdY+wj8R740gOPYElenqgkv2BMLfZGY
TzBrHCNJDk51VhVvPMEnR9rojOl6qsnJ0VstjeauroWoEuSmO1GbhBqp/uuQgKTp
adYcIkdALTukYoxFwlWhD4vwv+TRzuMVnVYvgntTGikLed1MCp6VyvRp13WBkla4
NlFu14qqw8ynw39uQTesyqVf1Bz4oRGyou/kn5I+4J3DwsRADmgmhaYI50liv7rL
tYP0bMrt5UXgsaBu6mc+8RDC3B5CM1CS0M7wFP8oFZlOJD9axjyb46GRGA8WyMdL
4gwKZQ6pp/QmwpAvAcqOQERIXsDCnGUBMt9XNjXktnLdLBYNajfrkZFvppac+6q8
ZyRq7fhH+TWjvgSzojfnuMVnIVgTImH9AFvkpvm5rblDxJ1l5pREqMOa/Or9dCVS
UaQXL2XkQFeVacIIAJ2F3tLkfxM9awme3XJ1pAD5rowZNl29wx2lXROvkOYnjPaO
bjzdlfME7iJC2pQ3OBof/h69mnNssMt2ymS1XaN+HtDkmltJ005any8oIpgSxEbk
fW8+kafWPHRlVZtcp8ikHlITAaStn++8wOeuRAZFAypoftG5+UnIErTrjio7EnV/
ILWFMvbfy8WSOo4r3ZV+L7vLfCGvOkDNO46I6ArJBk+1O2wh8Oo/nckkqOZ5QtQB
+KueBBRXMV37QF6HIhzpOAM0aqryLbyrAwDu2tQ1x5za1Oqe9b5beuIlJW3kJZ2m
2lDHMuuslETn2yf1H9ZfQ+TQ71l8Bw3YEKeZRUjczfVtW84MOBpo6+xHMjQTPvJv
LWfI73c7eIvWcOecNjHM16tpFaqKagw0z357fJIVxMWHSP11SqwTRP3Wbf8JiMiK
28FoyCqv1d3ak5HQd/FEfXFtcYWlWkUkhwg5tkbwTyrkwa40zoM2u+VOnMh7S/KL
dIwXgArCKzz2DiJwoooHBYUMpJZi9abJ97Fw9EbMPmHqBpi6nBHK2hx6Jr7515PN
yJmgjnzy7gyHvT0AjCH2JKR1jUUPLNx23gX61Qs7gom0MYl1AWX+3+ui4NgXz6h+
B4AQvUHAjWCV3Nafh//hgOy6aRq69ByYLriNyHNG0AcI38cNm9pod+siS+hiNW4D
/59y8bzP1aSSvJ0V8zOUp9PUhqN56jCObda9sW1htlquHYZZF4CwmsLL7VTOuSQW
wdQSgWZEbsXceUyr6b7j6FyjZnQw+9fD1HbEYxqkaOCJVZps9a7G1yCC6PiYAe5e
QOs7bk3RXYSug9/tpPmGjZ6suNfgBcxDI2FrfisGL+WrXI9I6Vqg3t1n6Ovy1lmP
FSh+EC2eVB/8jeY1j/LVZ/QU1c7/sIOMnGxDRlrTJ/kaMg2YCibJxaHhNUJv8cM6
8TU6T6xH3NXHxv2MHoLIeU2R0irr9F+HwHj4lCZ/0X+TE8+11enSlV2YMU9Acua5
X7V4byTCXpqe3cI/T6OyHUEKhowURlq6QZTg29fnaJns63+wCL6DF7/9bh3JIKM0
89GKBHziqyal+Kjl/eaPOvcdbxwP6/Ikt9KkyHaWC0PETJtpetbgx1cT8ktxv1hc
tVMP8EllKLSGagu4GmByJinRIzthjUunitg+wjeSLt8e0Fsv8Iuvocd7YycKxPvR
MPehTxeAdZ1T8s/23A5DiovAU2Mxe2EOsKIkxqgGUpqk4YiQ2j/14TS7PO0abwMC
5Gu8QmfpzzSreyo55fFzurwIqveh6EormclFNtwbisWfg0na0InmdwL6Wvx3TYs2
dp/b0/vf2TlmEvpngUGPxnXFN8vdOyjevhXx0+OFtg6RbmoUpDR2kgM0a2ME+IOw
5lziZM1qgNdt/KEpWEOAbOFwhzzXyI854KhVTbTzx2Ke5UnteIyD9hqhgD9KqAmc
xHhu6Yve2QMZfTijtd6gMsy5LxIMycBBJODo7k0z1q9syffFO7QhB/Hwsjf1tyoR
prNvri9PKwzrkxJXYqI1CW6noR0U4Dt2FNsWqsMgQzTunFWjq0zCVlaYq1Y50XVZ
nglE+hI+Nk2R085TKGnsiM1ZBpCRsGC/+iS4RfIGIBWp6r9JP7sOeW8hPoduJI/C
eUTySzWNT2VWXRbt2HvezO/BY5Q44iXh7JgZXkXOVjl9dm12rrZ70mKBz7LSAuoj
U2oKxJ2Dv/0PpT4VZ6D0DU7A43Cj9f1KjejYJ2lf+UIStbTt69VWl5SAebpEwk0s
OSGPkli4kXwVPIjgE5sCVHJvLT1oPUK8ZiZD4SSqc2OjobukA9/Dtf/aZ0XSGvHX
c1qslDFcsmH+RlYNPYd9004qcFWyfesTIAj4FVyNsOBoE8Dvm0qP9bMzZkq+m5WE
zqkfrwg5xwcWA6poYDrJ32eoF1xsAJw/cEq6SzRlyGCHXD5ULWCEKDZl/S26pvMS
nN8Dx8txUc9X2pzTm6jv6oZzPhLtQm7HNbFuU9D3RpE+Mb7hQQpjBseoJi53/f3m
IaHF7QfiTlbY0bcPYtmGgao2e+rYiZvo5eATTopQXmfMTWvgSDTrMkHnk/z7ffga
atq8Gx6xX79deekuXR/3F5Q9cMI4+9dp96HV8h5d5bpuqUErle2HzDJiKVohY+Mw
qBTYjAhTxIRJxkuF3hZVQVykP4wkstpyeDgJcNM7/MD8EKchvc/xgFBCLjUeC/4t
VkbfqANL9iKCJX2G95lX+BWaO13XV84W5ZLccO1PGN4UjyThj6B8jyo4yV9dokb6
2exq1zoEevaPpkLiNFsTTik/l2UE9V08BXMXuS0Ne4P3qLnsQRPgchyXmFIqcQ0d
JZJX38V9he4vgTGvEqmbGzxMpi4JwA1n7L6lRiRm2E8mMGSKJAyL3F4Kga4DAcMi
LPKMhcFJi3128ftTNAxz0t1KDyOq64yewYBwxCWgqGRkCdlFKiyYB/vqm4EuMjGY
JZ1eKBie8X4Z2bYoWLSAVOaFnzjA6sSDJ9mCvRSTkO/2nYcU+gjvSYZNqAYMxCSZ
/Vzrk2zBJkU9aiixKhVYOZwrNl2R8Uzafv2sG99X+dgEozzK2vB+VS7UUhpXq6v2
tjkmx2BUGrQIwTBdaeSfN3/eg8iMWgcbPsIWgcb8/7HSnVJ9zq5szVnvcW/Mw8GT
ar7e89sjCZawOhKTGnpx9OIdY0SmpZWeh64iiQENCylGAkbU3PYEmzEIWc/b9BtO
4zfFy88QuwlRpP4ocuNVlBOLY4/azkBrZs+b84a1f9zOCQviqH5+ht1pz4ajwdvX
ggJawOX2CuaW945i1iKpCb19mqF/bBbsXOvACoYuAQdEcACxQ35yr573gZ5ElG1h
G5G08dpgayALPDitAX4uhOYEYWa4PvxT6yeRS2ttYDsC/t7v005TEXcDvOmhcSUv
XXcsUQB3WYUcBPWjwFwtIfNxOneXtlNal+CuClfCvuw6Uk5AlBctJDVl+gUZxPJH
pFRm2Pucilbpce0VGybAgymooY7bJTyj87vZu9AdKxk7N2ncoV2RcYJ53dGgc0RB
Oe3WKZTF1nUFfWGrxMzzXQTHZnMz/37/8nMJgYm20DUdzjIgFrS6Dll1kyz1v4bk
ePMMDTb9iSQomzd5MmbbycPNe7n9HlDTzleCV0EAaoo6sdNZlpFyYjj+RSL3M051
vCOnMUeiQd0F0vqJYd0F6UpyTc92O3WxrtVaPpTffwGb/580IZH8c/g4pzlh28MN
LcH0ywku09mKOu9Jct1HxQdMFDjn+Wq9yVsZCxUnuZFzVqMWSLp7vuns8ocdYzva
lD6ZTsEdLMGYgoqNtVdrupN4d2R6gnrqDUOaNCakovAsHPqb5aau2D/ih6FMrhKo
BwnQm8jhU9P0SYkrSgsbC6j9rr2lNfSVOoyOjHGg+QMgkwC5u9ziMJiG7Hnr7MiF
bx/WQoaVfKkR6Uo1+RomIAiTzQAn9vYEfuQyN6kXMyV8KTL99q9FBcxvOQvoWksr
EQLcHCo1fabK3LpQ24WYlPvdUaXtBbHe4+tXB8A+FgCnSrl/6+9fflrN8HMdv6rR
P2ZRtKHWsBqYyjRP4lHjwVu/CqrPKAEtHz4bS9JWnuutLTSOSraHkwqW1is/zQtE
G6CNex8lbHjU1+7z/XpLkGaFrnRYtDOGxhvHxAPmjTEQLDi6/N5bzp1UsVazXeSf
yRR9OdLVDXeLuebQ7dxUPZcdSCpeTHsJUhJQ95g6KKoObnJ0L4dz6zYAL7fqRGh5
G5Dm0EXM8AnrynOSRgtQp25+NhIAB8klry+FkgVYqhZfzs11kIYz4SnKqjkwG2Xf
P2MxS/AmiO2SsYuhmj72Gn9V1HZa/Vb1KUa8ZYfMiyQTw3Wt35P+wKm7o1hNz40I
ugLoHn0kZ2AWFDZOt+srzivPx8hYLEKHAsVpn4iPfe88a+6M06mrniN4A8CGIBOm
xN0HxdM+iwSgZp9IIx5Kpt+64TGrFAuYtD98COMjqav9qjQOvAXE9ZusFarTJ2zu
G4K3tmBsjvf3/+BIAFNSnLrW9JyyhipBAotJKqNBxMHApPqPW8UF2cOOTEwNJ+Kh
LghOijFHp0LF/121JHNWq4Y3GYgYm+CdPe5VvcWhPkrd3o1lxSKAkAcXqh028lu7
EtCkpNOqmPEOpRMv7x9YfNyn1Ap3utiMtpYgqP+ZUvE5CQmHWkkhSdaNx8bRXpj2
9K0YsQGzmfrvmC5wD8o/nwU0CajgkBnbekYdxHGAyCKq/QZEjOctgtR3FKjMG3H9
IQYd/TBAMaAblfKJnlOa+6IcPFcAV/Ks7PoLthUlSGaFi4hbhXE4ejHhFWpJxCDp
Pejb6y7Yn6RWKoqrKI8HGpAt/fLZB+9O+2jFHRYymXXQtNaVC4EOsWQeXltY0OHO
922KDxZ4VyBivTUQNAqdHjgfmdeVwvTCEPGna6NvQ5rstDE0FvxeQ0spCHijXqyo
NWUkaV7osu5/fHMJizmZ5Ck4wb+rl2nM/qE9QfUqZ7ldmyLwQG/+Zup44JcIuPg0
ewh990DAoy9WmBRNM6v2X9RSbuzYsStHATY0tiftnHybHP7AdWz1COEjE9iS9Z7E
JzkIiO2XWE5ROwZ19qPMvomsjJeOK6Qvf/HuLqSzUBbJ85MClgAv91NnrnpwqA72
kg/IxGJuDU/belilwzYqq+O2UjVuf5xej/DC5x3LaZMaygUvjQs/2kLGw0HoxJP0
AbWST9VEjrK8pzW7KGRMZH18cFAPGOlBLr7c37F3QwSxfsssm666VzAREkbLzlPU
CphABbQiFOwHNqte8qkLpSEmbREVd2eSyIzxqKqng32E84tcS6sGGFeyKxPuxMQq
s1IAQCXG9phCRxnX3TBmrh+bB5VvQxYbhoRlrBKsP0+14QHBhysdhMfe7M0Gr04M
Sy4dT33qF/dKF0Gn8vAokpxioGAkrUM4KYVuqQOAOwejHRniIvdQbn36wQc4tMRn
riN9mxS7o/s78+AVuVbAEIC729aXwxNPgU6mwqfsaQYPlBHf5w0jCgMKgZ/5pgph
SG0BOszg5KpQHAOdUaUDXdIgz2Ld+PrJvAV7DThT4ggSCb4u1bIc8YRrhyY0u6nT
PbbYwHevGYfCSPinSSq5i3TVFnhxg38uItE2xTwqFSKa84OvJAEWrA92Pwhm0NdF
6AMKo4h508lkOPFY8AzNnqmhiw7w3vJy8+tLyY4limk1KPmj//SCzB1SOulP8gJW
I1Xf8D3q3GlC+3cxzeko2hZGucC21+L1/Z2Tq/Ygz5bXt+uxXzHC95Cl5ZP+ec9m
GGEfpZd9oJhbqLcM1ubirMkFeeTE8A/vgLg3NsBKmOit6ksL6AGsQ0RC6V7X4ioa
DDIzYYr6F9zwkHBWOx3ynqEyyPuogzCMb5ItGZmZ1bRT+N+4uuX/vtGjOk3RRNNP
bKScmDjLCeeSnCV7N7v/rLDYoofkMfo+hLQq/zoRD3IC2JckDabFDriXECSt22UK
Jh1WU0NXdsCbkZdlBGhxqvlOdfhFxFLkD66bg9WusRKqzOhj9RbQfiEcMv2hnmnc
NNemlq9QwlVJUw6AaEQs85gHYdHi8HGMI+Nyn4LA22qHUJQTwDnFEg/bFnV5oP7s
JvaKGqCDl1p3IpbuTIvz3ruuyKABJb1tOCpypgxpvNjI9TEIgcCbs6W6ePMKUBNk
ogwC+oJirdtU3dTpGeOSJfXOjzFKX8NI0hF/ARCYGEOvDuhsQdkizoQdnnqqXhlI
F4mzh28UE1dBkvExWFEXOYuKK9SN9AGRLbNg1Y8OsSQFdD+C4V9S54Yy0U4UMs41
AyXdn++bVNV555/ZwmoLWC/tJ0ACO7WSEomhKYbPGYno+qPqyjTxjCrGkVXcCD7B
dJnwoP5r3MpG9v8USr+qoBTQak/Jq8GNpOWrld8bmKgHxHeV9Vvyl5HIvqhJRRso
y0t+WWGILWqB3i7zK4XwkqOP0DAqmsTISZp5x2lLIhtwGIENSScJAsJHzai1/MxV
nspwiBazl1gVPhXizyu003Z5eYWp2VejEak5FqZ1dfXPIpGUh6M5wP0NzKA3HDSh
Oqj0LimwiT56yA48ZPKUjp13NkxBM+kxeL0lxNKJYmN6nvzPJRk6mNEkQseHy9Hj
YB9+6yhsmK9ihDJkRtH5YJQPlUg/e8Gwx9o88o00WuX+fAacn09j8eESQd854+oI
OaLbRVQzflMfFKd0MBn1FerECHeS/gQPmyVXxU44wqmVpBEf5PGf89NeulCE3Sxe
ypdPD/4w4PaqNFmE6q+rCoyztIoMfkDRJ8sQkxE6ZHrPZ/+tnSJKtDhaYY28+ykr
IG24yUeDkC4VoTwHx/G3cvoRkcEf+9LNlm4PZ8KZnLYtunjFhFvcZCiLiYZ9kNAm
uUnyJjupJfb9/abHYWadbh8HoqjnKR0UBII0aFnr2S3j6t/C3BkpXPuUtch6AqBE
VOV8PnOp5P5q8x6G9PETDgmhiSvYHEnx9Vx79FeCN5WJIgGWtkjW489x2J/Udi8G
rNEEhG//a9fZGxfwF5889z0WzMWarIVEqE1rBqKu0wUZuMyEerw7c/gWhiaPMbQH
K5TWN9az981pC5K8zMx/Zkfb8mMI48E0RaDh1LxNDraUpqzEbJIMHkwy6cUw3oj5
1RzrlHO/6zZPSN8eRcQNBRiTxxMfhncpvmEyND8N6p1ZYsi8pXjFMPeFgwkRA/zo
e9HHM9OYK2VWlHqR3O7/oGbOON8Rommb3eDsrTxl3hhtiRWjoCuqWIOV0vkfdZXW
FphkYKJAg7j/3tHDlJ/3UlqwF0Fv5FCX01woVAYUZcA8PoXPbBml5VmH/IqsaMdX
zg88BwhkVCwEwZclPFyfSZBzhO4bOE+RadDFtBmF8onMKSD6N1lzkcD1QAn4mOcN
FaGFJQWujOUUFlqX4UKtiHrBPNbgwqW5b7mdPM5AYQz7eSpSfTKUrRZuY4CUWBgP
S0Q+3Dk3UZ58dvpa06fGUdQfBGVLKHSbfp8xbA98q/HI5PVtrahHe8/YVYsnn5wr
TKiala32Z0dZgRRS4nWhLWFO+EliHymmqF2CG24VYy3pSkZ8TWCEIclqDY2QSK8R
w6MjA2znkL8ckv5WnWuQy0kN2YL9xFSunjEqPMquYiuBMEM4ioIebKh6x88GOqEy
WLDRnn+WlDuQSQdlArqY5KO+Tgz37nMVL3UHuumQkrAV2f2NLuq1KFNkwc822X5i
+ooaC4oF3NgPdgxkKZMyYNUG6xsp0MVDKFO9syKqSKhlegqbbLOzBo4M8evblDXC
SextH32fVbLsBsPe8YW2/H4niYKOYospMqZJFotAk0HfUErTwjDgCZw5CylsxVwI
knn/vffSmkcfUpkL50x3H1DUAoVSjari7BWvyGwLaC4G5tewfA+QJMN/7vAUXaAD
rDAGLQ+FqC33v6G0xNABEVfuXg+SwyCVcLPn/ktD15BqX15vWP435QKiunKf2dIH
d6q6y8G31dECdHOpKXqcigg1JYWn856wTA8Cd2u7UYszenanxWoEkTGKDIA7e3MZ
Yy+dqn4Hno6KhyJ7b99a3a2QTGGbEX4uQySuV4kDsH91e5SmaXAAuMO+2PC5Q8c7
Lm3AY9KxTC/yC+jxMLXkomA7K6y0w2WJcvIFy9IxyTcmQJaP7yljKbId0I7wZiLP
Vj5YViAqaT9V0ENc+NpHNp6CjMPp093Qb4MsaRR3bx9bVOU7JM6O5oNQH5W7r/+k
tABBx+EZ5+yw58AldcVoPHKztRqwBviLFQgpNVw29rEeOXpJQpVsNGnE/uuTP81F
7nK21MBRAY/k/FXETfsvivfSxXL0aZ6oxGnQ7di1CSjpqjx/rl7UWXbZE/XM+/lo
5vbLej0aRLTxnBV6fr643etuGu7NMsz3sz1wUH1DSeQjKcUs5AU5+kgJJRHVNJQn
X0jIW3+86ex2T8nFhTI5W07U4rIvALxW5wxTzratKoXCThpBWI1zrJjBhG2iku9T
8LcpUE/S2UXHHpe9pSGSeIkCVOw7bpbafmMOP/EpC6GaWyhvIj2JSqSHVQmT+vKR
AfaYkMRaZugGX/hOvui9gIvrkIM08ltAgYTI4J0FB8Qny7b2p37udk86BI+xAZrc
TM4nBD6lGZ9JG24w8wMRBqUzE4o15cmC4bCggfxeQD5OIF84UJfnQyC4eP96taBq
d7Muiy2VNf1fPe4g6YFB4OCTKOyGsM+KT1ArX4HwsAty3CF/kcqE88vx7sJy0iuK
7570tM35i74eI55MOb5IoaPsY1erGPF30Y9GahRUBi7v5BIuXSMaXJo+bbPyrLdF
zgiiuoRc6BpiUogamiMTx0gCWzJ4OcerKQQ3EY24dn2FmkWw5ycoTOz8pbGxuagW
3ikrZ2zrC1COTKjOXt3bZBnNf2rCkDubH0SbN1935xi+2UCORcriMa2ZeyiJ4m1v
Us21uPIaBtjnpJsXi6uXtPYID+Ljh6D2dX36fgGhrhp+MvMTWE006YUUwnAUak6I
d/WZskD3Pj4o0+zsqPZ4e5l8Xa8k97GJX6zz1Bgeff3DXX0GrI/vDoeBCJxW+BTq
hWDL22PMXEbdQJdqxli8m93n0EtiKbLf+PAQ/tdgvZ6qDAKkJvYx9W6lVfj+84EI
e9u6W+P9F8gk0bwem3xRZ4+7dnz7XaipZt8z0V8qmdQOxGlmNTB6Y0cu0jE/Yt/V
C/ZnE3yDoHG+vtteao8crpX87W69NA2ZS05gUeCoJWwWmMh+EUCe/760PpL9ALDf
mVq2PNeWmTBIDpKzEfJ1zZYxjIPXJp1nxfhjbK0E7kvAMz10Pmlk9rYjwv+Fmcrz
G4OmlkIRYld4I5sIDb9ELqX+x7aSPGviMyiahdmM7SL4jo1Tyy2q+3aYjtPe4K+3
oXUnitt7wQ8y9NbMnk3Nbd2Hm2JIDarK7qCHtJKpVChQkWMOKTB5DwiqObSFYS5A
WBBATT4ixhqiJYkN4mUMmCdr+fThmCCNsXs1N5cLfllkQYqYBZ08vZeQ2kUQlM6C
+428/91pAg8PLtRSm5dCU4bHMZRNxAa5MjoOGAsnJ243jNPP+bqAwu1iOTxMYVQm
z+8WttnZpzoLKFh8vbQXPC+wuodGuCdfwn5zout5nNUn1hmHJm9lx5tMP9Bbgamk
ohZfS/WMp/hrVpeTKvJA00UoafD1NOh+hZj22SrcA2ptSNvR0GOe6HzKLuj0dy6m
kpk+ULCxo/HgCLsHL3juAPpZnNZmNDscTZ2R5NAVZ1LVK6WVj4SVxbokglqf9FOz
jONfB0y4vG/GPca0Y37WfsJ5rS0+sJl+kOx5+27OPBSYPu43AaR4D3jTGVG3vlYl
rIm7wMsvL0Nu4uo7PJqz6cTNVYxvlQuC9eTBGNx0hifBaSzmSWGAmzHUJTKgBZPy
rOinSPIDoJv7vm2fgE0M/E45amrHaBWWg16gPQuP75jfgiHocG3+oP25ZKFBIxRs
rnCPu4LRuw7xdDvfZhXyPlS3PCeUqwBCGe4eBC9P9LO871Slr3N9LUldQGP10ph1
4V0HmxH+WMNkfztsd0ZRusojxZ93NLlsz7XBhqW7opFE57off8QF3UdhbOr2G61G
fecobEIWmOUdZu3mSnTVMdS60Ik9bnhX7fQCoL8A+2InxFHGZE7nvbs8puADmmhJ
ApRzBiCLo7RCcR9fHuM93aJGsepLV1zja55wGaUMIapzSmdpOUrQ2nY7lpxhwDtw
tfSXmcn/4JC5XsCX0eUAi+HoOxLd7hpF+GSCRRy0zqmhNYU+Zm3j/eEbD+ygYxI4
Gg5Y8UCfWspXOKgqYQO8NkujfBL0hlwclZ/S24eDRtrKVKPfKtsJIGiUcSZxMr/J
yuTuhzbYsUBfevFHPqZs1TVcP+wEyefrBN2sx0H0ReGLjXYvxSX6BhHthDhLV8A9
pPYkKN+C9WJUdAPvW8PbEYhTvpi87kVSaMWhjWdIeWkVNs3EVO+595Mn601fHZcb
7VBRFuq4AXOKDXUpeLkk2QHsEKFEiVFqeNBl2Zh3w6mnxWh7Op9tDUh44F9k/C4i
EadC/9xQ9TCZnsQtcEX1QRatJAWHeJhi11//7RBHZwxu20ICIziWZ5RqJ7oUxlMw
m6OU4MIElaA+un48FHS+lkODCTye32PHzPm/Z8DH2Zr03bat9tCVEw6Kj5xxLi+S
nFIXIldkdsjFPGextp6OThaT1+aSOvodT8qGzx+ycLtC5dY5bRwLo6uL4RYekJYp
R0wZiPzYgD4LO6ddrzJ6Tmbv15MOSSlow85eMN0w6nuAOD1mYrCVN0y22TMvAU+I
ZWL7wXwkaETKhrHEi+84Jx0/v3WWHxnJPmDpE3x08wQvv2PIIx5DDtVXqtlyk8GM
DhOLGMuU45DsdPZHBupoBgODBbNcl4iX+n7okLOzr7+ObRAgk2L7op1nZczDy3uJ
TPxCz/UvtUEO4qFLuCI43ufmLCAhevUB06EhzCPzw8WM9IMPU5klpZbw2hzjFl2K
7nrJ9XYdoo9TUAAPtsOCGFyri6eh9Q9v8ZEMbJStP723/DPtvcoAM3Cwgm4YyAry
M/r3UnufOiicZSa4fwRkxKdLa7p5LLUdX1ikx5xrKssxEvklzKktW39bpQTXg3Ys
1Qoy83lE3hjJ5uev8sNDERfdqzfUA1YYCSeLDSQez0EanQxvG6ZQuWi4R1ZdJOZ3
q7uZr4Zb37+qsS9zYmH+6ZGc/u1RXRzxR9OAxV2+PxiO+UgrYwXmOTgBTbE3r1d5
U1alC/fyXc+HyjUGXJBFdwcjZkclAePyof3CUlyE5xY4FqilZMi3htAe79If5exT
UAZ6lxxId/G7Q1E3zR5cSvOJCxr1oTiRsBoa3A6jbqwomIuBci1eOmdA5aSJQRdJ
sTZJA3Mv45qns8aW2Mo97WfpCs09HVPsRo4TpSw32il+sjpbakdUoE0ThnX3vJtN
vV4YeKFBLblONm/EO9fS7CI62MXUjRhxhnSloq8vtktbZkFbwQ4zoHe9dazNESDz
2MuDlrYwCb07WMTd54X5klrq2GWNpWpPpPZb1ijJZ2CdveM3phDKSiSO9bO4W7tY
ISDW/OCQQuCWb2T2qa95mvJE7j04XoxZeK3KJyP+LBQZwBJv/mLqXI/JYbKJY9ev
Us1PH8DZsNlrflmk+VQ1SVGZ5a5ic0IFtr8PF74lSkoy4lR8ATUeDjoqdlbJKydE
w6gJVyqjKUajMgTkoMZZgHrcpIdx3l1FwMrqTTJbxABSIU3gPJ1EINmFna+iZZpo
xXoIjknukgmOIdjk6tAdfCrn73EsfGxZLm5FAHe/9/kISgWZcqluMqf5ZSstQnT0
UvBaui04SvhdylZhoeZPdP0WdhGwN6Vxvn/fOp+eCmqWZEWHzEJN3JsAwGBlZPvt
1rpvzuXhAV2VVMIr511go80B3uFE/ZFaKU1NrJ91Ra7TPDoBeu5Jq7LucZtVmZc7
OyPv+Ssx5AEgWPzj9K2Bfmt2BA3W+dHiZZpZrSN0n46b5BnH7LC1nsVsUywd5Kp1
qx9yfIvYbtquuIO5LE+t2ftszmYd4Fpyj805lVSWvSQDkusFE7wsnOdwfIyjYIqa
QC2nwpi2lGC1tNuSrIgZzjDm1xyF1Ee3yaV6frDf/TAv/aEIMSbwFroOdtkFlziW
/XbjTCBCbc0Gu9vObfVfoltUkQ6mND/cXoAGXEohNe+rBfTJ9ugrTMB8doV6mfrv
/uQBsibGp96rfhwoUMvo7714ZqzMAB76elMyTv/gEVPDhVcCylfx473HEJzr+BLG
kEiJFsYjCkjQsOl3GWyYZRBaCkf+I3LuYLhRHbaO1UMVM/POubfmeeUcd4bmNMut
cS2ouiikEgHpXix2TQsrXt27cKeUT6oKrENxF2z4ih4GXbgI7J1IvxIJCb0rX4cm
jKFTOkQAJLh1r5vnjgWoqGVCs5i9QYdKfqbsSUY+9HV3n9IN+7BzaL6snHRv8EOP
ZSZLcmZRycjZYYJw0Qj2CC52dcnlIMxQx9IkGWbVHRLfqEY5Dr3Aqhg4i9wE9ijU
l4MoRCD/Hw8LF0gunmH9o6ym8WGzSAQiH7ug9V3y+sk7YQkNBQb90kF0QAQm6Gen
u0U0bSuI4fruE/dd3oVDzpaggfWFWL5kpXrCN/D922hlqOKlY6ZmzHXBx64eGO5N
1ltKSY88FUnEef1CAtBUKDdztJSZVud87zouqTN5zdPaS5d9eom+rZaozUpVpo4b
x03A1eUYaITKOOo43sNMe7Hsg58VEUj0yZcldiL8R+wjdROdiGCy0phMY6O+cZov
lRvncb1L3naY3cOW+P1DqAQdeBOpb8rX2/73WF3ieqcZogj8aDwUS3PQ2p/93a25
4rZEkynwMSWURGXf+lVDoHOVRiWJ+6Ut2W9BiS/T3PX+pg+azCMLyzlpVwiIbVpn
xcxi4IFEjRwYA1OX4NBUnY7K7o4t8Zzlpc3MQEaTGGwoPgq+d1BmGHNWk290J9/W
ECCuYspQlivF3HwjO6ghTvm4rF4B2lhsnCbDcOwq55Y1zwcd1Y9xU6pr8TkuPTx5
gqrWu+5XxTbMkWT+oUxBloxI+BQbPHYiJMpLE/tyXJrqs6G9Tv5WuxH8u//DpzKE
Rl6NVI631xQ17SLHLUQ32fJyb4/irvFoGHlc2XwVJjctRf7KAPYDhGqtAbxpZTLo
wVtU0YtmgTtg1vYD4WMwqFf1G15XDLfz+swg9Z/bnhcqci4wMNjDliaRCVDNStr+
jM3M21NexFax76SAEbWgFoInDkjg3poFVuRKZ1iA092fpxXqROcbHZXF/yr38Db0
LRo+Ra8lKJZBxyhm9pZYwUXEzeZhxSjOnbLmVvAswfWwLfeNSb8oOra7GX5ZMs0a
4Hf0q6K/foHohWJc7MEIeMIc2a3ZvzTIFRaEAwneNH98beRDAdymmuO5OapKPTQG
MPI58oZRDSRJSY2XucOLaW2ja60BHsHTwNn9Oj2pr0j6i05lbZgJv3ijYDF3Sto5
Hveh+0oHHfrEovLE/PIcj/+YlgtiY/XLj1nihvcH78hibWeyVAXEWSDflGuMQGIW
OtQ+KWEpiCJ0MWLhiMuy+RcgNYvDFbzyNyeAji8wE40AmHhQJU+HJ/RHznTY0PK3
4GGlr0WgcWDM8c9hzGVx9jNI5Vo58yUDZjtB+PEVEbM61n5irTPr8zc7mgVFyYsO
AoNi/Y+t/8J2C/E4KDIAToTHDIrx19LBu5qYgA8VuNhN7LLGWSl4+GN1jycplGhH
yBXY5jojlZO0M7GeRyX8276yu2InWu4r/rojVpBhgF7mHOFnR9gNspmDXYyWG3Ds
jo5DQe/9QpJzMxg4zI6N1xY2tnw+fN+x761i0/ABKAoEoUgtniHKscjYhBPOk4ch
tA0y7ogsIo4EnLfz8GIYqa7ktrpJxOkU6lrX6345IRuyFyuQ6/PkNmqmSkmXM5wu
p6dlVPnQXhmC9fkz7BVWKAkN2jwOVRxaVwEh1M0yp4dYCVM91F4OxHldtrp7WGRA
s8Edm0wxlF44N1qyhjyvBaF19LBiSA1Rgk4FLYD1upkkotcthDF3g2DBQkTKPm+W
Nt+xJ/9IOP8VLjLWO4n1UkQEacaae0UCA2ez2tmAHzADKhkBtZcDbzw3ik8Z1UbQ
ssZV+htPWYA+H6NFO3lF0Q+SalXDD5tj14R8/N/vUqn3qldlzG3UZnI4A/aLZ1Gc
1CcMt+57uP/6sjcJJoNJ/2rS7HUmpx/pNTDq2mN+dCtNmdcNANJOAMAhjofkCdc1
ivCNr2RzIeKiWgEV8a+Sj6gai9lFbQ0UOvdqGuhzvOyamNObSwtMEY/QZZm6CVR8
Nhsinf8WoqyEztwzLdQkdKB2zu9zNFiZ0U1ite7ZRnJATUsmdLtYMtHP4ia16BK8
fAKqtqULeRGZWcprb/68J/kHsWNAGBN0AcyPKwDsPriiBlHGcDvf6kL0+fCKud4f
u5GPLN4enPLLMs2AdI7gsJGKhMfzw6z9ixGFnU5X3pd7KNPEn9k92LA3M3h7+0gf
GTP2QEeb0TauUcrDp2wrH3hAVMZXvxhNHhvYXJ1bRtsIUAj1BymziqIZ+1TAPiWb
wntxT76FuYyO78Ffc1T6p1b9JpA7j5bnUX8CbMgoxdEuo7m/oSMtz9nuH5G3PXVO
i9/g1XALx7kQiGtXWz5nrsRdtTdbM3usrlONoxIm2SwUXJLJrqHq9HmFHCQ7KZoC
d1NTGe05U4Mc8H/dgO8kiRs46zUcw60HedVR41KbNU4kceXAA3ziX4jeOXkNm8rP
YkEJaqejhsgXZnGGwg3jA5Ewk6+4xdkvRoiyQKWQ7Jr4Xe8NSdcrSVW3R0YssEFj
LPCwdxKlFa78xcFaArp1hGOgA0Yc/LTqplMuJQYSEaDD57C2gHl88W4aE3jrKVqz
5m08woNulGwY2Z0oqIvivA7GHjJoc7+eVhNjbjs4uGXKC97VBhgkbXk39L2/m4jg
8yuXSuHSuVdFtascqrzCPQLWmShB6M5TcvFsINeEcroqYi0RJBMO+oaVza57X0nd
JiLhXkvlKso/Hm/ka9pkYFfP7JoQuBZeIHUneFgQVHcU3loQ7bWYF6vh2bEnQUi8
28iSwztw68UF5GD8mb4PEcT5Bs3xGcrlZ+Qtrz4mqlX5cQg3H/YC3ZBcTp3Gh7UZ
uk/n/D+g4bLSppQS9JPWbbmxAmJDJNFyITyH6HyTwB9NjKTzVdJO3DM4Bo7/AvnD
2HRNev+mcII+/a+yBF99zJFRPonB0e3U0G+iaiP/hZB8Pb6PGvRfhw7yvzpnHAE1
DZd1O20qzzjLK2buIzjJSN6Hc0vVAHRUppPkAYj/1HRboD57ygM885w0UTESR26i
CH3ZV6ixv/Dv+JzWI46Gas7+8B8Ui/vxjML1spohG2tUocLl1LmlPjmpUep6jHTa
HSQsBY/FvPljQ5rYrrh6MxFnB1Gh4q6A/VdM7ufnWO+QIQovG6ii/ePmyuAYBVTp
HsfFIFQnInesoezwVK0Lff5WvnmuKcn/Ks9hqEe34wHDeT7lGdSuJ2wJ1QndAq7z
Yv5PocObsd9IkqmXh//vDl3/Ial8cKxpy9Pfwic01y/SM907+qaL7N/0JSwSlPoR
/gJEhf6iogHfrf1ZjiAgUil+9mWpfeIXqhyg47aVH9tvACMdRamJLsln5xEKbRkL
JWQxqm085Vrx4FgZTDbRPpfg1HRhHFZ2D1eM3WmbPPYzIqnvgSc2EzP9nO/Ndd7B
MEfEgwD95wUVHuhO7g6V7+d32zZUfE7NmgJ2J9enH8Tc7zz5PlDC1eavFMBGzI1R
BwH8SEDg9/C4mBwvZCHm7wc+LpnpYYh2O1UoYa3GX9CYFwqH1j41a9+QtXjkdZXb
fmWuZokpzDXt7IvD0sDUxvV4xuA+6G58bHeVRZyK6xrTSphkISPyB9Fbf6vjs0A2
tGVa70KWEIIJCuMzAgfrl4FjKnBBkyiZ554Qm2Wju8GCZ+qWQYgpBnDlrTNzHD7H
bKn55DHrvlfUsTMbRQM2egdR8gC5XDoC1irmaYm1Ys8hQjV8ShIeVBTqXVVkBx1a
c9DYClbvnmtm1281U0t9XiXUctpr7dR6kR2pn7hMuLX81P/MuJwLIfkn30fZ9EWR
UZ5MJkpMYfr8alHZy7cfOtgZqxn9MYDPgq/9ZBczqUbTVMMgw414whPTPNKPsKuV
pR5uXENr6CVcBL3YmAAuTQOjXLU2tOZbiTMHjBnbQfXmSbQALIDexQBeBis7peob
ambRQliGSgw6zaPMgqkEn9+LBmim3jS0ljHMo4FfqPuEpicfM0tYLes4/Jaco8SO
/qLBiYyz5+mmkkUAa5cc3wUB+pxnn6HVYSlXQwE6XM6LO8xq72THJzTmvrlLPNzb
vsv96ZaiG1Vd+x5kM/2o/uc6z0Jx76/pgksZzGxwLPk7sgOPwXbMiAMNVu9HrRxS
FOrAbQljFosZT5RMpv8Q1ai9ws1xkkH2+9i4j1yklelzjmRMUOb0pjzk2FACFFYY
F/nvFGXTkeXoRLqxBL6Zmk+YTqDlO0G6gy2o6UhyQc/cq90vXfgpT+gVuhIUwrWo
z4JcYk6YXUmoZ7j9l0BK/F03/HNvnhTYDP7TP5VhrUKRo88sTWuizbFj4ZpdlX2x
KCh3Sh7gTY4G0cPCrM4or2Z2UV5PuQmVwX0vlyxTU27Cg2Sl/6NROzMLCIUa4OYX
RT9M82PkzilN+d8D0a3i0Ha2+w4hL5zFSwQ8ONQl1ceLcMseTSCRhuXQOxNSeEwn
w+WiI1bzkIgdLAGXAsq4dASUOTdBe2O7c8xr4y0ixhS2NzWwwEz+5AyNjWsSF3eH
8GtJhwC2Nw1jheIxQMCfqohCWxsxz8gVP4J1kvv+zDU5dua6M5TcJzzpNVhmCi2b
4lcx/Lb2WoqCMzDJnqwenjpVFQrLOJuFPmK0n+N/Jed8isXM8CQe296igtWTlRpI
rAkzUCrYPvI+28sssNW20VRYYv+BTx9XmCWeA0En0OnMH+9dqHEn1SVQ9Vsz5WrO
k5d3p24UuEcktcofFOvj8teO5ettABkuyJCWXrVodEdWHEMEnM6luBvvwmWGPYt6
7ei7V7KyZKGDPCDbOxLRjnPKz+vK4PwYtCifdPwSQ1JrcJDmheKkOon+7WmlYW+S
OhEj7uJ2vyrbwyRBSU2YTYhZFFDjOwMt2vNyN11dfslcFPZ6oqcuwwE177otHkFc
9z3RRCyqphUNM0PhnRQsX6EwrEVyorDo+0MrNliw+gxOWNYEGLVqdoWj7oSXaCNF
EQ49zyrhhoiJevsAbm768oiiKPP8V6h434axsr6vLIQ3zXD11ntvOZdNyKmgW6U/
OLUh/9iPCwV5JHthJ4KJwpL26G50Uh2DDCacfGFXPxnBInbZq5aQrWJhVpeRDQQZ
gWIjAQTMSGHCKBjHEcaW3W/zGjpPrm8fIc+HbCtxb/23mCnJQoE/b3TVC2D7cSQY
gr8u/0E6lqkQoOZu4BmULxaCj7HcqU97FaPGmtcAQK5toi+J1rwYMjDinU8SYcUr
Ak63tL1zh9qOHEiE/btNbfuFoACcIP+myqZLDCMTsmpIpwq3YRSjAvR8zwcNaQDF
XNfsFR6neToV6I8Qfrfrh1jpAZUAjShhaPBmBf/DDMSsdW5I5bg8C1tC2zvpXvdX
jjmsWcLHv04ifNHyig8EbmM52Iq/cyBH7mY9QsNA6pDhc1op+k1hWh0mxxBpvxN7
TkxgBBDlg4T1LlYkKCkf7pZHhqsCxzDH2EP64qx4Hl+jac9wjWGdjm/y86qvty8/
uqdA5BkPWrcbrBAegd+rPidDxpplDtc2KJDS/SIgh1MuQFBWJbOdZUFsHDWaywEb
0dbo7PTOGCLdpPrjmdTKxsxHU6huaC/urNE14VtJFJCWhgpp3nMwK/4jsgtBa3lA
F6+8qQ28dNhYJwhTzfKEJmm52g8sz6PXOSMBVWLokXa84qg3Rw1jvX58KVoVDNFD
XvxPFmjz31oBJxKuZYqe4FMoCEhale7Hi1znU3R50X1DQBP+zH45eHsJl0zbfdJt
8hPOTiAEffAQatwjI29sAGTfNXPWKdrPUfIzC81eWe2LPJo2nWt7EWdhEdJzNS2X
uKN6i69XtTM6mpshHyUSKH1LVg/7+P8GqReXw8j9O4ei1ANyjf2raDpVJrbxKWuO
pCVnatGhlVZSHH2RqD9URYI6F/9jaJdpdaBdwYlBlg3SFCGkzK2YxXkJz7hMyKEL
OrSIwkyFTGUoFl35+1X9uIGYBTszlKk8ame2etXqjPosdf3Pr4c3f4ISUW2G7AnE
HyMRhivGnxeT2u4TU5PInQRbSxPcsQbLYceE0VSnImwJwX22/sg/4EP+odPfiKEQ
XbCzgAjMZakD9kpezWpoQhVPEBQRN5O0ZqDIpmoviTB2djVA4H+LpyYQynlWJcgm
gR6Wn2fFunAoZv85ZGhXvJpF3Osd3k0JITV2WJiGk6QVLNmCh9JU17rZQaBXlGSH
`pragma protect end_protected
