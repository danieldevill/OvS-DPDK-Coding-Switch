// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AhCXolpFVm6tN8pfVTwkDJ1nO9YZuQEWDQ3bKUWc55keYcp8Eh8evNJjWpRg35OB
asFKyCWR8RA4/G+NTSA5SjRlpKH2x0a2rB7z/5oHkTmk7x+in1Lq7blAle55C3uE
peHIXy8luKcZXRw6ns1/b8hr1TOEvNVdA9vGvYp8elI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6944)
2uGsULiJizcnpgtU6IsNpSHVMLdM6aI4jKY20PnLpm1ORmqFo6XGM7GQhll/TG/s
kXCEfNZxFUqx981gVQ5SrQQUQMAJ5YHmsM33EE88sE3b1xj952/hMNQACUkvorQW
1FOtg96qNxVaJ28dBxk2UBLq5G4eepuC2JDv6S3j+z5/+uqmeur6cKIohJM+qohp
uHb25II3Z36hvN5223mF6Qe6IDHvEpoNr39z64RTBCK/KeEfGwXIfLWktaqS3rAk
bX7FDn4YdAIl/MPK/EcZk1bMcaqdgom9cuUA7Q16Doc8WcgV06+q+5vQrz+lDDSF
Spy8zuDgIZ0uijELLhqEcfjW03NFaRnPJvvU74Ry42xmwB9hOiX+UQnzyUx0AhDG
/f8MVVJ4NC7kL4h6KpZSTtRyY9pGDYaOjkEMJo5ZzkT5lRHvJLCBI2p1dffHw55h
MT/2lm5PPCAfk+f6dW3qJa73ySOW0cd+8mfDdaffAHHFEaAW/AA5lGW+FVZIVmZG
19wSw4BVEFSPAUV8OmyZtZpnwLdwvy6DMZA6QRzWR+RtpKXrq8WwR44nt5HC63j6
t+zg6Fq8MquyetPZkTtdAgsQKBDNrq1FodFq8NF4nBDEgXhTfCY1pVN998XQoO03
JAOIC9dFIC/mtxuM2u9lB5b+29Js6GX0oOSI4SCDWCViWtYTlM8F+FGMK/QhAc7E
IHbmVmwup+5WAYyDTEvV2L/d0dGzcCoVvukJIiUwTqaVPFEPAZ5KLPDQ4UyB3/Io
VV0qD4j8P9XrUoT/LUXAdmXh0k5KIoBE6PiIqvdjCrG/nNB1EUn14Yw38TvlH3Mw
+wihyLTyykLXp8uPyJQOgiOWEYcPrvogwOXUcUQv0WJeWAdvxxUz3Dcen5aI84aP
c4F9iddFWPVD8cFHggDjdnyIORjx49wLVByFaoqZRgdVVYcsTKisvn6I5lpUC+dI
uNQaASLGXB1osT90xNYtiqV3r7pes9llmHISGLdr4LXYVgGpYl5uLNPBOWTe6cXu
+NNJMJ3W9XtR43FrpC7DyY0CBcyMGcWKEdx8xEQoBueiDFcKBz+aZEI0/8Crk6w3
4dYgqmSIfyBQtF0blvzqdcVmCNTcmGNUP0lD/OYxfs0XUopRX4GKLkfhF0xalkBd
w+mh4HVnFmL7N8SNEKhoJ6tFF0vUHR5Ld5Ue1ERGJ006qKnA+oMs6EfKwQ+ud8UX
hSfyyThNqcSKc+qdT/tZ38z7ztDKtnJ2EiSDgx4dYqxqz4GaD1583cMqdGnSFpYu
D+iXMOnQ+/ZrneJS1kE8GSJHgsJjdybHJKDyr+QyYHA8ZDHXvL+zGB9jQQ9UB5f+
O+OG/UZOwLwf5cmXMDblJU9creS55W5QWMBuYZSdgbQIIrHTl2tpZTChI36T6G4t
f4OmOxwoJwroUd5/Al6kBP1IxDDHaXzLk/qMSQZ5Kek97GyvnxY0wjaHPQ5at2FV
TEUK7ecJ0+/JV0EEfnJk2B1m4gxoxOKymkWob/aqH0VF8tQmZ2e6Fg5RJCLbdlv9
IYl/x9h1Tbl2OImnOsnk/y/2TXBwINajc5H5HqpbTB7xFijdMl+Vf2xpTe9wqNMl
LsJqUroC149uMiJWF+iG0q0jmHzlSJkHW/ZGQY1G4KLCtQDbcqnyBJ9Gd8k5UNHE
t6kZv/4dvJaGX8zSDzyCp1u5QiPQKMvfKyC49S949zv8kGCQxOlUF4zSKiMZUFOD
2Y+EI774PantkAoevKaaLXqk1xA8E9hDU8Wav/UDYnEK/QUiZzmLhuwI2ascHSfu
1IEHa5EdvRnC6phC+4gw02wykxnKuk4BU4gLQy6xjt2U1jh4qmUdxzRy0EuWTd/Q
IZaS6Oz+u7Wrek7OhSoMLjWD1k53whJGGGoK/1ESY9YPcvItup6ue1sU3RYHBJRX
QQz+KbEPZZ3t9vjSqZ2EeXooJFyHeKHTKOwtFg2TPJGaMABx+u3sh8lQPdiXBp9y
Jnrr+qdEP1iWaXnDB/SJOFXOd1P4vovTZ45/G6P+tePKftRJ6+6e/wgrgcd+xu9w
3rTniMJRTYbEVBJA+33suhJcx+CRH+MublxJmdf0ZHtSfEXC9QU6/u+lUFIHv/az
v5ZSnlcP+yKFvkclhEbYjoWxndIbhsqXvhsuuXXhJk2px9IR0e007GbMHZzD3fzW
ZmEqCXYtHKKxhjDtCv67zgie9oJwJ1HbW3Bha7KKrZk4sMFNXHjD6Y3PhQhDaX9m
LdPtn6s+4ZYPR1jqKlE4iQO2XBMHW3eKAWoaxDPOgfbqkXp/yhOKNLJm9tcjRP0Z
05pwrsVN8WOUntl1BJoRVYya1RM278hQGMFpfu6q9xXXyIawkl0mgHqdQgZJ3dE2
aesCXNugHjfwrtpH836p/fdB8ElYWznh3v/dOPGohrZ4vY7cJseL8CV4JUPdPO2w
GNqMsC09+8+gcU7OXgjjqZA3fPDiJTJKT1aIbQQWmz06Z0iasi1VaSOIgzr97ZMH
jJpuhTIW5PavHahdCNRUc+SPg2DY/rM7iLuOAW1o79UbCrcZ7VskgQkRBfzv0Cl7
qr78/QGGLrymtUJuzXkL6WT6l/EwE6hd48kOLTSykfI8vPrqk+GrNMyIoXauuhiO
GlWLS1jH4h/UvSk2+HNlc8n7BsjJcqPkMCIgc97bcSOdiHe1+MnhryFZxzR9sUBs
sTrwrIMq8JljLHoYe9VD78omD23zvxzzcCY2S1ewfBEtq0FeQyIky0YAHii5iwV2
YsgrdTOsvlTz/5b2+8rTFDyrH1xpByk6O2zYKWXVQTrq9rLCY3fDasvmUJvRkC6G
dI/f+Xycgkvwyq2q9AX+5LlSunb69vW27z5bzLp+4Ztkj8Vspg+VKkSxL+BtQQ01
Ui86IstxUwSdtcJsnOK4bTKCFdeEhkOzPxas0AUZJ4jObwKTlO3o/mTdBZbuVmXc
4C3lgr00sGf75R8WsJ1v1MMgotbBga5OsH2Bjy+9FG9GWL0EUCHWj925WmZ3vLgc
QvTRGiPTsuqTuAXt8gU0FPsTXrSFferqwQSbF7JTgIOh6UaM/6HezXSgAxQRHnW3
h3akjrC3rnd2u9icz+ek5kMnqtzpJjh3Q3pS531wSUPXqfK6oWbKv+mr/ifgwNHd
c8BDxX45mbDXvMdsCjLc+bXJ7n1EATEBS1W9D7xLUVNodHgKW1aA8y63adRHI5Gs
McrJ7UoOuqzDqIlWrRX8teyhX0OKxnx3rX01TdgKoEcaKc673/McF5gHWcolJ8hh
bJ/f09y85AXXdoa4VSAhm6a2zO1FSblyHm8vAd/XKQdmc4CwWPaTHA9zP2DE4Tkq
nEMwPvwDolRsSzMS/WTcrsAlGLnKx8JQKwYVd4P7n5Tub0jxxy8JlQHla0YJdNKg
dMGGEKg13I6v/HMeCQm7UtVxcOjJzTZNdjynEdiK5A0ui+kTKis2I0nvVZieUX/v
xff8irSd7KuFyusTaW43r9fUhFwmPJaBjy5OxIshTEBTKNKdjNiUG76/p3mKWWlw
5YTu0cwh2F/EQBxEpOPOhhyi2dri4t+1ZfKzG6mPPeQCMybqGLkIYjnn5JgFDMEl
q+lSds1e4t91j5Tbg61A+symNGNndEdhMgktl5jFdjAGjBVRTdZt8wPK9X/56jz9
ozCYPUnrFrN371UYx5YD+7ibG3lNzQw11YNkVs3MGKJn21r95Z+/eb0zQTKEK9x1
NbXhnqZczU5lHu3+aU9PlCPnkC6YKBhhgNQZlTD4m+HQgHh9P318ywaxQI5StVJs
JCYeGLdlfkoKlh6VjutTxowre8xjz+VYRptzG4sKglQ5RnFgv5anFCfKHrcpB1Ce
KYbnfzYU6PhpCJ3t2X8ULB5l/CtzhRYtQjn7NzyRGgcANEtJVQlNB17s62fSlLVE
PK/nOuFZC6SBtH5W4TtIAriGUh7zqyyN0MyhKtH/MQ+tNUzMsdTbEMaPw7zlLu8u
m+VJhKSSXWHMvngpzb+avvbEIIwl78SOtQdlDhhs7hYrgqyoBIDE3VzJFroxgu0M
ql1NiJ8px7g5RtB21F/cFt42Ee+uocf7t/02TLy/o8EqpQZYLSgs+C5xvPq33x/w
m8tBy0SFPB1QrMTO51Ev9kXTkbSDbjhXCKgQkon1RlnHOaViuuhY3Oyza2lwfQmf
Df6II1UpLhcLA8xV7RfdmrKTdQWA2m3qABMgTd25XchRqlFkgku781i+jH0jQP3a
yw30lu6vsEQjl85WiUOFsITaaCIV2ZPW3d68ok8lGAohh21nFFZP0XtUViV/ZzLO
jRD7BEs3m8njLzgYmMvuFiZy2P/tmRgrndSDjEupgE7jgaB3qJZZsdAyrrdcwo5h
xZLiFOqSFjctzx47eJhFy5kUz835P/xsR0UjKEBdpvQt9Lg1PIClJwQ0xeP7iWwL
0SqIBgdaNsNTCucBCul5aZnrP7p0JKCymWBkpg2bc65ZrHOBbkyWa4LMMJ/oInqu
fQqG+Akc8sZPTiXG0HX0wxKtOGiSDmyactNviDUpxzjb+5WBD4C4I+O0VghR7w99
etLDtzc3v0s91xVamDBNoG2O8YpAgNeRZvmIIEPj+Sk+yAKmonchwnM6QMuCeye6
Fae9+Ti0dQlKu9uBADLgBt8TYxRIUBuHxKsrf0lP0XrVUhWhmSQWuOQmZZE1c7Ah
Qwge+rOEv/fDE8DDmLqZiH5uUie7pidIhpWa1IpJq1wLyg0HCelKt/0iTvOCpUqn
bQvFB+Okn0KjGOIal+euSiLOzqiAmUxxiKCulryeQ4ko99Dr7IwVtACYTvgWm4gs
yzA3B3jUPcURNnQkX0GUbQ01pA5nDTMoK7Z8V0Z+327Vg1/i4jXRE2Wuvc9S9+8s
/oSlwrY9NC/Qh3rhkYPh6DxGXKGL2HEnJeivObBIup3yhlZTH6cLs0sCTmIS8HW+
IXYicN9SDPQLPYNpq3xCUBYaWO0cjuSxUcRf8VapBFt6sfAyscYgqyRkhf80FG3v
b+hlo3glGE08+z81hMFfD3BgLMeU+gGrGuXguq7pSF3OSu+Kc03UWtUNOTv6wu4h
JLhvNHX2HiyDf+JyxrHAeMxpC1NFXftGmQwoo3R1uuMVPhgh0eHkH5aCpZo6SYXy
487epenA3jvU7RbU/oB3XX92V/04bL6XtTmp3yh40aq3ul8CQhVlE5W7ZLFQupTr
nZU8IikB8sHwoAn6BvsqmjLDXPiuqYXddBYIdItIk8b3Ogdjlim6YncDprOaW1Nz
Fj4Zu83gBXmzrxkm7PPS+uiCqvBR08m9et2/+WohkJL6SoLrF7fYB7qo2linYMRh
eBPmbcIEQ4zAiD/D0BoPrf8h7kyvI8O7b9cYIuWQk8hk+RCH4spOX4n2Ynnb9nsg
9fUsh1d9B1tumXjwodtytWwzXtlaaz9ijpTsV8JMB7qf6ZFZ6B8ZM2kzLXyNwURm
cjiWzydIu/c0ysZllu4i3B11Yqki2Goh+KyypQfV1PFZSJLVlDFeLkkE//tCy6JY
sAV4tR7jpOgnAaKIBX/AA6frhvLp7urXaMIhzcAa0Vbpz52lpndPO28X37QHjQGl
orapcTfnxgPlX0s2Z7/YMWBB8/t4Y02OW+6JAwUX2Ei5EydnHYJRDIGEq+b9NV0R
/zWfatcilWu611ljrFtX2Xo5XzILflXDLPi/vfipm1Mq9+jn5/IOQrOvL264fUUb
Qnua7GHgBDMzCpRQk2vSPgum9E5MEP2MupJ0Cc2AL4UuPh67Na1lumZ75hPZVgIX
sMKzCaAbfsMGMVy+tJtaqD6DIjnqZnLujs7tO4r1uhaZmDjiXq7tNow1yhZB7COM
gPQRD8WoT4DBrGwfNXrkgxUXhr9PzGs3FRQhBhhPALm1R6HE37lM16u1SeZUVcwm
jrgIKxRxuUgwmKpo+qGXEYzhPqWwDQJ2LuihM0BqaU/K4wKFqrrluWeePlg7Ke7A
wFX0VDJ5aS149k7cTU6374V3J2524e4H7J7+RSpsjASfrMqU/Suk2BW1J/GmMdht
7MqGp4Aco8nqavZqVPHADE54G9xbiay8tGO6GX/QWhnYeU27367HIj7ygAnJdHXR
J+cNq9ViJC0e+Gt4bVa2nO1VlEkwcs/uX0TAIj0l4R7Glp2rnow8HqldzMRZKBvl
RNM5Iryy5za+P79eCeExtKs2cfOqK5ASseY540Ave6yom572XED7DqxwYoBZ/ZsD
6J2ELbX01MSpZEePUzGOLu+aI6w3/ExARls04IhsigMCf9x+K8CjXriQRPEQY2+c
PkYq4EDCe6DtheL6c5X5FH5g9W0ZgQZOPIeB2nrqdf6nQhbMhH6MhLy1U92/FnSG
KLXA2VsvbwshY6QOjAd2EdlY+nxSswUCK3C/3rjhL35hnB37SSXko+3jDPrAs+Et
SnyxQVs02xYfBx3o/ugaMfPvGIsNoPUJYaNy7S032Gn7tBm/fYiBd+JVPJDwQNQL
Iqg94eCy4i6EokTBQuzTzUQJIhq8GaqIOB+Zu0qW7zjT7Awcg61yXfN6gIw1yFeL
u1lxnURamhpXOgz+yODjcE5mTFQ8jWfFDRZuh104yd7fKAd4OQoS8pEeagxGwjii
Oo/K0C+ItOH/SO2RR6X979BqTrs3UYRPQPDaDxUTZ2y0uS8hfRiVjLkiZ9Fb2lPv
ycOzXzMMyViokbLUM3Ey3apUymGJZyGaQcGNEmDRY1yD1bN8reB+gOe5dgIv22p4
Om5nLBwV3upjqye3Pb8YbQjkQ/IZbfsWrVANFj3uzl/0l0OYX1SmJT1tUtG/4pK+
piGNNRzOZopQIYGHizB6NUleQG/U5I8/po1APUSxiJfwiOTRk41bKnAYfetxcE97
QSeZGdux5lfUnxDecG+qwROi2ObN7Qx7KYWPsNMhqTQIlqhqU7SH7C+UVJK5KOhz
A9R0lilhLKV8tJ2IXVcHV3OzXsr4PqOGTZ7vHda9Pd079KcT4JxHzpCV5mwkWgXT
OLlu/f21Sb9OriJk1hmi2CdmZtx4pUIK6V9066X66lKoS1lPKq4XFLloYnILXwWC
JKuR8YBrooTzVG6yJvg6gByAL1e48PaR5CWBSolWn4qddbG7Xh+5Bgamx4+3k/41
xDhfx+2K450MK+B+4wFskJ+LDgjqKF12h/DJTIl+wWbuRNeEX6/32/JP6DBV1ECu
ZrgpsO2BEzHtDruazsbE9xKLEQupIcZSbF4X4nuYpIKKYTGmq66/cLHQ+EvBXchO
3K9XUvZK1q+6GvGDR/hekOd0FM5us6B0LyliM8wxQjgTfbn2nGGrlZgPLflpgO9G
rgZhfyTedKjR4rKw7Qxto3QRJ/XVQRjfSNbratufb0Oo3z0UKWyL6fAGltsDIMun
3fsWArtN56AwPRygE6hsbdUg+WMm3zTDX/mH/6qazHLbvIZqjsFbO/hneInKeoe6
7lKnn+GX2PEA69lDnQYs9nn1ItORe5VSsScK3s+njVRUpcKesIFqIIlv5W5Ql8h0
MNlx+KugjeFSIpjav34AWOGV5GSD6hpLFmpf+IvadWx1JDrbKxNFw7wbHxZnL9wQ
MxDyxwypcAN3m3theDsZ+oNlx35xB0ZViU3lyu0M+OFv9xRduIG9XymcmGJx9SyD
HmLuK5dG0ihDCATh+EuuHYzsl9pmhqCEvKIUJQMfxy9ZFZ5gRm+b602ueDRZFhh/
F6Mj9Gnar2iqqc8KUPwHxPE0TfmG/PBK1txns91i5HSf/apS80Xxiybn/ZeZbZbs
4sdn9suI8ybo+yxCLFlH1R9VQ2kWxcjsPRp43v6v90y3df7oxA6/OzIX78GKP1Ox
MQdMjG0iTCQf8pkjtARm9FdN2lXUAYPirXce5wkoGlyXO8mWLjGcuJAbLYF9ZJo0
NBV2SKYJRBVEqYPMwmfx5sjo7SNsMbz9v8FXzqiLotqeKIG2gKBwsEpRnRbcvqPn
Khiai/u0DEnLPRBcLlzWPdr4gn4pXOWGZ3b4F/dYxOnSfEhQb1OlGIiuv/yCqHGT
+lm52F0sqexpklxr4/j4Y2jv4xrkuV8eECW3ZAPMIUZDI33VYeA9DdJJ64krsGPV
KFDarD64rNC3/PkqmFLwYHK5Ei2fxbSiAbyDXuY7xXMPB60SDDcDHcsWZFRm7cso
W1CbF3+XFSRUWaD3J8qUlZTWoNa1fCwbIG1uCJAyckQ1kuFtZZR3AV9BnnvDSrid
57fi998slD92UHUCsDz4Cda38XM9SseecpjBHdNIU+7BXSK9WIwuUS0fGgJ9I6kc
iH6ylztozQpSuCpUJmkNT7oY91WEDj4Yv07ok5ZtnVSUeYxNbDWIPtoXYJyduwPn
LdBE6MXScMNjmb9ph8GWu+RTVS2alY3sHC8RGbO795Gm2vW8UIOHEvdZcEoEEqBe
Uk592vUAZeGGYTp9pIA5KAPRFwfwvS6bDRc6ZManhgXtm9nsgQen8bBNVtVf1jtU
f6AwLbHKY0wo4CEAmATetdwoiKEY1sDJGWMSRof3XnDAcoEhIJBAWbhvIxdAxW5H
WdW2LZWpsyH0xzEuAjw/IJussSIqUWOrh9qolyI05jpHmlXkBhgrNdelddmzBVD9
S1gc+9rhOEG7QHEPn7qvlwsfvpa7I4/wzeNWKqlXnCldQ0WBAcI1X+pKx7eoEd8D
IE/4w6ZsSgyEokvMxLasCwi60khE0/wW1VKxkhYqDpf6Q8YqsXk8QAAl/Z+CdD1S
ONzbpYFN3vA+eT6kC7E5ViTcBglDd++3M2kd7/5AWTvSpKvAzxLC77hAheXE8NlG
APsoSRWtof3CMxRADzVlluG/kN3nKOwoh4zcUaHwpQEIbLnfKAeYSQKrZkoFQN69
q5XQ04+GGyyKd3Q6a8BgXwM7C78qFJzFbV1GHBAU2EjgWN6YSsfP+B8QXubLuOpY
LDnhj6ulHj72JM8PMUVnAYU9tQIxSK5HdtkyF9V0TeiYKaytriSw5JKulVmsB9Eg
k0cIRajTsSPjy3ptx7V5hQNJJm7X9bLfKpq8wVhu5mdF3YHdDylbGAePtwW0ui/h
0AL0Gbahw3/ykgdorZTvWbYn8KkTS0XzdsPhMC6HaEnqv2Id50QPM8RaniB6tAfs
ewq7UUmYEc479aeu2ZcA6HPHzRcLFS65EeO2TJ41d9H2bjFAqeoY2YJkheDuIiLw
kCcezD26FfgoQVdvTVXjBelLqf6zRpg1YT/+vIvgtYromxukuj/s1kwJCmu0jArC
Bu9h9M7zMheE3Fq86FkcCOMONDOGsJHw7LLLJkbgXbI=
`pragma protect end_protected
