// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UCOCRMVwQRawMJgNQCU8bJhxZxBi2CwheRFQZFwHZnmzrQwmFxbdZSevYM0WnC2t
d8qmlvigfbBItIH3a+E15kNWoatbkba+6809Ew+bc7+bEDMBCejotzSnEOL1HVTU
eSXR2M2B6R4/Cdz8xWXgXKjvJimIgjWD6TErY6Pt3TU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4688)
PgNARHHLQH+oskT+rj95OoZFVN3/pPOHVwyJ44MlLZs8Mlk41urQwNpC5E2A0xy0
s1OonQR+LG5fWjI2Z7hyeKe8ZUcH45mG50P3tO0ZLX1ZAhKB3xt92U7PKCGcg9gc
d/ydKOzIH0GZ9pDAdTIhLXWNFa7ftSB9DnXBq2cAbWaB2enmX+m4QleGXoKwuAzz
MFgdYwgoHJVdrfyhM7Bk96/wRT+aunQwnERfBAldjl87xk5SOdJIIF8x8dkFayqz
MQnyWd5X+W0IOAB7McG56Pmfg+/QJB58IxrvtuysCvNCSb7EtLmD3KBvlZTuRnnc
4U2vTkQbjH5IfQDekn3z6xqEXsszPXdMUNz4pRaMO9rE2MmGHpO8xQLH6rtm/YSi
eEWyfWBiNYrGPmXDaBnlowj7LeoIvwZ7dyQLigVKYDiLvzcYKri2Mju6MlljohR+
AfoGmtzaB+62hmz3kdKUxBJgTHvbCP92jiNToZnK2Vpr9Y2F2QGA9GM/0qUaS8KW
j1t51nT5y0ADlhimnhDyyBkM3bP4zEi2Ven5VacN+XXba7MC0iLycbYEJXEGE+4w
/mUZ8xTB+AxZwbU5ovVVONJXQ6ZdYkk58ewZmZkfqrGmMuQA1VagiD8A23wXrIwd
3F8B7jJX33jfpY+48EV6CIsC9D0b7bj5n7PCpzPZzYYUtvVWslHuLa9v6ByOq7vC
Wi+L2f6n+hy4AXOItdvWaug4ivs5oFVsHLpgIqOfL1DeMMy+o2dt3L+TT02/I5xK
+2YxgJ6lHAwdnwNU5r8JdDZij9EmxXkar+ejhn1C74PPVHfiiv7n/dA6SD9Dr4EK
2YzEiExLPPpWPu7OrZ4flEzjHrcN+Ic0+gE6ZxB3iVAOCrYh453ojjhYzDB60OqO
HIQsDMvWoQPu5RBbYBCNQyg7xIdRik92Cj1JuHnbaXVHPzG4rDA++z2IbzXfpenL
AbpeQwkmXoxUSUChSmiCvjHSysYLBTnqLGABPri+sIPcDhtuwdEgIoNu6RXSF3cS
9CrW4QYgaGyLWxfh+K5X4f+DsFYtcH/sL29Q7Vw2Q8bfXMt25sYgBoHktgJRYy6p
23h6lpsPLiJQmoq5GLAh0+FXEJTzbY4bZWy0/Rl2EpQDUjFUtqowxrPGNCEhU32i
eSGMpfMaMoq79xnrgXSOu+fXzPlry6ZgWWBNkSaPyKK94sFP0+wKIn/YCLhVixJP
56s2Jxy8E++MhOn2Vbb+6eB5G2rQtxtdC6+iWP8hoZHL2QxIa4fP/lUFARI3b9KL
vdyk924G95oT8wPTuuvnJKesXV9wBXfC1o8Z0HqflFxENRYnUO8DISshg5HflQEG
j/SecPr0Y5LZpex4GphEEMS/f5m0iRdGXlpdNQIkuE3oYUjUz6peu/CXwPTsekya
czQH9WsNcGhN5aY7rXc2MfofITkTsReeFREdKHelj90WAcUnC1uYkSd+ouFR2umJ
d1wM0v9Gpg6twOer5u3/beRN4Rk7eRUbx92YfQXbpmBau9k3/8wmp62NjMvdI7dx
3k5044DJPj0xKt1bP64oTwmMHKny4lccK4NN5BuiH+GPl9uT4c0s9HsDFG3tWkcx
3cA491hyWhEJ/s3OgZaAr0xuui0yyYhzQWya2eWVyYnReEcqimCtuzGzfQSziHJ7
M0Ozq+xJO7Rbx2FtWN2HR6bj4pxcGZD0J+r56CNsdIkNJZBJ8heCkh+dF++COtNX
pKmq2uANoR2TucDpjUSL6NeR1bwg14gg53sqmq9P1pIpreuoOcvTNB3ESglx8C8F
i5r3hfqdkm/C16mYvSK7ZZl9rlyl4pHsx9voCaCJbxXmiYyeO02LqAUDlRkhTh5t
lb+vF6M5f2l28TZd91aKjkCAtdF7bLak8tnAqS41LW6JaKm4g/mYFGKP6sHwfIkq
t2edbF1f1Uy0gNDAOxfr/wWAQQKgqlugOtAG0lKbghPNsQevL62rd8j7tJw6e+4S
iIcN5SU6ljRphkUwVLuEMsY3MEy4TQRG5ca9YTXLrYNfpVt31wcyvdsZPPHLd25n
8k7vi9L8jovKTnjMO1iEaPlUdeGkFDSVim+ZB6ODUihDFbhmoQrrAS0f5PCor4a/
JUgyYpAtJHBHjJz7FES+c2wqToFsxp56vsx1QEWc7dRkyeFmL+7kDb2+fYGBoND5
7dZsf24GMCVkxAOOD4JnRu6yOUmq0eyzrVUW5o0/z/1KHn7rS3PiQygW47cnSKfj
64z4RsYm4Tiggs1KA5+d0pwi1elx5BdvkSjCKZpHVRSxmOsWoHRyVJ7eWFWvNAmX
8VTOmADaAZ0jNEl48oSj2q59HS75Grvlr1fysmjHrszGBCvWDuQNw4/lvlaQGUJp
iGjj0Gd9P1WgVxs2AmQy2X3xjLOHvKOK+b5yYKKv7b4gTEKEa9HUM3Sxp7KCl+Sv
FvnJsmq7vLPoFpys5b7bb2gqd6xKBO23tC8dGKoOqnilxM6c5jXwv1dFaAPC/d/y
v9SwL97HFkU/DEoYBZehtHEhdxlyA/byVXayFgU2EcbfItRpEwNMpk47vMCdNYHD
G2LHm27wFbu4loOC86FjQtacDbegnESR7F5Sy+uUWMsuL+cubPVnq2a/Zjz9MT2R
GqAp6/aaeyTjUGb72TUWieoUwjBiducqmU6EnDJENA7h6ihLt9MoXz/JT0wIvRjo
hvwd+TyewkkYAUP2v9wskFGQfvFdkkRbQaex4qmqQ1D5IU7Q4JhPexLSwoIx8548
0Sz1fj4Bft9OmcWb8+/NlUthpwS3Lqp+zco7rZDuO24sBtQK++X+yz0ert4LLpvI
e34xr13LC4VZ2E1jeEsMxlnpoYjUVKPP9z5sCpiuYFpcvxzlYmvwtRfO7jx9W1YR
ZDCw0XQNnAvYNF7qiujcy2xe5HzJ2qssE8cSh0oBbM0x3YL/E75ktn24i0XjeTgN
2R+HwLYQU1G+zoxb+bLt6yb84DfxjcUzqMtvppNUUCLsoLXplOztXU+2K6f/HnWL
lKP/yr4wHOUazkBgMUrQbDFjRSV3D69zVNG5hyEyqPDVvr+bHNDACokGv9t5l3p3
DR5ToDTzUQu6SIvUk/2Q3CJkkbk9BCxF5nktqiMlXoNYf6TtOYd4SDkbWu3CgDBv
N73fCAkztrA8FWsIy6RgzRFXEy0hkYmC0r0c4E3G0tGeSjp2Rmtwk+zuDKN9cD8N
vmltGqqzGk6zw6ToslGlxyUlpxo7YoNNVu8kjiwZu7zzXdsSdngFUdmzSfKSLxYq
+sJlvLTICqdM4Xxu4ToN3cuZ0nsapDQay62+VxmJRZT9Q30oXF9HkEij3J7E40qq
vldFNlqGD4YA65EJBMCFqba6/z7/gyanmjJxaVdDvJFO6n+NI5CG2j2fM7TcJa0P
zGl/VvuxB3/8sYkEcljdl5BVTNThKI5Bhl76900yEON1F9ESXAARPwbj4dXLyWcx
3d5nF5Ay2tmxZXccvyveWu6kkEfdEP0689tn2XzR2V73wQBEP33hTB2r5+1Vukqk
+GhQX6OjzyEmM7hO0YAOLpAjAjLHsyGQpX1r0iDGLhJHWNXblGA3jbvZGO/TcLBy
VLW/hRyggpW/isI4ehngjOjcwfLzgrhQ/UJ0qv9H3MUiF55z9o3Zz5XIEPocuj8F
GCR2OjficlgPM5V6nuH85knTEVHjNc0XKWP7a/KXUJIaqfkzP8wSRmX5WuW+cPLq
aYRQXcZJIm38uv6wTpW4qnCDsg8s1GwxvpHfrJL10hANcD9R89WAGfRcpAfVS1lR
uuXiI74tldJJJ7KuJ5+NVROj88bjxgBXWujM8yGkPH/bMuOMotygZvEZwIo94knV
o1MfznF4WKagVSow0v2/F5EeVdkPW+ucP7CPLwvMN7tXRXxcCR9iHStCdvZUzMLr
v1jLh4+jCWupG3AC7BmcoGAiqSoRwCBWEXbGSW4RysaqMv+71cCAD7ezePhwuFyY
yzEZwVihfdSwmc5rmNkV9ms3FBSs48HNChANNoVYylnG1DK3rx1jnwARsZSHaa0K
ps/mUoUeXKLkJpeT93Ba+jq2AxHmtFcrlTyv6lhHsQlpfc2FTD9IXfLIcpB3Rd0p
q4XIp28mOwIazyp57nzPpkcNnFak823xBoEWdCmpkknnDW9Iz+5BeeZegXvpfHOT
dszuP4e911WEs1l+Dyu60sKaHvgV2n9PNOziMWshuWJYwkJWRyQ6CeR23thWsKrv
d4os9WgkP6Ywl2jlISM7Yj1GIzr/vxt3Ss+HfAAejZrlj8IOoneNKuENpezoP7qp
VqkzVnK5CSTAxciAin+vsCdIEBPD8VxaiaFbsuxOrkt25EePifPfPED849I6pVJr
J31iqDdkTPqYyl3k7qpFWFSprtNeakNZLqDO0YJhTgK13QxmsFaVF+wD4Nbgauxb
Tus51Hg2UJvVi8O4TTMXJv7ZkKWYDQOrUel5a7lO6W+721Z8CXtkzKcOMRSpeOh1
zCYkbt3+mb85u9oCPEon4715J71eQ5LrB4Gl+Rp2ikCTm8nWbaBc5N9K1lyqgp5i
68BL38rYnxVTD29XY5cDo9EHSlI4IIxwqV7YdTR3YNbSCjFgaYsSdUK/rZ/hh15h
DkPcMFfKY4ljIAAYNw9fgCyA8RZuBw2+qo1juATO/Dy+K4Q6QFq9miHi9tJsve6Q
Ii9/v4KijDUN2S+/pCkf6KspFP3LLiPF7Jyw2LobFDQjtQ1Bo1wUALP+sS9GMM6P
KHRY1LV1DNLCRLMoJpQeRjEWpSrn1y0TNA0/vvDuF//ZjGw4n22yb5KUVhsxN463
DAaHpgzUUC3V7gkeWDZ61GsSY6G7SigLWXDE9jSmCEPb4vAipVtIJ70o3pWu6Qyw
0h6o0uf1LJJuVnsRFC38Td0u9raRj1x5oyJPV+qhKjHcBUfQkhd4HeeOzsFsjd+e
H/b4TizxeJWQZo7E0IZPo2LOUZZt/K5U+OiZJW8xq6oEnHmoN1obgX15YCNUZZGl
4dPZlVnaawmIv0AGZxSnO/2Bqj1sty4CzgW+NFXzHeyO8oNI+QQCX6+ssHw3W+O+
C1hP31cRBpWD+MbnHEzKIQQVYNquKg6izyH/vM36Y7FS+GKjDQkfMYEuqEiEpsXY
zTB6CWy+dziVng3ZMWTA4rVHk58pbxqCpuvk5Oyuw8dcSuq+UpieGZw09Vq7TtZV
FskJ7WNrUYNT5nLKpEnSz+j3b96jVx80g80kR/dSIFfZtWBW79J7LLH42Zf63ZVO
ol+m37Ezd6y9NNtZGiNaDZ2EOAuBd6oGFjF4JMcDA2gcWmRRXVt+tbZY/Cts7kLV
i6u4Bi2aISsW+uLrrK+qtH/PfuSupTrKV0ktWI9a9C0+/frhOBPkxnMdT3Q/CvxT
8u9ridhceKxQQzWGYkLk1M8qM4GUSzAhoqOs7Q39BnfICEDpwH2pMoc+LBkKwCk8
2LE2Cv8ZbDCu7BJAiB9RFyoFI7TWwP+gMGv+L+kFeLtFZ1n07WZoKmgzX0VhKrZQ
5FjnxevIoTPZBI5iTHhatbu4K00sVl8/LEnV/TECHAU8gvYVrAOsFmacTjc9hKdq
VJ299R3bkKzhC/sB6AQ6z7A1UltmqivlMjxkvdfpGGPWTXm9e9KoPSte7ATNCP1w
zs6WDPu5+Jl9SNGRNb96xxdg1Jc8dxwAi3AUG4ffZMCVOU66FlEJhbNTQpluZRbn
q4pEKdHBq4V0ZOVJAEz374ZCFazuIYvEeCIVGjvjKAn3n9JRLOJro9wW4+50O6Uv
+4xEyr7cElTSS4NP+6cfj/DYIziq1A1zZuQBRQD7QJrFGsdhDoLbG0EfFXMh+JNi
E2xfkK+Xc3q2mGIXq+bQkcXGEN1by7r4zSMQh7LlHzk/59J16gTpuvqgXJcqBjzC
LO0feJyiTC9lRehiUeRtutI9iUKook/NGdJ/6FG7qUEFj31/xeY3wT8dopA6SWcc
x7byLbtgcwi1ElXiz79LSMEq6//293FPk0/IhSShUSacfWM8OB3RW6R3w9OE3/Rw
AHT1jboFhJYwPHgnhQy9kXLcbVqdcQxSeW13dbppjRWgcFe+nhGqBECnSKoFHbxq
91oNrZZaL/Lbh8VQgfmGaSD//I/Y1Qf6STaYieZ2LMWz6GlROaGgGBfjRdxL44FQ
Kvb6/Tr4j1Z6e5BaUu+PrYiXwaFyd8ZsCQxQ/69CTIPMFmA5eVhJfJWRhGfPBSy6
CQaxZoDvtRfY+0zuugJh7DTrZMArnwGVcxlOe/jL7cA=
`pragma protect end_protected
