// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GbI2Vk//goZSdT7wcvolg5VVUhuOe+pxiqAIFfsppEyuEK9ykM70oXeur9/vWaIE
6/yhGnn1GgjYOur0t764okVOWoR/Iie8rHp6Nh00MyxC4E436z1hvWtUmL52KzCS
qj9umSZSVRURkTuqTtV7LaM/zL0WL71VOgtYCg+v8Vw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21984)
mWJd6jINvCOoaxIe0tMT1uONb7UDIRqXrZLuQhGqh8E/TIqAAcEsgKkYJStA0INM
4TcRQhwZ6qjSy6zIPBE/R20M3wjaDf/R8Fo2VNWp7cC819dJi0BXJb2/cU/eDes7
y3KEHvXuXa6X+Op6iQc51VuWgc0ZRSsWuzc8nHDpGuysqLnH8m5/N4pf5E8N4qik
J0mHAjSPYFaVhcr7x4IzJE5UughOpV66aI9Fymsi8JIZj3INyjw3Fr57PeWvZnyP
11JbH9MRoLQJb2AwbacZtDBLcQogRHFRwftqk7jJ6QRDzgQ1xslwNnuMpQEjqh85
cP5MUiJY9gjd+mHAU390vi0A2iVMDB1CEOX39V48Q0vU4QA0ty3nsv5GiXC5ofUm
lbcHN1YwQIiAuiq5Lhv/Xai4EHPzdul024EvlLBqG5miPkrvW/JzZcGhqB1sn7ej
ar6I1rqcH7/sHl1nUl1wL3gzJCaGiIOmSp5wMqof74T3pV/WI4JlPL+CyMuhfjzO
E3VUB9F/OX4+Mj3/sEolQ5V4l2a+AqxdutSC3H6Z4K6sp95iCRKM08dswch5fcIj
ARh73abVnyR9rqzeyqFoawKHsZSfZHdmuJGJ+5ru4ghIrNttMy0Qw5rsD5S6ZK7c
2ixuNpq87RNAulEu/dm7zp6aOGNTD393WMPw24y/NmnafWm6a2Uf24I+z/H6benS
YVCmePT8g9Goeu647TS7z/Krtpy2QhuqFyW38YV5Hy2xBhE65rsFrj7/T+aJoNjp
vUcUBwKrW/YwI8aMwcGpLemuBd5IZqRc6auG37/2SgdluwrfhLZuUpPJgjlE3UzT
ZAzx1YMc9kjR7y88hfCak+7sHk8e98g7SbMAQZ1Hq6y4LI3EazNLU3LBpTttGGPX
Hg2AD9SVlFDBA5uquZVAv8ppl9sE/vqPh5JkVzzHntytPHkLvKRqvoirXxOyV3KG
8cbYJ/do0dUOx9YipRhQ6YVlbiuf2iRbK9EhvUDUECV3h1n9g/gfpeoXE4WvvrRQ
vmHVoAe6FYw9gegKBzWoKw8be/TZhysPpMlW4i/zV/LUM+GOv+RHVKu8wjdB1+6A
P0UfdIP0jxvYelkCgWUeW2mAWPFmHrXKXStVFRZ+4MDIa7cy5TTOswqMW5v1pOqA
cp3RE4S86oEYi/L91+EMlKRc3kaJuU9UjxXurTzW0HE6IRq7mMQCwZHg5EEfqULx
TpSOpiQ7sBZjwLdnakiXeg+BFh1wFUdVh7PEY2hNr3uYdXOO8Kpw8JHKFts51JRy
Q4+u1uTTPSZu2NHpSU1tgKYFj5bkhvS5d7gDA2ysWUmzwLsV716JxsG3hfMbHD3E
nTwrpkCrDk99gOL4qk/G/nJW2tbBON/4N4e4Al0572rOk0zOlvHgEGPEmKcikw7g
PiDMDdf1OtowfC/VnG+y30FylkQh/gv8IWcD5p+dWksFI4p+ClHhnZSyUdQ1C98f
Q4fhnWu5V9HJNnDiVFLgbwxgk9MqQilxddfNYsfsznr03+RkfeCPjz1L7XaCgug/
9ymG19qOL8ELGl17yzhA2ohGX6N7Jhv/GYRMnMdzvxmbizy/+ugXIM2w6kKdEPrY
HmoVij6VZjynSfk5KfaRx2d+6GTTfKmpaWuYTEjN5GPkwzs5A9baMBmUGo2IGKn9
aVm7Zai5hirwByr4eFdYzI2qGCqnJQ3CLx6UjLr3/0BlBhTT1fhGoZZGqfeOtvbx
zr2jL3BbIp4ZTYzx3s3InSRjzKOjZsi4yeWJPDhWfKzLXw9mHX2+ovp6fdYrHqgQ
BSiURrP35pmNSfi4GTVd/mXpsa4OywXtMsol0Bl4B2fYuK3nn66KGHSWmGBashsI
XiZWHpa1VslVEjobFC6yByZdg/2CKgqAeWI6BbIBX6D/QoDR2ICSY7G9kr9Kq4Za
QxyfxcBx0rUW9VCDcmxzpSrbd/2flVIi2rN1PwyGb2S5DcHg2R+tqZL29g2hwoWa
wevkhtsvxWCZyCL02Qs/MoPo4NzFDvAvjnuXgQmkeTHOYubRd6J40+GdhXgd0F/d
aS++lZHDq2a+6ZMqmWyKuxT7CV4QnRb5rDBvecoCdUurUpKbalypADsU4REwAgBb
4amP8he6YdFvI5zNEGTiSONR2iRYqTjg4GCYf5SWw0qTTVfYfV2rt3BKQ9YIEdoH
6XVSsx0iEah9NahEqKJ1jt7OhgLJQNf5B16FbrAXAKtakAfNyoAjwLGWDdnD0HtM
1uJf0OroQohs9pabtPq9BA+GvhJAGEn0BZtMf9RaN/DwZxl7bInQ1+2bCCzoaDsT
gPLKEG4LrSteO9ff04SQ16cMwsXY4Vx44FW6pw6PkVeHKBx99nQ3kn6kM/xNDijQ
qftm6TsCWs1tBL2YL+AR++UKzx31CRMi5UHV/5nDIRXzyMY6KQbUppKQM/o66TRg
tIno+59yVqylTSNCn7xU5Pp2mdeuEWesfwCCk38Ungmc87y3G4BS2/MPAV8jrpBB
IrpUikCvhuvxJrJC0Y4rge8Jiys+HZEzXu5W+Z9vbhwTG1lDagn8OqBQqcXkDkwX
aiGUX6ZlN3Og8YqvFuXnlLGYVtdN5JkWnVrYhYfNABICKOYa7pdXXk53+w+5ZkeT
IaRF1zOXH53nm49CZQl0XSC+PJjWPP4gud1lAOpNmkefWaUOV6u4z7j9e12gjrvR
XCjawwZ9q3i+luR0LyaNaCmZbBaWZTS1DfrO2+Tus1d6d/+jfCV1p13gVAwy672m
IKZsm6PR1VJ9dyGr8fzQNKd29x86SWWbJdbuYLrbiiIYQJcl1pjqDGqHWU4Ad+bh
EHpIlg04P4l7kbwhibDGEOsJBRKhV/Y8jlPU5J04bcTcLKzZIkEqTXzOna9KgpCt
IoHI4hRVmwRwCB43nMn3lFD7b73VHVvE/oKVYeCjiIkHrfTFkjTGn1xQOLN5GPCK
OPl0LXrLV2f3Zmj+Xq+iIdjF1EKTmDLALDryP+QaAbOFtVvj49oiYZe38G4wP/K4
DneNC5guw8VSD3unl+H8DqFywVT+tUmvrsZwXcixwIr5goulVDSmz5krO6Hs28Zz
UcegrlazddY6kMH2KvrhiqrhqA8Z5CnVZh/aOkqd+Tx5vXjPwzOaS23xC3eF+UJ2
aEg7FKUtvJROUrXigJCb3K3Y9PkKzO3u49PDCLsz/al2TUCJdEsJ9V1YI6x9xwch
xx382P+yt56KEd4rmv+WjmkNrK26mGUllyJSkV5xmmS2eiNNaUdzdlV+yoCy2E6t
fhNyZAnTZNHYyjOPi2K8i7DdGVu17P63zCE8lP25LvrKsCO1/eHMmmUcsk9ntr3U
l5vsYKr7f2y0szAXyarcWJA1xdqA0CO66oT6bBzgpNEF4hPn8I/VZeXY1eKHuNzd
gLEy0snxXNZS7cBvbroOJQ/YZq2ktd/UuGajWswPRCx+2yXGl6w8kHeYATNOaX19
losjxoXT2GdF3gk9YufhT0tN3yaHIF4wo7jApAavwecwSqtxpniy1wGYJCaNklKd
AyiLLGWV8NtBYZ72z9S9oMLA/sl7NnIgtqsuRmVzzSmUtLj3RRHKdqhcEGfZzFmf
yzFf6Ym77KDUEtZaSQmUCkB5gTPxBwBw8YLHuVcBxu0Ipt3h3Fixk6QzgMuU6YWG
C5Vqe69GF5ND0yK5NlE1aaVfe5EtAtqs+fLspANS8w+f8gGjdVbgNxlq71dSxTeJ
QdU+ubhfGtHIM961VCw0DIo0SWkKFuve76UE/izJcd74trwVLBZsrJkSOGFS/wDb
1zXaLqjji3uCMQWNWDxn1+N10BxYnupeMMYPYaQqrSpPLvb8db6vs+LOv5T/wEJp
rrANcCy1ANGNajofXhuwzRQF/QCUlUoP24XJE8B4a7XBy3gYi45xD0fIrbdoNkNW
v4RTjOnWc6kTPp8svxFORj17ETq6rAgKiFI/rB4c0zyeR1YJwXeh0fyEapTrOcxs
hyoANMPxpKR+wq2vZe5NYkc1bA7z8eeQcnJiAkYHjappf9JkteykNi7NgTlBvHG8
yVBHpSAkzwCf0XJ3k1rNOfTZr9SCAydBnjjtenX84KNCG9xFbHEDMbJMCvftDAWa
WbzreANaGUI/dgjn0rbzXgrZbyBeJt8j8yLQs5oxd7r+RDYYhW/b1Ow5/IRAf4CU
hKGtrgR0qDZaEBUnWz7fBaPjw/Sr9omLlXEbtOM1fEzYcsv1G9VtZuc41mDv4nS3
B4e3U5abrb0TCLKfPD0JmM0+KZVTortty1R/Ru1bFk5h19Z5eTQ8tBa9eH0Pd0a6
fC7nrtqtd7fLzDOSTvGREX4BEVNPcTVa7TpFO2+KhEmU9gBmOf1vVDWDR9hiQcKc
hxv0rwXjk4jDlHJNU4Iqg8tkIpPXDkb9BETzSXl//9c2up39WhRDgc7jBgMMhdpy
61hUeOfR/iMXltU+huifLS3stFZM8GDzqcmO0mnohLqeoI+Fq0EmKbz2r3x5lYtb
SueflwyCYLi/GwVYvYtfcJLna/BmBqNbhDea0D2Vv+UGjzdh+Cwarq8EdwPNvoMx
TICUk9XrHHfPFx99/EkpICTwDVQiuW1wWi/VQJa5vpzBrkjuMWEa77mzCuKb9LSb
U6WSht/bqx9GrU4LNDG7NJzCUC6FCXXVnWrWMgU/Hxs3QgA2x9L1IWlxDAJIDpga
cEkWxgojI5hyLrSYzlBnP1c4g8HC9DAs8qyKerKxdyuhecQza3/+JCTy/tpMqeud
+pN2zzM/LYpOCXcCaVDU0HGHc235iAGaf6FU9JcxlJzR6XgjsVsRHiFemC6QLLdm
77ETtrO37ISg5yLv6kIwSzkLrI2hm886+P5DqGf4ypQh3GRwSSjx3FV4NOb9lNg0
kUQjvgzDjpaiuX9QAXGhdZM9ZwTtt4wlPpzJAqZ1gFnP5yhWrnU0HLNMwjFIH1UY
ZliOfMgUAI95Q5S8G9C9t/kYOzaRO1K2GjXGKdFom4CAYKa3HWAp9pTVbBE4DjJw
iS4gSSsH/MM8vlcRzptgaHYMaV9aNnqDM/UNYiPvXRHjiufWtYddpwZTzwmjbkjs
qxIxHCOE4QOCKSANIr5jbFWcDmju8gwmcRdUEmmF6uLwCkclIRTPXyuzoisfn7yT
wHz9dFvaUHESptble+LcLJmKWoiUPeMMzes1JH9xaktPzuNEpIOIFS/ZeBDsKABe
B0/31YFKTiqo8M5n25L7YauZmshUYo1eMHkGGGG8DbIAdrlnTGGIaDG5bKihCIUQ
UxYsXGtBo27BVsHjyFSN0VCEuSipOwYpmQqzp0oD40S7eUXw4mZwfBNzjQ9jpmsR
PHPgEOlVvRn/RS2q85BYdIVd38K8/5oeg4K7RbYzbvMzuv5ik3FQTbzlbWHcempS
mY9iMf5yN4apdScvXRsEhfH325lCMwpA3VB9gyAf2aNyzS0uQQyMUAhZCh3NQ/Z4
23ss7tBjqmUCk/kz/5Qb+dmqP9MI/cH5WNj9fbEkgsdfhyBL9CN7FqxrWlpjiQ6g
q9I+ZN7rBO7Zw/a0piizJGJ5OT3SqkguRqO0dYRUdLfwDcZqI9YUov2O+V5Izzve
KW7kMVFVpcc8PoKSW4FTdXDLOJFCA/tGY0m9X6v4CYhr8tArhyePLmr+upQa0jkf
cXuhVigIsFvIdiZRlYn1nZ1PetRqktvV4rG5Vn8KrzcPQaQ4Qubm4nq1WaPKPqgq
eB63IYgY748u+fnqkf/WKEr5ZMLrM8Q1Z86GWKCIattfg4j81wAwHREW1oQF10AR
1HbKDhaNDkvqxs99J/9bQdKmtBmS5o28YPFvgRlEbK/cXcX7D9eCfW68b6pY5CHR
jx4HSUPJw9/ccUYk5LvwQ8EUGihc4DnWvi1rs6dcDzzVBVc2aX14f5RJM/K6Y5HK
bB3dywZ6Q/SiV4Lq3m176xxRVIMFzT0WDDUh/gwt93VEj5VNurkdGYDZjOaTlgb7
VGAr1Dm6dLFtKy5F/awLfF/r45isitHrPsfq+vnGhdjT8rZ9zyATJNhM8t1bc20z
IMtmWOXfgBDtalTMxZmltCiz5mEFbp6pap/b52LduiR4DfjJBgWZ/x83lw16hWDO
4mGYNs0god6EqlxC/D74h8yB2U9DRyv7qIUF+FVe86YlIUa2Uizq7zvSQ230m/+P
emfvX1ZL0dx7Z7bRQEXZTawlbBKgUv+cNAOZZFGGkeOhuGqfdNRQZ7BwtO7AyGtc
QqwZF4sr+9WjMwzIvdKHiK2Yqv3mSQNQTjAid7GNYDTo54ejd0iXBc2qLagbJ53E
E1j7C1Cix9rK+NbIQCvQ0VHnOuRFw7Pco78/4tPyc6OQDKCxSfTneR7ftHv3NZa7
DX2oyuScU4b3KxKzaqb5p2386ki75BCbrxPS01D3xUxHm+LbpVpj9GPzmjE3I4vY
Y8ORkYZQSuaRHZDFxufvnJ23B2b2cvhRDZMGNy4JNfh19dgFE+82l0WK6NfSkz2F
jz/UyJmTsezPkgvIvDHnKckI9RjY5Rs3j9Zm2+kzocUtfq/kj6EYjenNlZUa1RXm
ug9hql3tH1P8D42/2MAfWsvooJ7z1X4vIHtTU87WMP51mJqLYYzs2/arTsq7XhZP
vD0pRsd6n08Zt8rk7kVWP4ytkajjQslYKDvgQj03foeCHj6iDpN9oml8XixSJcp3
A7TIlCkgXfQ6dekjuFmDiWFEhkYsji0yhm6hEz1oh7gF3FEOmUaQE/imrJ9cIdd0
Hd6qDVA1f+X4cchQDdEOu4BX3jsOVoSHTMmY1jKn9Uv0hVj7eS+dQ1jIQSEyx13G
Z5Cg73F1IFMA0eNviPUv5gV6MqwX+evVBBaOhGw6BdNc/ssRI38b7BbpaHP8YpZV
4y1hNkLesKtenIwq8Mfdpb0hikjHId1hbNrpV6wOVz3CpsL1y+Gp61OrqNzvaP98
oqjBSGbH46IlVTmC8GWwLrg4CLUz9PDkOsXGxHxuNKMC+ikJfN4AGMZg7VYxcjVC
Mds5N+m5yk+hRokJv3r0eCR3HbyCyt/82VObfAj2t5glIc8OOZFy193QPn65Ze+8
42Pwsqi9XcRGhQZHUGPCRXgAWfRT0Vpr5PHiRwrRpcniys1t8h4kShBAFQn6ln6O
jxot2s8BqPbzQPnMELQJWV/JgdgErF2cbXomSAnvryYHRvMrZTwLrr4dajSc9Rvg
RK+aJUgZdUUTOEGZ1VIKYKh2PvxPtEwnD3xgOhfAklY2u5BhtXG+mM0NZZ+MWm45
0ikoCqcagzr6DUjuLZB2jEbSUNPUf+2yCeICZTqqtTDotqr0euBAB2CA+eQgZ7BG
S2zTEJ6h+8tzZwHI+yJTJHnzkMh19Giqpm6yzARPVJuqCOvBW6GI8rO/pKlWHg5Q
M5t3X3KDgB+Ok5a/qOo8qHdZ31mImWmNqTvO3i3xqONbrXJQqODZPve/yzRA9YU1
YbEXSKuwcKfG+hTxfdjyHkdEAhE8j0tNYKAIKyFC23VwLb5ju1WJD79237FNBbSL
d+hDzv6Gh/PyjoOTF+On2lwe4BlV1LdNnjNBDlRVlvlEgqbtS/v9FeegDt6vjyM7
KVMcW19mlf2fgAGpSHAmOwfDNvlpON1gS3thU2JA+SYbHfuc1LvKBmDWcxOdD4cI
BcdRqiZvlc/rFDhqBgYV8kUQ3ixLV6QW5X6BXn1xL50kXnGyIU/mLvjm99Rujh45
bxYdUnSc4j2Mx4nNTzznjIn2dS8xkWLarP05uF6/8ne4hELSHVHaKkFcwAZN27hk
HXZNehaJ21I3ljIDbuKaougGAWaazfMRaTdilI2oMuQkn29C/yaVAxwPxCac4C+L
IlVdPi8WcgXWFdXycAz+O2cIoCcGMRD9CEUUDpcx0C577JQGttgXJ60EDUSWnkUh
LTRX8/S5CgaHwsi+t8rPHks+QM1eiqYwLurj1ocLarzClwIxrw2mEZCead3mjvCm
nQ4AWSi7LGWx5IUHre876uoCMFYaIp/IK1uBPkKiXa0zKGtMUn3nrEZtONPR9pSs
Ltv8fLSMiacITpgAdA7/4MN8XaO9TKvY9nhmsw0z/fRwzS+k6bHeICdpt5pd5Mha
MxI2PW4QoRX/en608GeDPzTka+VO2c5dpgEXAzUB2LjZ1Q2eGqGrI49ack5m3o1w
dX3SmyjhcibXyuvYcXu9L+oCV88wT6q+luZL7gnA7TJMrxbMzSbBz8ISwU1YVkqt
LMAeWJ10Cui64BClEEUfYYFG2tFef9SdASlReCglF8A1OwlO1cr1ZCjQ6+7TVezU
DIKUzdPs5V0OfPVTXNvxKdZHcr5c6T10Z9+YS7tENwHpJgoNPzWYc09jxaL88t0X
F39mMMSSC1ZH8jzCNP7s+WwXDXS4acN49AIbYA5bXRGxAn47kKA9Pulk8psyHeR3
bWX0z9xLAo228YF4Jb7E0CFtsMA0Hu1M4Btjnl2JpgEiwiHnXhV7So03OeUT11V0
zHmcXksMyzQEvHFcLq6MOyq9XYGPkaKP/zrRp98edeWnUuy7smdVWUzbMZvvruX/
vIqVa2LU33r5cVVzv9fAKlMgttqO+zX2CS8iAy2ST2iOCGJ0hyVNxP4qauno0rbW
NcUbfJefI0mGpzUXffDkOQTAUXoc92DWrQV569fAbiAAiZbTo3r5RW/qTofOJzr5
NQHYNyWA7Bv3H98uoVULkKEGEGzuhvMfL56ny/fk0nb/+g3lCVbos5+zJs97IZK4
JrqVGd/+rpV9Z1AKkN4MDxkL05cMpxSE5kA+KUhC/Kg5wH84WhmGrt4YMuF6Nq0A
UVHJ3MaS1Pwvhs8GhSHwd+bfdQ4/sxc/h5MP5Q1dlnKalQOdyqq2H5968uXX+TxN
O3LvdoGpQZSSSsf6ijOeNZRXelL4uGFG3AKMkj0vyCGAzBsCIV5Kfcb9IsPqLDKP
Iwm2nPzbuku6LRqm97qU5UW8J6zl8gQrrL4rsyVa0oLDDUb/MNUrkRnfq/36Rc+I
3R8MG+nnePdBl3EUR+c6AHEb46RTJqJlcooWZbgGT4YOi/F2DadAboaFInjfwZvX
0QxGb8o3SZivyiyqQ/0UfEsgcdbG/zDTTI8gQef69u0OcE8R0fimmEz3n3xB6jbH
4rIQlwWsCImKlJD1nUFMlQZxCDdJU5Xb3f+Tk8e07C7+1rIInmr+bZ5DkUkNijbX
jdZaC4lNFSqXOYIDrRlkC6v5wJ42BmYhGRYTaeeQ0UiEVF0eV6UHhlQCDGyBg+pv
ggyvm3J2vP3DaC3yQ/GBzvWqeW2VBXahh7QxD/VdTwEFKFGoLbdM4xJJHxD4FZcG
XT+QFvyo05JX7VEq52inonbDaG3Q2PsT+w9dq8Ejk9hWCnRM/lr83E8CCOw9WivK
sKZSUHmEoBf39laQ8UVICSUj2bKyRF2CqbSh6xsVBSfBcvCfow+Dy3hL81Srcbit
lYUkAUAHvvbB407rgO5z4wI+ZpvzYQIrl6DWstRnabZpnhTPso21BiTPdfwOMS/A
ujosUN9oUR7yQ+fqibqnd16U+sPkA2Im0RU7AjwbgeGm9b+RSm9MnCxIEMWdTQU0
ioIWNnfgeWgEUQHZL/hI/34c3ri7EffX8cIzzSF71CA+7OEIHImAHs5OYZ0sjaMy
NV5PZwuaUMbzr3HcpdJsO01Ac9p78yCYAIt2+tZNWoCxTW9IRwfU8aer88rLYpi3
4ZzEeWfxbGcVm+Rr0/J3c5iVeQYyWlvuXjSOLBu7yPg/ebSSKcoSvKIUx1ZJDM7O
YQTadcXoTGdUhaw40ET5Ajk6JNQMhIM0C4gQhq0E5VU483ueyCqR6dtkOQR0AxjV
UW8aaVfTI68wWGbLyMPWlOoegf4jZahVvRP8AfltbLc+LQkK4C0wsJvMPZ7vaa8J
V+5DtPLUMpig7AbNnjHgD++akqfobFLln9eNTGrU5vY6RbWMqHVmu2xfZQSNWRk2
SOOX/pVpwvFaDmiNOI4Klog9YlUuTLPyCo9unDwHfDlzkHOymVXe4+0tXZYZqL9s
27srF4YoSSzMvgYbEPEO42XsbqBGG0PCTrynVv+766oD8tmPt+fiK+Ukx6ED5zLS
VJKcPbSNDd+FIOz1JnizUBynu1YR8g1Go+zHhSYTXCGa6uD91xc4UWGenexK6/Yj
3rZ9xzswBkP6jA+N0ZDwNglWzRNwBu/YrxJ+NjY3XRvYUyu4b3lyaLUeiEprEhx1
LkJO0hLfnvU+jOx8M2/YD9ajsPhoi5T2HalLdicHE93De3KkwZrUBWu6NTSGd9Qg
bhEjDmn9ZoCwGjxxMTSJVzaCvdbdSzEkosFA2Yta0VGlZO8EDXncHttRztAjmdSR
3I8THOtnyagPwwmI9ceO3jocBDoK1604m1wVvm8mLm1/c1ckY2d+TVPsLqqfXidc
y7lYfGyil2syfRNdNlAsSlu9pUjSY1rpOdmGw75x7YK/n+Hma+aL11lBD8LUujBf
aHL7AOYgu+IoXfxSTCOdHE00IB0vb9MwuAE1mnALJshSeZeitsUqUoa7VmRWTJbv
LRX4WwFoPsypG/IcVQVBAb/Uw52lfsj1nrqrNGixY0XEvDh6xd6Apegx59jbl0tv
WpqhXbW0XFwdT0+YrXlxMz5zhFt/5I6bSZQGDMwnGxFVR+8NVvdrP/L/4tMVYUUY
JBqVXDOVRadixGeQtMZlxb0M++Zxk+4pk846Ze9YZb2ATodxd02xtE2jWJSEmS3O
t5WpOAAHt21q+1xZrePw423rlEVIhzQIZ5L969FdmsyxzbYVenqZ89lENP9dZBif
HUddMPSycgXPNmbPqVeN/RoFQ2facf2dGslJXLCoeYb/WTC8Omj6TmslnHuynaic
OdPQs3XXH64rhOEgIVYQz67XvqiSvuB1M1yfBq0mjFjoZwd5flhjzGziNoN78o7Z
Q/5QYFpk6SC6P5i2QXo/xT5MnMmes5Jh/BlJN2JGLFs9UajveSSyshJX4o7i6dVn
MpvN89+kzeeRCjIewMg0HEK/H356OxaJAZKph/J/tYJMkHguHbUImu3CWYLxwJ1N
76PloCnIPlil5mGc1ufnILjxCm1+3Ha+4hvsX0ApTsoB+1x+E9xyIX9UW2Ud6yUy
sfhapkVJnaWg9R3ZXDnZeguOVnuzga0Fq5Ftsn2Hy2qxLkpyNTkQQexTMWVjvvyP
5OlB5LnHXEhMBUMY/zeoDfgajJbYHCMyn7WeXNhcuNikHRx5uQo1Nh9T6jMlIDZ7
tueyaRvZJEZfi4PkwnudDuwqN51R9YVplym5ag0/SJc0lw/vishmP2aDpM/lqpFX
RdmyIhIz/LLBICrz9FTDr2cB70MzfONcmqxXs9NYR8I7xW7tSwJEcAouiUuOyRmc
yDAcEI+e8QfsSL4F0EddWY51reZ83xkRZPvCvc+yh76qIN4iI2pfxJm24AOldxEm
ifg+j9kzi6VkmHmWSlvLcHpZYAhDqW60ZNivvkrAUhnzH81TS0DWS1LhHrfukDGZ
P34AsCfrxs9zS4I4n5L6+RC8cfQRI/4p190MyZoTc9lC8zeXinNjEZBAPAxOqFTM
lPocRKkN0OsSgpIGonDsgQXKVwm7RezkK21aWhTkHvnAffHQHJU+q+7n0ADfn5tq
U9WrPcQWNbTGtEqKN19Sv0dMpkzQuQCJ6iEK3ZA4bc3lzIWV/El/9zdEtXDavyTZ
evzjUqnCtx5a9uYgBV6JCdvfQAcvcY5AGbsEXfz22K6TVdkrYN28ex46qwija2fm
s45p4VncHper/cBu7w/M6sY0Oeee9NjZSSKUqZG2czx58f9I3oFniswn+GPFj8TC
VIBg+Dy8djVIruVh3+fZ9Dl0fDFbTaO+Q3jd/32X9D4IA3t4iqF42WL3LXcl0SpQ
Y3yP0eZGvzAlQFJ8TQgttk+2yoBD61pp/g8Sc4ribbFeR6/zLkPsz1kb1D2ECTmO
h3aNZ4jy+re12lspXwzO+GiC2ZA3EUUiBhSQ14QfCnGHW9fMtSgy2cNUhQYneiTJ
B1gkM0BGNhdptgE6LsdwKyiY+UN1fplvzYw3dgsZ0joTcaEM7bQhFLY6AFluq835
qwAHU6jgO9MMR9tRa8QnrCGVeBA/j5SQi2Y5D/IWrscrZfDjfxfXY8HgDAYIEWh5
s29IOmvRW5XfgohyMBCulORi6bibrAusaKrQrqzEuHzeVy0Rl8TQv6s1e41MVcBr
54WfziLu4LtJCwLfJhj1YIvuaICmPmvFTTnAK4g+FXWGTy0StoDDR3xsU3bDZ4eY
au1u+Eo04vsyqm7RGFgU5M7lor73Vs0trPwSeQ+bQGlC8fr2k6sskX81csWQmrfS
kv6wAyJZWCNuhZNwY7XoTOish9Pyihk6ByQ2K7W35nEKXChrqKKDey1k0ysxvMqN
Q9z5fW5zel6IaYX/9cUDMA+OKfXsBTGV9daa7mnVxnUVD3MI5t5hQRmEoJFvFhjX
2SekwOM9VB3Y01yfwLpb0m2Obpvyd3Cg9qAstoy11yND3ZYo3oVLAvYjJaCFUYXX
b8+B4T0BJlgk6wPPXTU9labKtcXJzPLoGUYCTGckL4ExJvS6tyYgBofhKwEKSNIm
IZojU0zCaf9uVyuWchvy8kKPuVKxYWElsYfEbNa9ex/g4QgXQ5GsCKVU0RPZ6rvJ
kdxGZuwg1XC/MPq8VaYV8Njf6Rz9LddagZTFZ8wmyeSE6IIwflmBQPWWZ+/DtECg
JazYE1cbtM9SOrHkh2E/p4YB8juATcpgXql9yKMkhEIKdP5Qy8tAEsTyBXsZGV2i
Reh/VgwcOTBdDFy4j7yKuQGcd9iMXaMnR82Gq39X3s5tDCqj60wr+s6jYnAJhq5P
jvloINsyPkYJK6bgY20eZU8I9Dl1JUIpLUjtk7jgO4JZhYKKXKCVWjSC0/i/mXqf
s6EygyDHgaoE4VJwAKqB1J86PO6phlwsImua54nTB75n3Uc2SJZxabP6JhxFzb9X
T0Cdx0TP5YgDc3mhXndOj3pRhyiwk6I3MTaJdlyS4gfGXNqhMbiZNmBfQblaifyq
YynxT1Lv85+KER/xwT05lzZr8DzHt0DPKKEwRmZ+cQrMQWJGHWBaGeQLwI1FJPhu
0MQOIl7l81/4hITaXmY5RL/l/nfOZ1QZndmZ0qXvrMOMa7f6sNhpNze13d0VO2uu
ISRfATt2sxNcXEQEHotdsdw8P044LwY0KYOnFFzRX44VAnw6sgdyTQHGsT5kYFsW
9zI8EdW1J6MoYI77fOFWMNCI4hx+jlPevhYjE/TEfiVmNZbcbSf3xCl5dQT3QNqf
ZZox8hIusMP8fYQOOnUg5ridXLQo6AvJ4qqUmRdvLvZI+xsTnfqOJWGSfuA43/u/
QPSMkJgve8+/HSJkFJDOhqXef1pYTXBa2OAznu4Im/X1tegRAUSEbU+HzO93ILxk
Bm3HETm1GJeu9e8Ekyk2Pv8IyJF2pRQ2P5mxEWjG7nByOAbmUG8ETXILjJN/0csO
5QsFnP70Mo3z6fT32Eh5dcePFGn2fcaAQjV5Mt23A4RxJynrMoQ0T0sSBgcdRke/
gFLv2PzrOJbix7Xhk8LvgekTbNF2pjgJ0Kv5mZpImjzSnP5yZXTHLlAs6dBj9UQ2
fxAUItJdz1Z5js1DVl73iGyafx/cPLqeZFzNdIEfPj0rJob4gqjXAjfLUzQkEiT8
B+adTzZ5a6pV4zwrV5rELgpSByNm5Tn3xs6aEpjdzOt7Io8xLnomi0oMKMDLuk+X
4qqnEtI1kefkeCrG84iqbkgIFVTA3BHIaRfW/sPfD8qPumSV2MMknTWcpM56yODv
M4BKoFK8LXHiu+SBjWyXGAd236JJrQjRUNqe+znzorbEjrA17FsgJTBM0MPwCNFG
ULZcRNOZyGhmjMUnG9mPyn73q/0ihu9dzz/QnvO69xfAGEc2lpM3oPZmM/ojrh0O
T4bnnLyatylDBSZ1D3dpnMEKaYkG6bTPCIPjY1FCIvPSVc/IsEvXWmgr4cCBXLJU
ABJCQrGHfQuOQjCWScuupLRegvYtsFxhTJsdP/8KbdKWDIXAn2kEKY4Jr6N1gYq1
cB0AzI85i6+T+z0oU+RZOb0spIXIxrcSKNAZRxg8UVzGAeVBBuqbrmq50veXBYg+
cv5saqF7Hos6yFEblCLnYQ3sTY46Ga64nHOYOuyLLH3vCiMqmwvU83pcqcL2I+Ly
uhkv4te9uLPOMni26f4xoKn4nPIIby+rY1J7Orq2b2JHtNaHs3UfgaVYt+exwsug
4g4uuqg5qFO1bshtT+XudR2QvlWYhE6tMwIyKC2jveAzIlMF5aH114ABzVcMqKn4
CgXkpmnDk1soBBMy5QTGqoW5zK3WAU1T9noQHoUsh5kt9Za/gENBdckg4sfqXBg0
bTt7ib4dG66vlHbgF/StvUbKFwXQ6QjFyhox7jXrRm0i4phvIRUVCUdLfyyHydzK
HYcTOMjvSjgEJralDWhhNZQF/eVx5DTT9ZGdT9LeZQ+WoVdzQg+a5Fx1Yq2NxSn0
DUZmSGefE5KBMC061EF0Z0pSmMTvU4xhr3P8n5eHL+WfsGPDFFnQVAXI3EzQFDST
hmHpgW1SMZHLsK2F8HiNG+qPMOMDpXPy+F1W4mhwWLKilGSyJgZVRzhjTCaxDrGU
XT0lKMRPmCbfkajaDIcBcQs9NXnTAUHwXBlD3RErR7ROq1RcIM8X6L2QvQF7i9O/
evxNCbsSq6nD1+w66x2udvFy4CCcDVudeGmLewuiu3dXtg2QMYh6jSOJ+qfXrTTF
hqajidyiN19HJpQWa1Yigray9/nDmBlTPdYAEvZ2hsXczGVsSthcQzf1EajtHXpL
Oa6b/D+YJbXQDclqTe6SMbSP3aTPbo+N9RLUvit+FnguW6y0PQJcRkiuuZAckcx3
jAsTgKB4nldZb21joFwL+/uz5Xp/D6YWhbLRZymtmh2XRPqpS4Il4N8Ktyxsz/nJ
cRPmP8OzELWelMVPKX0OMGIOj6tTDXruM6B8Aoy/HvfgLP8jsY+PVE51fLHwQf2F
rC6I1jX6x2+OgUyDuC0eFJP8abM8jv60vWKe1p6EtDN4cqIcCRGWb9CBzFUzJ9e1
csiPX+ck7hBempMBtEAnBmLRjXXsjptZhm/+xGUbDRdEerFVmM+EFUNsykhNHfda
SxIwqAXuTCc0asLN4V/TRPDbR5JtusEYf+EW4/T9/7rPgbUKQc5LCiDNWjm8X1Ya
orw0vT5T9kFl1VS+c3aA9p7Vr/Vn15S4B5OuRZOdwiLjqr3SriuuPw2Hk5e4qbt8
ymeydEQ4EcWA64UFEd2nSq5RdiRjWEGxyRukW8rMDAXensrr3fUKBU+ODU5by7lQ
r9l4uBZXmmVl813Oqf5Kxn0v7ENJWNnDvBU9upxgVQ1zJupw8jJXnNnWtYeqDTyW
ryWE2x/zsSqAB3jRbTgpVgISU9xZSFo820SdmO1iqU2/aOxMn7IfJ1sgEpO3qfuk
3wqM+u3mMwLjrPi4b99XEHupQyLP4cZfBiCvRjLbHD9znFSV80bS7/bxiRmr1/sH
amuXLJGwlSQ8vpRqgpRsvzpgnwca7s+CZs/jxmfBhIhOqFDWGun13IwOTV2ShWpG
iMYBSofElZgJbAB8A4hyH10y9FGgC8s8af3isbCH6fWRhJyO598pD/cAhUXuG5/u
eCbHyLl5gysheefYV+ayDI9//CGs0DOaz4Skvrye8DVG+3KLDkbgQhvnE5TQhsSm
g1taUhaEa+OrEqpb4teT9/Y8MLojyu6ZVSROIp98Fp6b+RptbEfHlMjFDAPYoM2D
QmDtKDgrpcoh0Szg6at/1oQFFK+wHlXBZWbGfmTFYY/udSlxosKqT0nCvzpWApm2
o19LIGG/2CiwKGwwmDrTw3UNEp2EqBB++WM7itabLwS5IQlkmXMZYi1/ernzFFe9
hbpcBTWpMh4mE4JXdZ2z/Dw+AL5iTJ3OkXEAGOsB/raMuSXc4uWrmxuNctEeV1/H
4JhfGzBMp3jooLcTrgHEI23RRg3KaqHyXKXn7UT4GFth9PCVcXYSBgJ8l+63hNcu
BkvYR0iIdqdT0YWaQhow5eeFneIhxqkUPYw8y5wMEn7KWWI/7280DfunzccEkDIi
FKxOHfoPbx1TmaBS5r3PcSh9SZWPtiigWipw4VMsVEVSU+sIwPgNolW3WqW9fz6F
/1aRCT43cEqOB0dy2pSCS+0/zGi1RPHJRIPFaUV6o3SEZDtbxiJSEEHgO5/IZJ8a
N0SZTjCdLAJbk0COP+Ja/ISb4IjNqtCi7bB7zAqMTw9malhrJ3+n/qbMuNkfynSs
0AGykcoHov/pSZgUoFIRck54+soC0s5pdVED5P/b6WAFr9obC5R/akFF2NU0EAm5
yEl6q8rX3ZBeB5mNqMOnuBLePOn6RMTiylO54/VLiajXhXDn0MV9paYIbqTCA4fr
m38ifAD/Ctym8n8ar34KUkqCZOZt586wIoiqymCC3CwVeteAQrWqiYyAtOegR3+V
s0hSzg2PFUqfkLtq9JR89IhNhuzFdZqFbSVM/qEhDNTplRagEDJ1jppoyKQv4frO
0ZlvV1YJ3mF4AmVc7pqhiq6ecKcH+IJOGxvrD24sKaZWPYtZRWLVN2rhDlrYOfTZ
aARki5Lo10I/MiHNd3iXfcTRyHCWK05msO8WJZa9OLkFVVF7LsdlG13eAWzwn9RJ
RF87pmjs49ep70jBLWqalM8CyFjzx6dTq1iSYxaqLdLKg+QZXxk3UluR6Um1Ly84
txSi0M+0vohaW9uX5LVilBOkyPdGd2y+DRaimcqvk4Rhy4WCX0cLOr40ZQ7OLkAP
tSm2djuq+doDhK6o55NL4bxJzT/VIgg0VZ8WkSaGYEf7koOnpGjFNrv/0lt94YzY
Pv4UmLVbDXC+g1f6+PhDv+RvFP+1zm/OBLoJdFxzghqRmwzO9nbFvjX3YqDnzZrs
uAVeC1+otjW0eS8MxAA/r+vHb54tZrzF9lqgJFVBWPwcuOkfpMgylW5GxVM9i6qK
/LVhq0UYV6JCBZrMdNuOvRB6Syy6ystjKUU9RV8bX8GosFlMO6tQtHXlLC2LWyeY
dUQrAX2RHcPHK0c+2MweLvHsavBKEQczNU6Ia8aD9CY1950st2TUpYEK4ewyjwsl
ihQxvmeqY/JmLkGqkPwZUuDQs+WYIL0u4hbUjjkZBdFZIhWdi8VGeYlopMVxVUcg
tThCfnUFCP1z2I4x32YZZX37vihr1Vd1kcgUz4PygQK1Incf3wvahCCDRTPD8doU
nQcwYZwc2jKrmM+28k4WOM+x9mWsRk8fSxnogEfYaxbYz2mPibjtbMTBVv2mHCbC
H3tqCgDNLopPm5FYBMthUwJMf9P7ZJtLz1LoT1HdaD13G41QabasDaX3UBKmCl0l
IERNkeyOtYqOYEqRMrdAujet8djG+ENbcVnAK10DSw5zNnXObPhuHWGbU1BNRLxJ
/v9jtPfccGFVoeJURNpggz2rQFHQ245cdYNPf6WN+UKGmgBdlr0Vr+I51bF6YDc6
vFb5XKcSkiHCUoALNzyZRTDqpryzR+CjEQf6HTK8xIen5fpbXGERQNdvGjGJwiF4
VSv+7LzTL9LYdpfk6OAUvlskfVo6f1UALjcTX3k52iE6TpfYF83RfQ0M7uTQOUJK
PjD8XNUZoFARwTm+rIuMSrJJGiIuSjeoVI4zq1+Hcmp8E401nK3qg/4i3CZWYVpK
AvsTDinhgkC8/UAR54nNdYaLWDkPi58Se3gX5ORqEs/TqJ/oaQ2gy7tkCRAXAmnS
6NYdfbl3tZCPMMo1qtC73S3cIjXYLkOHakbfB7nnvGeVKBncf9xvxeTsSYMr9Z5f
QDvsJHtPriOke5GLmthp4z6NQ4A4129KbgRfxQys+4+20lw6WREcLhmcQPWYyLvq
nl+kbsUcSh52XEt2it7iTsHGKSvr+flKWmdzJbrx+gJqbgUXrUJt4e9ULuHUh2sO
MeIG0I9l/X0CcTRez8XffDpW2FN4WxTivbe1XgcijZJZ6q1+KvTmCPvKvy0jVdbf
m7H2h1QC2QC3/tcgwbPlhiXmJeFZmj8YJIK+dkPP624xOQa+0j3t1AnspUxMshCH
XBaXd7x6hir2WQVbWSLtgU4/yE+GoLpd5dhsziAxQZBIsaPz4K/tAhYZSAQHSvkE
EUusOGSru2Of0Y/FtRHxesIYKUmjYE0jwVpL4Z5ApINNpDZ8vVYk/zP7CwXdb3sN
OVSioiT/ehf+dsaJa+LyKmhkatmRyIgnI7WbqiVMY9zN7TqPqbjvIRO8T4qfwbts
A7n0knwPA35fQFksfvim5099NHDpFXLIqkTdtRNUcN8KQHGQ539MuL4GrOYloUUK
UkCvvw7IXUuXiq0r+E93yGSEho6aaaAApWX8zsCjJcovBgpEnQlmtgadrWUwrB1f
BSEGy9FLowO9uQ9ovUvQ69ukV/jLwnGoHnyvcoIxuivP5GfS/cSI8HpxNKRhnpem
D0AwvSkxXs36fSVc4Ypc7nbEog1LT73XBmThL6ISUeMhBwHXi48cJk0Uml/fjbqJ
LBfB4gAdvv77H2B/bgyr+LpUTC8WaK6/yUEGNFyey7x2zYfWr/SCYZn9/x18l4lE
EvFmGG8Wwd26gEkAyw6LsVyI77BzXn2FiqafDvEILXFy7WouRetrb5hcIbFXiNZW
iMJBvl6txKOwIT/wulgcJ1V0+ibXL5qoGaoeJWH65rWgsqKdOpybOlf8yxW0w6/H
T5QGcZB9nxQnD7cTjXt3OEH4n+dzFrLsbKQQCM2RjkvhZ50P1Ax4iC9S88be91Rc
XD69HwgMUNCSfYBgUzHXAz0F61fBs2yUeKShdlY0WTTCjD9Zg2LMtBSNWTeGmmB6
gqh7fTgl+jJ7WlK+/U+fTp5pTY2l4MkMovzEll6Y7eZa12sxL0Q+uxR40Gay9Gq4
H7RzN+b0Yzg9G227/BHa+zksou0yziTmQhQiv/XbIi4/hmvRF88RsEBvujVc6CkX
QTpjUf5Zejl7pOqqFFup6HdPCaopryCXpUMziq1OSJVph84xNNG2IY0r0DDEgWNi
m+m0jqtDRwn2WmBQymPS1MpPL1p9ibszmNwxQOhXFyORwTRbgrkvy9K9myXiHALE
H8RrHNzakt8dYfN2Cy6GmslrvtEThDxK6Zn0vLsTIju4NHIs0Nb+jO8PJag7fD2E
9Z+ysPqhmDe/diaALvOjmr+8aFKQXAkMiOixiYA43yIuV/7e6qIuxnzMjxJNoqiY
FirPcN1MeA4oI47exS3SLsba1e0ZNY1Uj3x66+6+X/+Z428DL2OYm6NnNTZFcehP
zyEBDGzMCfnAfXswNniXrzqSjivvl4xjJVYZ7NvUYV7eGodT5PLaIkomoOqiKBEO
4eC9YWhTxqL2AwPLzTDwq0qqd9xt4ZDLbgG1AosXrffIWxoXug21J6KkIDrXzJXM
SbDpLqyfcFVnNWIN5fmPnD78W2q7Eyo9ewRHw8wLXNNL6ipJy26JFkCxgXog1gjd
c0V75BdBCAuvH/aLOOZBEebZaz0FHfqbRwh6ZIGesuNQsRbunchpKbs7EATMKGmx
wryJoGuucf92wYsgUTgmNDEl24iReU7mbHyaZ/Ak/b+0VS/0uTP/idFEFS4xSQKE
QEOF9cx9catSLjMW3w62jTUEe5vCWX9wNky/AgUCnl9rf71reGGGZxAP+VJ2qtBK
86gdc7nGL5lKvp78p0V3XAVK/y8qXxlaAw+ZF7DxLJpQ3sU4vUKzVZm/SO+lkDZV
26l50nibznnV8CT2Xyo/1uSDbnNylzBuzu306+E7Z2sAXkJYf3KmKn7+DFJFpeeT
IzI5hN1694AgO8sdGdBrY8Y1oFiVM+Nb19CwUDz5QCRopTKSl9VH69+vCq2fJ8dA
Qwv0NDczA0rjmftar5e9YWjzY8RfW3PWAeSzq/1T0PnUOFLVA7EuCXxpl2Qq8cmA
K08LmiQoAe3z36QzCBVRp67WpnLDcDiLDRR6V6d+i5c5lFIz3eQwPO0P6WVBeWm8
1L9yzPx3/LvDTR0TridVWVz9EqHRrAJg3Pu6+YZPf2tig+B9uHr3XnnAJN6eXUpz
hDHJQ9SlbrfdioiknqsPeDy2C8bgNUBxzkty+P4BVX4W3E1/NxONDn0ErVXWtmym
eJGEbTZ1U4KxeAYnT6nTtokS4l1KCVAYhKMA1vXvr3bwLGfPC0m9eZpuZhuaHCU1
AgbcYSPx8/YPzcsXToXiymUx8ZrjZJC6s6rTGhy2Wwh8Ahca+fjry9meAxzAqzVA
3uJubN1ELpREjCtCwOFXfnAQE5RlKU9Q4eKv3iBxsa9cEG9S5CnSbkXDfRW9u6bG
Qofg/yYDkqNSViTNwmbODJAXYN4ZTIwYOZ9vxHdPr95CHpOWAlr+cMg8CjrJ9mWk
H7HisTOvSGyifjq+5ENiu2wW4/OyPB3KWsQ2lioEJQjHsmkrLIcfokp5fj3jgo9j
vqWAusQEGB82TSiNGwnllVcn+w+ml6FN5MH/p1T7b13y888Vicu7ShyfrYn62o4Z
zOTWLoV1i1ojtozG5O+1dDdAyD1P1ukfWdspXEVMoTOghDAmsyjuw4qouFl+Yqwn
C2syGufMJsBkAaNHRaNtzn9jIcVXkXb1+9e6/WQeve0frdjliujpI5QhUCxezQ5w
DAMnsOQsVpWhu98RZipSgWpRKbgDT4ettfNhcxR/TldIOSLocUNyN8XHeGq8g1yV
9ucOED+F3Zo2nNR700VrQoxYLDWen+a4q39xjvXa3IP3r9azgPj80g7oJd9hlYaa
Vfqj8Y9ys+k5lPFOJ9tppIvHFm7Qal9IglVObvagt0O0wqsPibL/vU8Y44Diz/QQ
e3nODnUXaQNd0rmaWG1iThdFUTiOSZuhA15I+edv4bGZFjV6UocoLO7xigsx4iUb
2BVNsTmesGf2pPlxnkZITEuRv/0k66P+gbuYSv5EfukBl3tPwZEkiwAwXS6gqXzd
BiBB1nEZvGvyqxxtBqfwX/Cinla20a/jbalEIs7EtFdkoJTQgeLeXBOeUO9xsMQJ
S/LnSZPquFjea/l32GnkC29YwB5d2zsk8OeOQn41oBrb5pGoSqi1yWjyfgm4+wUH
y77WPcopEEuhiy78S9W6zRXTP/Vxf7HGieggltPwNKMOPBBHplrbTSIMl9vrX0wp
PKz8ZL2AzhkPSVuM1+AobUgxCwNIiD/oNqgOi2dnLaf1Kr8IfW0IsLfqdFWD5SvC
RFK2gyI1UWngqo3yp6m/wN640OZFmda/knrzd8DISkH5rXcqeQ2Q9diCADXQdN6/
Mn+9xEmY6TG2E5pcBz7rOJKgneAe2lmkIc5jyTTYvMxvJOb3bg/j+7RsCIFT9myp
v6v0TfLh1RAZKmoH/vImlBS7jKo9SnZHhOgejsQ4hDQLaAHexHjUGf88I4vqxVrG
FcpgzrG5mIrFiW/GBpGKZAKZOm+PPn7SLMWISOM0YPiGjLcDJk7UXGptEs4Uk6lf
DQy3BtUPgcvNXPJMA6oCwZuCZqp7z7VN/c61vt0LNuAJjrXSZWoK57eMsjMv2S6P
8TiHfSxY4I7bSvyL4GI/cxLX1P6xscP6xkFBa9OZzDslBxT+TK8tlfTRw2FxkKb0
VWKJgxw9WfYmb/VY11EC5KYDyrlNutgZbB/SXkM+chBUPoIQ96TbQNWHDD74vOoo
e4/kOY6IOjUQIJCPsAVMdgVGahJ0KBGzZwpKJdfkSL11aP3KKY1KZqSwcGlZWQjl
rfppXgQ4yYyOH64l9nbTP6D156mwUAdtabvNPvp4SRQVGGPf+enx87XZ2ROcIFKu
LGlrCMzAz3PqmpVfvHqz5Wo9GOvK1IEtYw/w/khVARvvVHcHPZB/5jlS5BQjZj62
ZPEL6xrl9fGm5O7WpixcqRttp07Tl2hsGVaxyQ4kVAXeRJEmiUGc3wkb9FTf7ymq
TK7QkgRdNlYvgIGwdId2fZpumPj0IIDC2Wf1XDn2Xc6KmcxLKcwFEb4gowNPmI/E
PFUOmJhc0y0lh7XNrPouVeBHelKaXw6gkdOPZjRKdHIOK4TlTnKnUg5CHbdV9I2E
5OE92AFyYmvA212wCNe31HDSczkq6aTGCVrjcYRXCcaQDYiI0WVCMHpvEYPhnpzw
bv0y01s3CFBvLKbteMBnwSblK/Ef1wHVqSVjcQDCxS48f0oJGLokC2XkELbl7vzx
gUQHgNG3BaBpMZV440dba9w+jgY3jQnmgL5eo9VIaRr25USr0KKWdPwhzawfnGfQ
lfbuxm+oN/nTilDP1wl+yz1/Nv0/C4yEuvxY2sjRcU51MPPLMmKSLLcfU2XYi0rF
9u3JLR62AEqqfwdwHbWF1jhp2jewME31f8L1Im6XRUSpSnLz5tVxqXed1Cn1w7aA
n7Mhzvg6e2Ql6qWajNTnY91ZpUpBM4Kn7OHBvJs5vLpEHdclffZzvS2SHyHMzKpR
5gzr09sVQZV9mVgYdW+S9a2+8zCVEJCVcfZMaF8v/XZ6on9F12zjfyZAYSrBp1To
kG6scmKKvjg9fwcPxkc8dosmDZ+rj9MKZiuiJkzUl93Ckn4rHZpz709Co8IRxHiA
Rzj3U/rglhlFwXkv37ZiRhVbeyRjysBPNycJRtLKjfYC42BFGSCa9OiElKUbbpRX
pupNd9uxmE9h4WxN62In2LiuMTUiIqyYoqgb+4hUzGCe+EGx/oGgRkCvbxEjvDqq
o4fXABocn+mrgnCGh/9QNRRZBkQR5Y2wmZMLTBiQHiYU51hJqQxpVjnMAhRhTm7X
MMTwgi9EjqLLTNs9bDVtGlq30X4SsuMCr5vTy+5bjiXv6S+2TdluTE7LJQ/KCt4J
qRkOXJ/Sn75rTuoD73j5J7KWWuDM+ojKed9XDY3x+UFRRhNLK2Ptxn/gzK3xaJTW
bQpkP3JnBsRwPkNqSPV7OcETNPDAHS3fTBfOxpnExvHFwgqytI/+3TI5D+Hp1N1w
JnZIDaOLsHi2bFXo8av/kiBzDrR2AKszHf/Vqko9lyLalxMiDvBahMuVHxfsHzLq
80ZvwlIIfTpOCjqXTY2Uk6FdlnD8i3KcJUYu0/PWIhh152SWDD650kJdsjqbCoh5
wasTR4eTvs11A5FoBow80D4Y/YhtzCYnMUKAzl6durJbTpd9TyQDh/qgJaA88se0
0MSwR6yc6Ir/i3vzwMKKy+MiZ/Jt5pEPBqwyun2qBI7rD03tg7enJ1JfsKKzanXX
Z3SQpoJnknkL1DAsYwZqzHq4lO8y2Kd2MW503vyTK/hOQO5V4dEDWiBykfJYH7pi
7ibvAXbnwikqP0SBrdceKAr1ugs9YKQJO337qUhN5U8oduKYqZwBaEecK7Sa78cz
EgmoJruxdKD/7GlAMkglZGXQsu1zN2yup9JhLBpY2elyMYKX8vql//egWMSkatVA
jaPOE0VjxkBObsik8CxbilHKThz5922DcvwIJoZJDcQ6OY2pdAEFDWZq+cpfeG8Y
v10fN+29JK1YfKbRYkInlxFam9zjjBtSeHoc8sMNYK7uOBj8iKa2V4fApgKd94sl
a2daMPglDX4oNtCFvkCjteyDDwKdDXvPkoVRdlt+SPBcPN4G/JG75667WfGOnRTh
3sTuuxOYEaUlsThcQklfq+oxQ0WcY6aeyr/wDU7m8zPUX1pCGDMxHogksSuFdYco
WzYsegZ9X0At+QcjJCRj0eik1vxusDfHPXGqNQyI5HAxGa2iu+9QxUbeDFvo0I+Z
RMDZj6zA8YjnbLjRbcuDlR/6pdWwtkMGQhRSGmug9ma77QCl+tIjKX11jOZ5YRSO
nx4RxyWC1iL0718r6HbuCNV5SzRqYBKAM7Y8yB6rf6psLA/Pr5NOoINH5PN0dUx6
5yXBuiBkifTTSIammjqwvyMl75e9bQmwXxq2SSVVsNzGna7Nt1HLu4tJGESUsnNx
PxeiJ98q1bDa+ed4d72Awi3Uz8eH76kqGmZ8qt9zV0aYSLvl1Y0ZqF25EjD+oNqA
7SNI7hVxI0d+juaA5Hw7mKan8Wi11gykQVIGr/dTnuaxTQXad1sURF0qc15JXPRu
tDatY258X5F0Kj14BbBF+WHVpua+vqor+ULPlO/SUSsMoSq0lAZtFCIHwixjBhMC
sCG6ojZapoGsX+r1lc15zdkcu/ze1D5XYd4IO418LLBMzZfC4Q1L9SNmY6YaekXq
9KCeb36LR7b8F00jMcQq4mZGZg9+fPo+qGk1jVq/RXd5P6Fb4/Ac1Hd/xS/ycjxH
KcRczJ7DtnvrkiXYunUZOEqh3z0nepKc2B2SI2iBdE2bzdnan+HCIJhazMaQ8Faz
NeMiFMnm8Z2qPbvROYcbqQtvQzftDrKVOMHdu83nzpSaPm8SQyu9NoWrCYUNdmCY
0OfOMcKzFF3iynhyZYKfdBP1ckT3MJGnN6hXvWOI8NbPC9u2RIOgdCQyN1bqrSgC
PpwSI8HHC6+5OUaoq3YLmv7prdBGplz5Q4EAlhx3Wahn1N+Bk8kYoxavB6KLs+j+
yb0xTaPstXGsUgzJUk8XK1/fk8hVUwOY3objvPtMnpwChUd0Rx8prO7tOQjMXUh8
/jvMfJi1ZPk6y/+yxtXA1SxE4dFp65PTg3mj7IXKbRsHnQ1Fn5EADPZ47cHiJtFb
4tPKcG+DYUd4Ba4vVQOR6+mEKdQZVO/hZDp+EBFFXvoyYyq9qtlrvth5jUjDXDdw
Bbkkzdw6OVBJH4TQrZreK/rQEoFw4NwReWnvcCYPcr6woCN3/c7ML0H7KPqnCvKw
LbN9xwSpBIZ8PIPJljGpMpsmZ1+2BFHLZ8hpFCoF1ka7XiaXOekGX9RGVYOYe+Hx
FUX65aB5yYX0PLQ6Dj58WXBVFJ7grMTGYeTCiETDkXMfd3+GOXpJQDDf/4hjNUl4
w6TYZqo/jXo/Xpncs7Fii20tQ8vTUOUIRgEboeoTuO1lkdJ4jYgvlw+qZZmlmUa1
kDJCOwRCEiV6f0ZDvKOcGvE1R6PABveJYp2SVVUMnxJ0tJR955AkAy+tCc8eUwV2
oJhtoO3SAZdLK10bK5BfwmaFUKjZ6P2cHxrRtJtzJBZk5TE7054Ztb+fQsvlTxBU
2LKmhA73ZybuwociDUP/x13P4gODmts6pD4UpZl902fObvGMnwGwup0JgRtv+sPC
lR0ciId6mARKttnTwmwyvhByCBJwyELx81LMXG9ordf6vpfugiYlu0NnZyqNwmuY
eJeMit1k0GaAH7k4k2B8JZOydTckXkTeWElt6XOt0HLxEQ6XMIuqutOdMcOOp4Rf
udOGMJbFDs+UMKCFJebr/1f+dsbUav/prL6m2uW9EqV3BqQTK9rdEpttOl/OJhy5
Wkon97evIuHOKPJGizBQtcYQl2mb0K3lBZWTSCiL2aC9lv7XQBfU7umtGcKzshWl
nWePpskJtHaWDvLlhmWuZ5PNhKWgxv49WKqPZbC5SSgQirHpzJrBdBJg5gIag+Sc
N3GAH/LqbUw2P+PkMaRzWHHdfHxpbOPX1iKXPtowRjxre1QHqsKRWSgNQCRq4dE8
zD0pJKq8QPjoUlbOJFNSHIiwiH3dv00GvBufEr4afS03WeRrDkfFoUdscG/Kb2Yh
LCC0MRX7wW8jlqqcqzagIl3wuiKsng5nTZEcAeu2Wlwo7MCqB+ouefKSm3A5gZ33
JvaM1hIibUzEcPqtaRAVXy0Sy8s71SNpMUA4MAXTNdwZ64uRDuJ991hla6auZSl0
mv3EJsZufUAmiOrRntVPgVLB8NWHn38zSd38EOBA1q43oovg24g7wDyDADh6Lvg8
y3Sh1YFJ6IHoMAL6iotByJS7DxAILnGhUw4Pr05pW53PlhOv7vLzH40P5NJRkSUl
Rr4oZCiD4wsyENFkAV11uNu4PAFRP3LtW3fsgjZ1o0wmDpEs8WbkkNvV84XaYxV7
tQXyR4o/CDtiz+rrbjBxBNWbBTe5Kj/e/BxX/knSC01oMPVTOOb9dn/l9ch36+Y+
SciGuqOahdObQ7HUY+35v+1Qp+ncvDyUsEw7eAsA9ZqIVzRMLQSpRTJK6pu0Za/1
cTFBuk88FLCIEgDTRmcetCV1ksLuF6zmGtO8irUST1+ZAPldTHUOD8iMfZmjq3Cd
BZf1h9ZqqwMnV19w97nbrMbspzRZXYIHj0cZgty6DSxtJh2Dk8/XIkGSmFvRWdl/
s4U0VMM/CWWp5wxaF94P1hx368qT7ZordKMzR5HOGfyxsptXhy9MGQ5wB5KM8jTP
HlT+44xFlj6xLIo1TgMTCNyPPRUY5RwKYSCCBLe70BJPjYLSjgij35mAEM7Vievi
AtSVYfdQtjoIucJUF9jbDAb0coKCCrMzRQQOUzkkAtavxu2oeIJQLDeThBlPZZrV
JrBo5mPuM/OwD1MDNK/Wgh36JIg5n6Clul8scwWuo+bD2+jF/v4a/ZZd6YCwefRM
dMx1+XjmGKI9wmteKLB4ziirtZNpWKHNNPcWyj/swDTH2xMqK52CNdjL2Cjwa2+N
3Y01zmVBLq5xHLNEmyMLNgXVwMTUEXhqqrVpyDBbelz8Mc7WsgsyEVlGg5jShrnM
eyDGo0ynvvXidHsjc8N9zZ1/Q8nvLv8nsKg9rJ9LgG6czZFvGAe44ScEaASMtNvE
ERzWl8M52c4yfniLm/bcqDyYUucxAJ6mXnLgtWX0YArrLS1d1KPngGgdSH0VGHl7
sMbTtFEh912iEGmtuIMTXLFO6Gb8Sfu7i//d00HdLDElwjCvIfO5KFIZlBRPWa5J
wILf+f72tI98caSZuWpCKcRlYh0Lux+hseQ6H/aQaQ/hOq4k75gMvLo91JNcSq/4
0FLrRfvNrM481isoANPmDxxeZE5Bk2v9qIPobWOZYmg5dM9T0pdqKn/WqiUfS6RL
aavA76FSytC3U64tNj7/Vh5hGbcTC2wqyl+xAHUpVIAmUKWHrRn+b9JE4sO0Hrbs
UVuJplu6XHreFGdgoq/XIbdOS71c7oArFxnIXArG/KqQOisqWD1UqnzgVEDiDBFE
ppwqgXHmtQX0zq6oIx9qgL50rVoqvCezpOF/bgjn9iBq5XYrIjQOvmP2/kqbm7FH
Jd0fFkEGL56Gl60ghNaxjdSq4TU2QR5WdMbHjlxxUnns56gFcpVStijcM2zioFgH
5rZO4gPtCzbxxZ1eo3JAPX3hSXw4yKr5F5J8k94nyOcaCdOV3rJvMmlE1fsJkx2b
d9FxG4GYcjbIB2ybOXZFgSDfXfCIWRGLL2EDRdAGUK5m/hN2cwSsYCrsFX5fcmto
33dDL0/aC1ut9kGZJHsQ0exx5RctakW+RxLosemKGnniIHggNo6JRX786GbqdXdF
PSYeuPw6eZrOZNNym2C4Sg8qh72zxsv44CNi4iRYOIv30YRI0fkDC9hXAJ3VqwIN
v32+oJD7d3gPMnWL2b3I41RJKBstHe8ORIUH90sAxJC8qnIm+k/+7xIc2Ixkjlx+
JIgD1req7hcSci8vEVFVHL1MvilVERNRrOlvDaLjuVr90EjRkUGihcwmfNr6zPcK
y/Ar+4dAyq5Ed/48G8L+UYEPhYYkVZubwTsX4pkgINfBkBmTVwa2z4N0MYCvCf2j
g71s2MlDCvnuLDt1kgAQA2FKgEXPplnMcF4oux0L5+is5WM0FkOxOTicsdJWkggE
keJa0MFWOM9hNdcsmBnYITOx7KpdG+5RzkC+SL3zmknLDArjSt4Uwd6AElkSWwP0
CUUAd5uBxoHwN4sZQBbU8wDJE2kDud6BA4Hw+/nm68sgIS7s9QM6QMMb/z1He8N+
qJAaEpExtM1BhmN64H6wA6F9eDwxhpP+4GTM8VvIUeIWQ7z09cRlwMZCcbXOdQeJ
qDIIthx1r3JQYbLW91cjqwgaZotX4iU5c/444LZ83j6y40fMbuf33Pnsl5J20X0n
pbjOIF5OaNVlUYeKjpukt3xiQqBvaNtMwkiXFijySl/z4vblLGBeXIMcwDNvJze1
IY36EmXPlDckq8pk6ndNouugdy+SskeLm9IpvPkj3kTKcVnaBU0lghh1MzYG0UkO
khe5IGrxCYvsXRuRDobibTgzrHUX1BazhAzV9dKl5GEl2xoYpNiS2xkdBWYmKO8C
hkFPYQ+p9N2s5m/DM0SLtcBFzDOJoc8YK92ZB5HrWMFihv9v6VxyN5K+QQh6TlzN
f25wFxxF8Tdzqq8+z3mGXXWOHZ09a6n1fPF7MkhN+7FtFBk6qjZUhUHlMlBluzxb
r0d8ERT5L7z1A/eOSzfnOk39uqjHb6HF3DLd9yGaYi9uKFiPaiFYYFnb7+DpV5ka
A6/C9ojrPdjQLAD/7eLQURqCw/0oOP0qljMhVGOmStQrdd8xjSjNMznYHf4VgnET
dnKrUiKr+/PzWferB9pgJ3rTK2zE5mW/Bzs7Rd1wfAwLjPE8jsUqQF4oC9jYnzc+
I8tMot5wCyPoFnY4ACdo/62USMalp10bpVaC0rKNUjXcuxR1s6OmcQU2TE1Q7Luv
f9ylLYFhuwSbEI7f5w2xjnRLMfVjAvQ6YinO+uN+452rhae8KJ9qMZe7QFVAlSPj
OUZvYHGcHhKl6RoMuxF0O5bB1/ndsWUa0B0tRj8R3vFjWq6ze6K1QplGrHmDeNrN
REmFMGbfCOBoUCPcFzBSZlC1IoevkX7dUvDmpY0G6+Z0BaJWM7yqTOTmdIdH34AV
NmEKi9PwvMeY5sYZ9voygqGq+P9seDoAJtn8m/9o5i3HXV+iuXT7PaYt83DZS6gk
ytYPXtOjNA+4b0jVaFDUK+Dvg7fTAuEKMPGWxKl4dVkI14M68b2sdk7W8tVyPw7P
fz4cryy0q7ui3MDzbcYiN0ChUnCQeUZyK1jp2ZbxIqQjBbxjVUtBpgRK3eOkVB9G
vEtbZ2k9gnMhS9XuROXTuCZdzBryXwHG035kjbx4UZpWigzX7tTMSl2GrzsuM9AR
UoqAnKQwqhY85DPW+5h75dq6cHTRO2z/g+Obc2JdKI8Otl4rhnqpOw124WeKgYTX
f/TDbLYPmKskW4aetDaqKft6YqBqwhghCX/qc7qNI3ma7guNTdsGP8NBVBpbg+d8
1tbYG/+xY4EKXrpR9GfffIJ1G37VPwn6McU/uzC84xRf6gHano0Ajv/Op4sMoqId
/TrwMyELfb0850dbtEOO/xpAA4OIb+olRxVcE07pzCYi8qV7QXpz54/e59Ckhj8q
FjPhGqPoJKRGXksQVuvxfY4eyVzDG7UhZVZghboMK5I8ZqX4cbD76EWjInwjk/l8
gYKCanAxY5pBmgJtpryHySGyj5hn6HoHoTGiwb5RJ29lcQKsRSdJIjDWGX4V7sfd
rKWD93kvD22IIyFgokLu4aFtWWWCAKtyTvCxlOy4OFKR9jk90CqNuO1wViMGOcL5
`pragma protect end_protected
