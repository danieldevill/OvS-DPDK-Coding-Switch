// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rPrpCR/z+tiTxIIGQKAnObzltUMdFyD05un+MVUgM/ddOQkoVMghnVbrtqSdekGC
wLYNgMYjPUtgN2fQyhKznT4Y/6b+vj1gsPb3i3eVKe3qvenp/zE8JYl9NXxN8sZS
VmlAlKXRyD6IQez4MjyPWMAipEodSVBcUtF5vTwlL9U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27680)
MBzmNoUMOHpFKN5DLjRYOzri7uUXUViLikD0nqZ5b4Ycg7Kcm/8L6MP0sdMB8bGj
zfTu7u29I5VJxW66S/9n+GGIYnGOYoRtTFAj+oH3nBw2Uv2mIJcCR6ogTCN95Phg
L+8o+7i5bzhlCb6xju+tKLCk3hYioeDccb0h+fvuPsFMIe3rtGWvRZLhaNyeBCgw
h3qcQAvXiQ3qN342jwjAqUADzq2+4D8ZPn8jFNOEX9Dmidu+a+ruRfdL5E3Opxar
spwu6ybU/4zZwolcizZl77ShUWCQx0X2YoZdq88JNiDo7F1TUK2U/HXZl96Z0jPM
hPyXV5S++ZN8krzMXn1mTXsF0pM4F1m9BrudmdfxHCCyU5AHaCXsoq9Gl2mqPZlH
4LpFILBBVqpU2j40I0yhOeTWOotlQweVHawhilB0+VSv4cm5fl9NfWXcC15WiNy9
8DuPe2wkKXEfmL+3omlvkX4jLTAXrzoHKOTt7Y8n4IX2Px6YUy7wfz+vGQ8vBuPE
03a5SKP+VMWy3oIkqPhusa4KLIHXdYZmSfflskoUCzs6IEXcsCCi2aCp2Hwcw+L7
OZQVnnme4Vp7NKgYpe5XzTCfnHXsZQG52JqV8xu4TwV563PVVGn12viT9sIM5Pvt
PbKVHnj61r0sA5N7mJZgabBKliWcrAs1YIByxToDycgHCiSV0SajKPFucKJ4Psn+
/z9hSh1MTZ+nPhrK5+u8Q4+nO0UB5F6eCgCUGVl7nEJ+aYZq4ftBODZmz+iT3gBh
Nt8/aLfoodmOfiNDxLBbpDAtO9zffm200BYUfSn0Wmnxxru1mQgq2KYvnGFUydkM
MP1N2JS4XJSsQdu1WihQSYMCKFY/+Map2YNC+yfJW9r9nVHtyPNZRYLPbiYDZjkd
KVQ1kSBCxqB8PkfU1zxg1fFrHVbddJ/uMY4F49a6M1EqvENxQVNIviWYUh4AxbEu
t0EzNjGI3pr3gS9cyyuLKWzDj5v0rZ5dIF12Kq1FUr/XuU1qpb/E2DraDNryTc3X
1/tGlAdv796LZ6owpUDV33nHwAV830/3lWuxQRdaBy5Gf8zgxgofaUUkvheSN/ax
Bs0S5iOHRpuOIKgaZiGTvLuvKRzYWKrlcUb/AYPWwSUuxGxMhKHbDdCL3RhCvoPm
CLXSOL/yYPmQot1M3fl7jehv8RV+9/Xlmpc28sVRn2Dc0EJmhAu0pkrA/0hUKY7A
92aLOqJ+SNoIzVA4jPbpyapPMsEXGlNwg6GYuFmdwO3Fp9Ls3AURZbMCxlVjD6Yp
b+cRNXuH1nj0XWumFJ4WdRMXNz4AsMxx+2Sm2hP87B+8Q9DhAwudLH3bSl/6z2F9
EL3X/eqEZoDuqhWTV721nbSwXA+9cvLqx3oVQe3uQ4toJd6qIBN+kvrkykhSp8N6
YGn9NbNnztQX73/X8/M5XC7Q5womi64qT3l3UZM1+nW3m9VWUNQmUyuYCmBRpgdK
Dl+YE36H7G0Mv+g9no9mthi7Ll9vmLeQieUqHLLySLJqPPaRbzE1b0ETePuBcpr0
7YCdA4O0boSFfE1NqWvG5Yt0U1WNwx0VxdloUDIm25rr7UU2kqrPRglhTsp/SZ7u
3cMFmqnwrElYr0sxqpJJPIMaxW+xj7vmvOxwJuXtABu6KEbnyiN7ZsYQlJwGsRJC
OneQBkJPEsIzahh5ez+E+qUP95szQT+r51ipFZ7tlH57mY8+F5J0xPkuMVj71wHy
4QYOFu2B1tl4f8HLZqaRYVfhzFHuIdcS5ab4UaEn/sD4kgd1hg341VcePqRwH8MS
WUNRgY5QK7XWmbo9B6wgeleEDNGHSOA0FXAZsLiQWobzI1PFlDo7Xb4izyw/HUAW
fMpWrywwolJneMGdp1t+tPNg8ZHL/rmPVgI5TviHgOhGB6i7VrZkYhLZZ2v3eWov
mz7x6NwNP8pjRWLpEwTe+YQFyGz4x1sD9VAbckRP8beMewKMqOHN7e0Y99ma6ToP
6uwIQzXdlev9ERfEaZNyHmc9SVAE60hZngul/E5/t36EjjeKKmfRRE2mFe8VqBcb
ksz7I3VgX7ThM2iY9v5wCrp64dByL+OPJfDuwUhvRk3LYrHSM3sld2ngG6PlsLMb
ntHGNifs8/5bmV7hpXPIdkXen/FIQu4JHtx1bzHDlRVAcYBW/c/R6zkCkfGexkrG
13L+PSXZ63pSIS7AF0ESguwl007kS14gLyv+mOZfcyTHqY6Zi3T/1uTxnkWQiB7H
gVRUK7pbDFQit2IBGEjK08BTUVrMvIBhhmlnz3JQZk4OsJhU++MRCVYNWeKvAbrg
frAngDwRHpfGcyHDmtlo0c8JjNoprgn+vlxrREYhUAyNjBOzdoGPaKmbcMFZzeaZ
T67LNotWFn4KHj7ZuAfV3MTmFxjyIULlUeLqTTQBv0SoTluGz5VZBAbcM9at18Fu
q/w+u7HtdrrBhr5rcQPzj5Jc07DY6Qe2rDEFQebZNwtrfB8RZNDS9F9JvZkq1a3h
TSqZRDZPykwT6tF7nt4fLByF/tdWof9ryDqh06rlPzKQHiuy7aztE1knsQWLg+2n
VZ8ECSrvMYhZdmXaNJ0qiR8+PfHKd5OEEMfvHiQ0SpRnjoGktSJ7PkpsIrxHX1Fv
j/1C6jYO0Ohq55xrN+mL/VicyXJhi51CbqL2SbVu1pYCrAXdAHJZKLW2Nqtpwj3u
jTy02msYnPX0fzWPWa4QEQaL9qQIiuY5e+WU0wgQOZMWBA339Vkygpv2YceF6HFL
fK6AmX/766KiIDJLBi7eEsPF91ZP7pUOum/aqoIvRZa+at+Dc9viV7QT76iA+0FI
oPFgI5R7lrw5abt0eovsvW4596UnENiyU7yV7h8ScdsMc70bX6FAyK4rddRsBfH2
hGFLx3fQpnE1nmT6cK7xJiGXGKIh+i3SBa6eeqmhvPx5U0yxGPiZp5NFElXuVkNm
fsCMCOm4O5zEzAub2KNo6OBQtl2iioHpnwqlULu5v9ss7wCYkGm6bwtInVgolNx7
+aCpxpIEUPb2AtasQ94P9mvXUvBEjBKHqfzRjWHaTrdxG2CALEEDtTAVgiVrXehe
vfQY0uS5p0+cRk96OW/8pQKR1GDm76uqQGV/4r1YoY1l8ceDHLiXx5OKIoJzeLAB
VoNZdmhRik237dtd3jVgcssSg4oiCKJ3YlEzHNkUlvdJEHLsbY3B4PgdT6T2In6V
UqkVrPzGcoyUBQcIWh7zB45Z9/XS0i3kqgyUTXE1m0CCnOPMm6KIYLu5w4bNi/Ey
4diHf0n9W3vhZOaCGXXErP2wVmbhoNZhj/A+tY0SljrLCeZYnIe8IuBX658Z8IOs
M6/eWTRoBvBPXC20ydFHLQ1RrNH+EUi4THA/Zexj/6GCm7LWfwJ+5tEcCqcoiQRi
IymCxEzvprEPJWwrqNQzLp4cRZ6l5DaUxGb5T6OMdJdMqvAmzdh25xNyaMzeE8/u
uoCDcFzQOccOPG3K4o0bWudXb4dN4DsLVAlyo97wdxEIKnBXF43q9QBZksNeucEz
HNFc3QySK63cKSoGwpBCvjtaxn/GdHqvZVW71lKS7Sb+mRpMtK7yIY34J65+TnNf
p2ajRkOES1nBWVCFnXNNXG100OgSxMgZ1U+KbBtbRNMCVV2S/5fCbc7tnNshdIvv
1BjCHhdBaMXhTuJXZBXInrua0MS6UglC47FO61dRv2zDz440crw6I2zEQYEl4psu
qGl/uSZV83hmqHbH7LPpITHFVbsevY6Zb8M7xcOeNedQ56hef3BfVZNk4xWt4u7q
q3XBtv7c1M8NNwDhA2TPj74NZMiWtFsCSHqsxutnTDelBPBklfkvWNnNt5L/2U3D
F9ptCY7yza61dwdbtDt1hN0GCr2He34HN+83Hw01D1DzTq5XwBgJMKEBRQSN47Gd
2jrNIpZpLqY2VnN1TaGegle2oZ0jPGCaRRJxfzpUgSWQ8dGporuYoqDaCA+yzulB
+Dv8ZTnyGLFZXjf6oRB+LlneST9nq7byjwFBdYq+Pkx0nnoEoWOJVAaytVmJzEBS
OQ5eXMB4EBadIdYopUbRqlAai/Ubkf6oXDxj9SbaLIXgr4f5c1QEvVBg9DYtS7ES
zSQEmfj+iuAk3HKbj5CSiwb6v9RALQRunFzTzPvWJTTONyrqmSlHUv1KDdzuQevf
uVKY9IGGylBGitx3vXb9vs/2+Fo6OfCWZv/H+HjVWKXO6YsmeepNBkSb+Xc6OV0x
hjaIi1bzospv4ztRDeqhJW6Q2S+KFW1xOzJU4PRvtXsxR3cIpOZmGAYS+BV2v05K
xXSaPI8Lt1BuaGiJyc97MvdCoEcO6x3TK+NPHmB613TEeMh/AewmjIew7l3iaJMH
9ZvjbRYOyuu5YjilgF7CuN8hKt9z1ElQM1h7e/L8QjApvOa66KgH0d4K40SDPrXk
lwktMlq3rU0Ebtb0ZTCoW9O8Rjc2BFXwznHSI7caO3p/VefQ+2Uo/elK/5iXBJCi
CDh8tgTNfdyt82aIwd3NNTEqtxi4koIiYtP9bmJroC9lT2/W39onaj0nMEPMOpJ0
wYYLOV8a89t240iAHB4yXuGukthDo0+nvj4g1sWpu9GcM81hNv2ZIZWJ/lJNpKz+
Q1Bi98rH68hizKoQFBMZCPGN/PqlKt/n/5JuEMr9Lfdw85nD+TmGkUT/QNP3g3zh
cy03Byd0sBhv3zqUYa3zwD/XBMFUMfhqmoYKW9MQA3YBVdSJLLbWMVWwa52vudds
CmIoh+LsIW2k4VCqmyMIylnXn7ZgifgFAcHmCDI3A2jZcJJXpollOQBTLQ8JlFgW
uAqxthV6kVjc85932Kzh+KJZzPnkrN7NT5M4kbNtshq+qckqiJzqWHot0BqcAQeu
0djRqN3C/IHkGR51RDd3chavGckPmW6dbiwq+N1dJiyVj+zIErgRfkOJe+jAOCvr
5/zsFWvesjgJxUbh5NBKGXXE7B3iEL4Wb6WCfy4+BPNN/MiYFaaDMhwZzEA5rWLy
8HEFJoI1LUY1T4frE2tFgz0Qe+F74GqWRPnqUMkcG5uLHi5U2C3GaFKA1rVTs9Bd
p6DapFAzcwQMdsJPR+Wq3PNCXYgXx83Gb08ozZrcLrBy67IM3ynenWnsX6Eq9Trh
7p16e/iTpoNAP3wBeGdxCQIpa7lKsjQ16Pc3gvSci8rm2XHYjgTzO/tWHGmZ+EP2
wNN3ZE1/WJmt2LWQ0tJoK4cu+zuaT354UxQ9Qp+ph0o++rC+B/ZDzjVPV2LsFSpo
dTDhVloZlZ5I2uDnsXolVr89LV6JKAnYAAL0KGR+KGzZwFjHjiT6s3lrJqppbqWn
JmMSb7GFSyzwikVBcW5zUbZKTXOU9xlpl+a5CGIZO+cf4NVZ5wib8OWC9SKdsLP5
WFos/Vf0TDiQPnY/o9jSc/i2nLAuCWIsf5NAnrjLHA7P+e/JBo8MKdbsCTWYcEBb
e2+LJMSYeIltzp8I+mASf1BRroLapk8romOkapJHfcg8kqNAA3MaDmx3Q51A2ecS
KiP4ltwtwZyPHfevrfHboMydW3DKpLkpqsDaWCVdJ3JSzJAqovTuMdQhYaC/Hz+c
FvEj23GbhgBHzZVxraXLtOCILcDgzbL3DQjs0IvOTDMx3Pr64mpAxi+f8+/zaUob
uiOr9VUvbQVKC+kZhq+bON9xns2OezXqcheotpkIWQfudADaz7lsZZVQUbpa2u5n
VC6QqMFT+NojNx2BHsZyEoQuAKEVLkSefRSBLXJimZ1jTxDV9w2CW8IUyjPGcfYl
pWBAcPgWd0JKJzBbXw4tDY6MY8h7+ABSuAfi22iA1gAy5aIy5fp8DPN+mC6qqf6K
ldr1eM8JUC4use1Y5NGVJd9Kq5V3m64LS/ojRc/wnL+2PBFBHyE7m7oeD7wgALu2
bNlbqDqMKFMm4piwI9AHLgRqo/5pd8FHFvlLI9Hw0y5Po9q3SfByNi1eHAiDWK8b
Wfjrh4Aw8GvH98a6CLwpqTVGf1OUMpwTYvZafiukeJtDEfTIv62ttfoVLJwlemM6
hv7U/2RVn5wDCuy34hSbiIXqGNWGRgJIU50aA6ogNlHUZf/PgpbnXwCNlYHylXD2
FzgUHSFY4yfdnnrELH77jB7JI8j17HvWP/yB9YH0RcfL8pSm+0GTmVurM2bfq1S2
Ngw8OFyxpLujw/bWMEkjKpie+wq33YD62CHkHmpIpxslLIdZh/yWGhnmNicDYYxZ
uaHIfCp5tCIS8Zc89SsHoo2SvXxgUHfAeJ7AW7YIUcRrhN5TMF4CLAfuv8briizD
6xvdaQk97tWZZGnur75eMrUSxgG+xE1YVks/B92lwe5GnMIcPBFBIT1GAewUaMYq
EcqVOACQIjdhByhMyOyFVQrz7U2JjX8oyCMUlUg0GfNeIT/Gx86wCZqsAQPkXVos
b80WvglfEPRsDRqEPjN2N4x+N3enD6dYRzsr5mzEU61rnWPiMSIa3UC8NwBujri/
IczRfpC6sNPFV5jgwlpjtDBVvo+7uP0WxJYcGTdhYjikrZfADc3pH5vEv27g/igw
V6CzFmySL/vN7sF6hCdxvsncD2pA7mI9srZgldQFy428Pz0OosMAae3ruRGbWNru
vz73j8rG71UGt6X9LfftszUDpBnVLSe4AxbJmUckh3jEyyKbiwTxK7djA7+dRHwQ
f8fStgjVcSS3f9++xaUlrSKV90qOAViyPeHPpXoHpyH/M1We5iEHpFX5bYc63zQ0
P5Gm8gUr/Bbzhk19bPzr4NWwI5QaV5gfqIwCHdcVh1WGw7ADz4g+rcYHNddeEg0R
VOfuG53tNy+U8/1punoJZeTKJoHNbncbqvgXcoDDfgQbu40fRDJUisUNiVOV6fnC
LiuQ2oKQLAtQ1f5/X0VQcE2sKjIWp5rEseRA5mNsRNvfeHdgaAyFPZMZ/dt8fotQ
T2SMWZ7KW/W6DFKvBTAAtfP2cV2KHmxJcgYeAg58w00fdcEUEUdZAU4kAUdhmzpA
Z8C/cenQtGM7qaGlIhERSVWnAndYtUJFrnhkLee/NYawzra5syu+kPKsBuoYy0XD
WHLxLIjYIesRxVfGYC3qVg1cS7aIw/et6LvJ8Ic8wuASAQbe45OJ3drNBD8ifaa2
1evVThKxrr9b05zpG/TFdktSuVNHFqx7HnYbqve+lJ0soDo0M6YBNTNIA6PuXMW4
8/kN2k1kEIpYJyt7bQ6odkiAf7P27YXQEUwEdgwfu7WvNSyHK+DmOc0SfvPJJd8j
uiRbyqmxDN8IW+wzp67if7apB5pHmO4GoITpN08kWoB3t/BXHnpgjaGThnaEsPkO
x6TYyyLUCq6mWHhnwS+tQQ+3/RO/tuEp2f5TG+swu+Q31A4l1CoofTHiW8KRAgux
MF/Kbkocl83iavdn1yRP3MxGt4KLc5m8CBAqmiAduSvBLJjwn8ByfY9quaTlcXVL
rGvSN9IjxaPAKmHGuIm5edowl68ioydMo1RGfxBvzBowXc0gEVlDeY7xoRTOEHnp
Ag9+SYGzZFHoqENOBPjpOAcuZ4UsrIRh+EI+A3ZrvU4YmzZcevoykJaqDvcN5qyx
ReGT7OFhRb1aVKHCl8yaZPg3teBrWlpPq6Vy5HZ0BQW5R45d1Y6kibZ4UXNQoALl
ZL6TQ0rliktzo3Sc86XsH7/DDZbgkaQTmW5fBNxHapw1t4EL2ULwUuQxD0lQCEej
iv99ns9BeNqBxX0cKas1SOLolZTHDIpgU/4IIlss1u07l+W1SuCuEk1Ky9uRrzmX
IXlAXsRfw7i3N5v6wXgK8oquDUFJ3E1ZuQjzxPaGKwjeAvU7mLMmEMbbz0nGKRYi
cZdM9RUYmP/FJoyf46LcjGHLDNWpTYJoiDhTVhnYTBp7wmrUbtOzZ/vH3Nfisn6Y
8vsaNZcqc/RZghQsLuuCpr2bEn2LCeIjnn668m+rJ8Q+YuGxCJUzWATvHnVhzzDI
jbGPVchtBGGVG4/LxI/2f5j+ssLOKZx/n9ozULl5ctTDTW8hnQcw7fjOKtV/I1tN
qFkOPU44GBvc/1v/ae8hE5xcXv84BlifPMZJlDAqYUjRoiAieyWzgLx40GSa+Obq
wvmhHFdURay6MjecY+i1lR1qAZCkDTttS1j9kOuCXYAZtg1UawGakEc3HHSoQAO8
6+gteQ0/vxuy/tPVhm0pojsi7ZTfOHar6xE7uC+7WaPVir83YrukOlLwpbzMpYhS
QKy+x1PO2hCS7ClQTU0KQVpaD5OxOjdKf5xikIJ7rlO6IulofS7Q2q0qqra6/c/H
40A/g7xFqwXZT2Jhq2TqjQYkFzHeUugsnlAnlNa3PwCidxJKV7bkqlt4zvt9wSFM
o+TqzfyE7HF+Q8OBrXz7IOCGHEoTCpEaxYgx37rKhIT/npofx6X8GxlUkrSUwSdk
wsunApbcLVD+Ov2TNflPkD0199xRm8pu2O7sOLaaIRwhkv34Btb6O+M0ZKEQRYlg
LawDR/oanHqeS51oncR2BA56SvM+y+atV+skeS7XLFjZooJrTwshpbHdSUIbO+A+
gV/LWWflSegpdgih8vluSgx5DnayJBoaAyt1PavRVmZt9RmTvjlj7fjWZw6ZuIAF
7JPIOFIQWQACJOpUiDv066pOLfMFDddLEV5KevcGaPvv7KbFne64qkKZOgzx17wF
bvj94jkuB1lpGJy86F0zkQekMHLmFMHZ0LV7njJsRjuBid+i0JWyhNnSLMzxJ5xb
xywnoVxKxU7otoLSt0K0Dp2/snrGJGJm3SFM6hbtzoUQAKhlAEmI8d74dXvur/7T
jlIUiVjcB7JuBvV14NjDcXjW5sirjGOiCmkYrMDlP4AC+lhRFK0AxvnwBl9gNLR1
+LAygZhF+5fThMI2KioKkmkY2oTasF+iWSodif9+uPSr2vvpDG3Flhrl1IJE/cVP
VRw+ssgPBJnaC+gzsAbqZ2+IUgNUjH+x7AvJS1/96tn89wqpgu027JRIhQw9Feep
5PvZgNcyQ2i/TLi/iwXUFIHWW7iMz2advQDzrT9QPhnP/BkN1ySzRhqOra25jJKe
LrcqVWxc7Zr2rtqUU2pvk4LiUlWLl/l0sTMmub90lygoYaJBI1wpCUk338EplM9M
pCTYeUkWxCYanBMK/vN8GWVUovOx1H5sRvSuj/Q2nv7r0x6QeUZmQdzdKhD0Is79
aq7o1WBrUqJ7BeXUZf4Z2OC6SJRiaGt7VqIAkC6gwAPCte2Hc8Ni8WLmE1X9acqQ
uKjCG6+tPV7NZYBBkGpB1AbFW1tXbB1gcphDx9y4buKzuK24+memV99s5io+du9A
DCn70RRDCpOdOYcUcxkJGy9Xs0q8BrHlPFxg3ixDlR4LEHIXtkZSD2oKYFa9fQQX
cZGPOm1DTJT6GjL/Fhz/EsQEtfwGjv8AilFK0agTjLa7XmSrPSVTDIQanGOnycc4
RaN2vF/rWfkGgQU4DQc6SSesjcQYts1i97aVp/C+NhHKv2375edaiKyyiJQ17+Zz
MI6YhCgMEdreeSeRZayrhBhDOLbuIdcJLsV910Rs//fjgL9dkojKpYmMpm5C2H/X
y/Ilz/d4T9EA81xlPD6GG9tTPpiVam0ox6ccgY45k/RL1yLrClzq00vP9xW5hn7r
ejnm9BE7fFkRPWfR61lxKiRBaTGwsDod00KpIYW2wQCHiYZ5XYpQcouQh/FGzDtI
p1I6ljh5NKUXx9NyIe8ClbEJLTxUxY8IcV6/f9hTJktjmef4tqMczlwWryLiI4fd
iafvX/xFQThZ3b5yeFQt97E6Ri+bGP0zdv4XcY6x7jI18sWluiqaR8ABy3qqbIg/
PyQd8fur67RmopUW9m68HnVmsGQOcvb+6Gg8RkJBVU5kMinZAaeNuy3Y7A5naz9/
5ikhNiXAXNxbzf0JoL10ooZh62G+afjvJl+97GbVugFpJo065xUf1/tt+zbAVBBx
eZ8Qq5nzdn2nVpkz9xSMGyPHXKDlkK3lqq34XC9ioXA+YW221kPzDwEEiAuDqRPo
TLyy1JaYP2+R78lNp3lJ6Rgn+h1CbbgEN7dgv4yIiV/JwdWrxrIQjrbFrsVFsjyw
DGhGob/yddARSXxu/eByVgnqRYHmUG7SPwsWBavdHrk0yUT2wOwdrKNICar0hVNR
Q7ZFuPGSmLBcvkgqg8IXbl0dOoMjLpTeFkG5gFxdLOsv4TMzVfgloOxgdK+YPHAr
sbNQv/7ETKMkmBi6Vw5pnorchCJYQVkiqXTmdWYLBIr5EGXiqrd4sEcnD2y5zSRB
0/p5Y8qC3FJIEidSF3LMCdEeo8Bo9Xvg/w9CFTT2uu4MEyzq7Trx5L/GXe/4DLNC
kqoKQ3T0qGHe8/GB7VBXHbHbYiZp4pAPW031SjNlreHQu4AXBt4v5j36B7CdrMfF
5OVWv/v4/VRKQ3UoxOxubu7dGCbF8fyv3OnlbzB5kDN7391NNYqNPLzOSXg5KWYM
Ca0QxiE4Vlq7rd+AVjybokl0Rh7cQOqPxvpoiKpGt6Opv1LLKzxIW0/oTDrcNGif
G/jhaMQLkltJFzYzy978xU3tKgw5autpnRBwrK88vzHo4sRfkxMphT5cUohMLOqp
NbfuvYyOz/IWsd5HZKu++fiQtUHFuCtzYOP6CC9Xxm1c5qY9RRJ2KZgEXWlXLoBM
AQh1hhv27mfneo4nZyn7tj3J14GuevNYeX66d3/r+N5BtCE3zIavqqIV0iPLPxov
43g+B1goVDRsOfiLgDBzTt1KrXRn57Larr2xVw1p5Gts1ddw8ickn8cBXAQ3u7wk
eh8G5Aw7K7TxsmoNdRQtohX3BWCaVGmUvge11wN4hMI6c3KHwPdVMSpX0IGq9REB
ARK65GuCH+TC/31+HvXUmqSSYAkmYrk2bmnq0cTOZHcnIfzqquovk7kUewbkhzGW
hfu2jyO6Ed4nUhGAWidwxPe8sP+yjs7rlCbTbaqg+4x0gowPB5q5pMrdZjA5n/ic
xM6q4+CB5mKhcLtbNh6rllFAf7coW5LpGl70MSBYLZLatXCuUtLN40XsE9qeVqbX
D2rhCa4Lhri4tWSfHSj8N3niNqfq+99KLeMOeHSi6Js5ssS6NisBpYan5fEW27Xa
gLi3+K7XPzg7Xzpgmq2lsWcRqKboswZ2b27cKXB1Ys9C1sC9MjRdoBRPDJs33+/v
G6/JVOXpDcOSu1/OXis7v3OxqnODH6hHcIh8h7WPjpSdfI3Oik1GHLEq7bB3d2VJ
hTltLWO3C412Q7Zv2wb+K/l28HbemgUXcAZRks+/ef4ynLEb+4PZqe0JZT7SlNSz
nN5mIivwLGQufRzKd8iNadpNZwEF3Qqa+Wsup7ZfA3pO4dofyDsFjtG5Jgbu5bBT
PaW6xXiHDa76Y0z/1nSUQm4qhyoluUYLr2Zo5h3H9gKNsTczYPfvoXDzuqyG48y1
zq3hUUne9JPcVHAkhJJm++oyOM/8aZh0AohtxyTOwOxSym7GPmo8uCDb5Z/YuKhC
+shWgaG7SM9FtgfGtlxeXUr5MsQTlGHVanFCn/WVo53tNNTRBUTUYDBjAc9zMkkN
zVeGsnjbT8QBlSBgt+JSTUBMI6fFMtb8ByAQ+vxMUlXk8xMfQy8TWow7UhJGhX3M
MSXHlI/x+YWiT2cBcrY0HBHl+k9PvXKN5RqpLKU4c50jKQv+5n3+vNdLe+3ceTJc
y+lZkm5UCwSAek9NOAjvRbF4Z/nNDoFWYqvJahLCHYBhUklkVZXkrwX3L/FWd4aY
OWQP4l+smRHFfbQFTCMY1D5h6b23gGpl37aP1wlfANEPnGIOOLOjC/Y8QZWrhHWs
7wjGLDC1ATgRKrm1j7GbLmRLGDQWIJoprtsfIGE+jnillhrYIeV5fOa478fJYK0P
e83CgJWK0m5Le+/yJWMdZK6XRamiVl8vxGEQ1IjTeTPQxBbUEHNA0BELllLYY71r
hk8+ijaTYmdl+KJK7+F6BH+6K8ZSUAoBx0VWN2LsK1VtcG2WF/0Fi1N6GCxC6yiD
znt9bjcIQ5fuDE7n+w9sm4koboLsv141Z0qnXbbd9PfkHJAytbSYjj1znRPO6URF
qkaxykhwE4cxIU1AaO4phRg9CvhN35TfowYyynNcAOtL9nu+n6j5qsYIpYNDRm76
fkfY3LGSqdYbKmrvi3GgJ2GpwoHA4VwU0pTLC1Aa3LJwsqGbxcx7oA+l8icJAxiQ
5k0tot/PxbsIlO/zCHYlRkVcoD874fa/SD5MjxUmcUg0hL13k8OgSqnQttw4nxN0
QngjbKTJ3Bil4nW5gbQ4jc7DNqjEC6a2ZX/GOtCH/5S4g4BfdDU9aJFw7ryzsyGg
QYsObLRbj9efAdfjaA6RlDq3PrnhbMHhvHbqcMoZrweNlefR5TGbMgNEmcQo07ay
FR7C5sUvSh3UX0QY9jqPfw4yLxYud6DraGwoENpET8c6/mxVdlh1uLI7yHrQnKkb
HzBGVeEzEmz2tTsJR25jbDmQFxdlWKhcQld+WNCo5j1LoPtmleOrPgNEIR2ws6F5
fRaS7/6XNKKjskSUxe1QE8LEXFmq3ZyhcLMJqs7N7CWDDCOo75q4/GQOSP9yM4WX
2k+Wl9JQGwLTjNtl14v5uw1XEqkrR9S36IK72+4DagFBokPqv0nVCg7hCOvhW1tD
FbuO5GKVy6Lc9QOGkaBSSBNgvyz1cwu06qJSkh+ZTArE+lxiP4vX6qlIx9xnd0dA
6yXOEo9SX48DdKb/en0fe+BKwEgXfjm5OGOo4QgcdqCcEayrGv5LAg3KYNI/b9pW
2Qv4zMwBiZC647pvaHZpxtic5DivDegfhcmRvgofSFP63D7LNanpnpFls1bXbbnB
aLao6dJoxnar8uCEXLVQB3OhkCKS8n/xMlSGsFeN1lnK9mfH2mVU7n3D0GZtQs/a
RdFyR5TZaQgt++/8mkytZFgTBEmiI2t78twc0P9PvEXLfhCsdBq0omkRHAyeWds+
3E64n5IxG7YxUgXCXelGVrDH/B5O/7vawvODjn5doG3IIB25yRCaLsbo/NnubKYU
SF0sYS8c0sgBXkjmyi2hd4u7pUVBuujnPOacREpAs8J0E2/44DeMtyu+bW9uXdAd
XxMKj6yJQSfyz5WKkHI7TUs91v0ogLyxlKMb2sJXVWrDOgQDg84t5iPjM+cKDVj7
3dZKq1rPbZC/IcEGyruaAiC+DvfSDUdowHx+HWcoU8jcKJKm9ykfyO6YIlYl/kBX
x3d0Whiaw1PxK32nAg2TITxAuhnM+teIXeGlNRSg7/hafbb7PN9D84TmA7OGyDQK
mgEdW+1bYuCeo04eYglkC6ExyR+9yjHaLrVig2s8p7plVL/oYjheKMd0H92UixlN
OtNzTaEqm4FHeulVbEJjOtNtb1VpDYl/8t087lZf9ZfZsY2z3Zi7wvagkbs1oaeN
4cGgPRMTNxQkahQ4IcFiWM4MNKj85Su5exFZz6BEAZxYuZ5qoaaqmeV/pT4ln2xm
tXYClD7aSjQ+qhFBGDaTdIYYTEkT96+fwbvyLByaH2w3W+uwdvjXkufk4TLpHaPP
hm/o/nYthU4DXcGGd+rwIRkJS902tffJfaCERKDvkDRcS9PA8+3uCvVufk5uijE4
s5j3z45Ks+K+/K9y9UTH6qiywuu/Eouqiyay0ie8yaThwsEwAIXJgfpuCnksJsez
s0ecBL1tH7JENPEabPqewGBX4zTnHRqgfTTYJHS3NTLAHTOKdPuUoQYu/RzHKCIt
7YcMZQtgs09go6eI4G1myVbBd/wF91qVft2ywxqEWbEdm2/AcBwWSprvSY087COR
erXh/uITrKrOZ0MFTV9eOCmZdRt/p2dMXTRgAY9v5VCdTNaU4pFZkpbh852fwXAE
2I0rxhXLZBX6i4neSwfIcFV39dJ4PovIJOamzQfOdBC9jihH039ixa7r2caaKASg
3jWJYv/5F4utf1QCxgyjm8Xu362Q1bwtvA1uq2MhTXbEk4t5NCL6Autq0QhtNqb/
d7YT8UNm6NmBWm+5hi+j/d1pshWFvJRiGFJX3n70AAdr4YBa507HdYEz3uE+4mKi
Lx8sRa2tOYyB0FRz6cEhgME+SS4ylov0m87upzaT82QANJ6HOkaJ/+SwXBWmWO6I
K6gUOkUWsQgcrc+emitoEBHXXnruMo6NpYyZUcimFEJ1x/ZX4NG4cM3TWiD/paAT
ExKIKiUoaLwikWX2S2M41xUZ3gPH3+7ecdAjjWpSuH1hduwOiQvG6VJh657wj6rE
YguYIiSl41Fl8MqHWWzrz9Rj7nzcfVG3ASzs792BM9DkA7SYDCkF/kA8K3Vj986+
PkVillpN6Vq0xJ16I6A3TRMPguYKIlm7bmLo4M7WRpwf+cMKR4m8Oh/zYj3wlQb/
vFW+nQCJb4iZpmg/QP7mP5mnEFZR5AOy+PSMk+KMoUANgpTYpbHkIMrWB0y9rexr
bbgzsxZ2OnlVQ+ay7iaV5C1vlz6qxOh3Wbw4HgonOsX9ddFDJww1TiMpeCh8Jduv
a00ce9r3JyO5PkUAUeCL7pCFY9K1gZWEFhYnWcylvItM7lQ/sX3F95tKjQBgvf7c
73exYOQOw8Qsycl1Xa0lwZ8Qa19lEk3jCBhNf8erJ0X1iLqPB16qQWQcSF2zc+z5
RpnyiTQV4keWSGV5uoGVA++IPur5Qu92jCptnLU4NzGFEWyNLnE8UfpZT65bCcWj
7yXMLRAeOjTeF4kJojnxCJ2V+zHuWHlCJ3U14Vtjr5+N3v2FiYhF5lBdMKnpccJo
VQnCJfaVtspq9zLkBFi/2MlYLYDnn19cN82HHa8kI/UZS2OvmTRkkgRoONimNIdH
G9i0n6bh4WrTMXNZ0tq+0HgFA4e8XHu72D3H0MMQr7nfTYL+WGUckY5CjWpYF6jU
tlCeLZZU8vmRdnEXR35y8LrMKY4KqMUBKqgfIjbLS2yZh4MDoNGrm7pjtMqupsTk
c/Dbg/GryJLP6uinNa7MK7GjHDXiE1psQMAF64fyOrGQO2jhQyikT5/z2H3iY3c1
Lj50mw2wYc3+w745aqlat9CVftRtqoRUJIddAqdfdCYc4z4H1rhAy6PjKMRYfEHr
haKmlQDiPJJ5PpqCntBAul7hbVPMZavHCKXNA4hL/sTFfbyCTWyerrWzwmsGuuJd
L2ntYt+aZCCb66SxmUj6AABiZwwnklPPvWoCw4AJYKcjN/gSVN55Gl4/QtIRzaVx
+PG1XvhX8/Jk/m+S/Y6uBSzXvRbCYQ2u1TSCAXwEl9rB0NJEvrWZL574JRSc2WPF
xfGiEWohGFiS4F4W6UxeIpiwkaHKgyOp1LeWDla54yHapWjpd3PXK+6kx7HbfWye
Hlbwe2kJEBTzeQkf2q0PS0DcuJhasaDc17+LksYqKx+jEMr4yYOViceo0p9Xa1d8
MGsvGFfXBMvRk0rJk8FsPp6ONXOO2cUmKQlfnVKWOFZlS7RQFLm7G0h0OZzn/mFv
NMTIlbzig/oB5aUaBJQ9ZREA8U+GCLGyHwcUIy8/EMdHV4O0zPMKPRZ+b9U7w/1A
jSnlyb4bnt7J7wT3gaguADRhUpZ2xC6KEjSXbyI+gRJMSEjuKaDwf5hCwrAvK4Ya
lsJE9SS2kPewKwlha9Lk0Pjog/ncMEF+bHoBeAVxM9Wb61o/lIW9xvT6uyoAPkzn
8F9D2asQ3Ur0KWLeiLw/mFyZCjIUE1R8p/Rz+SkQqwHYUdpBkWqabVHZZkxrKpIG
5VDUCJRQJpoKSmvDurCrZLP3pmLohcUg9IF6CSgDLboUb7Eq0v8pSudQdzuHNcor
7dV7MSM0WWAVDJ09iD4N6pfFx6XC/7raiiy5loO/s3P/jQHgCnUHAYYDtE0Qg5jS
Kf6GVBMAU70XNxDpttlHaJCvEFDBvu7C66Lk8NSHKRbJaRYceXc7/xSGYeC/nwTV
pFT/3MXRMOEMUrsf7JK857tPGN2Zi9KU/iZ2SkEu3ddIp0U0K/u3xUYZt9n5KFIJ
4AKNt6MNFHzGzZd3F+ttcwo4U7aIFatLHsjWjKKji0yuab5Bun6LUl/p1xXd7+5f
uFCWeXTJDo2pfw0UGX9usnGUpJ23GyOL26zzOo+dGa96fhAtX0TnVkzKaPqscA1T
434wNGxA6rj/5En07T7KzPRvMJ4JJ93RfATP987C4N8O1JdR138EIm4ph9ONLPjF
Ne7oaoS2/9j6J4o5n2/1ZZKB/IDEJbljDZkLJIf5vmlRDdVZYkf1HN2xhS4poLQF
Nichw9do9fXk8H4212lI4pJglQGHHRnwMc/YlixvhyjPGBEGcdy2b7TZyZPlmVtK
bVG8xO0uqWqM8pPPqnoKeX+2m3slwWCAATTrDdXZzVwelAhtFYJO3PXSTJnQKQUZ
2q4Wyn/juq4Zs/u4R6bsgRt4AOwE3CR9WylmJor/paDeeoES60lZUhSaTZH+mFRJ
N/QmkVjoi7zIsxmO5ZPTinqBkTL8SDUgMEt4/f0yR1oc37zF/sDVR6eSS1ca2eR8
RRq7DPu5fjH/hPChFOWQ2nZ77+Mrmxgt65YEb8sQLYbdlcE/sCxUjKylsP+gU6ZQ
D1NC5xxoU4a7GMmw2qG5QcRAEFlg7ttWoIBkGox9888dFy/kTm4Koj8CaurXzmzO
wZQOaWHTqgNVAFDR4QooIMvxUlRPfptdfSBG+HMmX2JYP3wOVsncs8/9+9eGgTjv
ebQoTp/2vTeutpjhOFv5d9wmfR25kWfkxLcjWL7m7RNbVW9h+sFX5PdTEi3K8v7U
sNdAVJQeuEMNOzEgPjv9j6mDutx8D36kUDiXhgjNzUFguQSdtwUrakZgWZXWwPve
cIHQOv1WGr5oBQwGRV3ZmZdcpseZH0Rr6PtHwPBVfp48oj6co2eH4HL2hbKlRFtD
wgM4ODH0oOc5A9aGNxF5iYTn98VHhqwPaIm9Na2kDYQxHoj8vjU8kz4j67WfuJPU
pLYjw6h2XOAVWTvXlqtXUtNOZbJjCOoZDUPmR+O/ub6kVoJ232QDSUtx7lSECwMZ
+c2dBk0s/5W5KYGU9FyvOkL6fPmhwGc1IIiqQxtlpflrCUJQ5ZEveEIPZxgyx7dv
3UNNIOvquYVzoqNxQGhU05jq4qJB+vjv/M1PfHmVp2uxmJ/ly1EvYj0odON0/gkB
ZYUvjHwMHIo3Dd1te9udC7YNQwZ+dW1crQ/DvO31sJeO8ke/t1W9F6xP+gXTy4rA
izvxwtBqkkD3KLU9xNteMl8zWX9yvpBfYLh119RjzydPRDSBzz3oMGlCFlygI8AB
TecwJLqtJY/RxYhyHsvXhwDM7R8AWJwWED0GxA52/eSZZyWV2U+4otTJq/watnZC
WIyoPBQMRuvgBcyrJhsplxte2Rr5R51pTwULSag+3i7iOkdbz/RsuES1D/3fcqZo
KN1QMUOXd6lClV7NQn8/MsDK3UjB8wbMySClDuUG+iwil0urDd0VLueHCUTW3Qnn
lVHil9Q2/r+M8FM5pHZUUC0mghg15HAu9YAnc0RU+fLTkiaRnuMzBtUp3OFdm/HN
of0xTmsvWXlM6roHeCTQfvksmhMsJspkTZ+i3e2vybI/6MDmf92N6FGof3G+aHYE
0oRS/zSQ8F7HDmRD4z8/IbTm6lAPZF3BT8eJfKtnKW7HKgVAOy/evD+OC0ZazMMn
bIfVCVzvvvOPoeRlp7LoxDHbOUjyAVxx8c6icU1Uor6rGZfJSYjGQaZEH63NYP8e
s/M2TX+Xwkro56FX5Glzobto7yWLxhA4nZy310QLo0d0Gkyh5nyu506ZajPPajxs
KtMUmUKp2x/kUApetZNqogmJGpSMVnEiLsZKZeREJjAu8Bt/C5ZvrTw3Xq1TPvJd
Wbr8KOJ3iW1LDzNdorTZkE96/ZriYYArtYJA4BRMMM8quB3YyvGpP+5JQGmtZcPV
91ak1Gwt63Zjy7rvr9Y5abtLscZyWt2jSGjtX0UYvP7sWkj3V+mj2R7548UC/r/k
SvjYfiYlUNSQ1VZSu9+2mvkdR8yauW7MlOW5L1cDrDpX8YLHrxMLtG/DTZdymloX
8k3Ky1bJiCek9v81fDmKW6oR+A43nEfK4ZER1JdxQgSUJkq5jJdSsbQ/JZtuuB8X
nsAmOiOdxAnP4lF1NT41d4IZzztMcf5sOAtNZEPYJ5HuG+Er/VgkINa9evkLJaHS
L4eBi19BQ256jShg4lNLLTLoIm+s9YkyUJcdTLysEsicyAuSPdBV+RUlMm3GaNII
VWOXrzi69Z+VU9F9nUsl9wAQjxWtak7Erp6lIkLJk29bkDmNWTSbu9OHDGe3mG/R
ChsDyfVss1dQdLVp2n04QOUAYW12zu2VnHzzr37MCwEnNevgBiNm21Q1IEemvYS5
OtNW5FsUbK/K/b7w7Hg/N3waUSlOoP100KW49qOKK+dgZEkgSiPhtFJDqs7XELls
Ce45YIsfqXA/830Dj0P8fR21RRlyYVJWexAbp1IAv4kBGc9rjMpFqx8+S7z1czAi
dC7lFyJQP/mSa2ESKcsxUg1TJGNdu6KbFumO1VasgzL1GLP8gwWGK4CaXGZJbJTn
gCT21jZLYLtP/RZFBLKCFOp5Q1o6u4EHl+Vzgf1gH8+ndK+znwa9KlMJViPNC286
8JM0kedXsMqQvCJjuVSnp9kXu9+wOT/UJqUGgKSo+rw6POq1R9Nag+htBD7ZKK/a
9pA4HXM+Y5cdovHihdOtOo46EnrRTqosdpLu9mDIvCXZCyKlY0oCK/rezEPdqg9X
a5cYU3qR/qQEBSYtzB0Z8s0bXNu3w4zjsrYdtU5x2KOTIPZbLYZ0RzxrLsEq3NH1
42xI3gUJGkk50Lx7nrKCTtaRbnvz4dJycp+1qBlxmNSRw1VftxiBUczOxFt1hMLF
x+M/uevGDGR2GSDZy7Bkox68IRxr4BGK2Jgw1jGxinDATim4DkdhbDXMErnMpEmN
nPjkCETH1+uO4AhB+tksrUveeWvBIVVDfS6ZreDOyQ/cvC1kO8gvQ63UU1DrHc98
sjnvij2gHotKq4k95h4QGq8Wc94MHOTQI0eoEhaL1cgi54VGCMsQFB1OhqujWO6X
1+0zciykWuDAw7VRGG5hllayO+RTOQDMhzkp8oklahKv1yys60xInYg0Q/s03RXa
kxeEBG6vE+bzNhSIMMGuVfXIPFrA4PoqV4Lxrf+4uP05pZSWCSbQ5Tscb7bU30KY
wFpW/TfiOACrllIXnml8/gwKiHAlZPjATiWSb5T5HU6LDD6JASwKNNrZ3kDhcMNA
+ijePE8BsVZWpSHh2FY+zgHOXT4NAG3f96/C9GB9dnP+/ImYChmCjGxHAMwwxsHN
32+L8rKqksDUgpsLbv/mFay9BCZ5uRtVUCB9GY8ABetC23mQ1HXDHZKwKpyYXF01
stFZAkWie54q8fWhfhn+txXTf+KNO6k1yPkSlFPkLAISp7D+YxGegTKHDCSKbXQc
1+GS7IRgGtt6WIHK3H8i2O/rP5rqjssPSvS3tLBHAjE5fhbMYmvj1sGaPldlsV5Y
wAVIZX6tk6Z/OhrGCW7gYsCzeyx0gnqhA0rAYTvN4MgMo3yX+nmZUdcjlpxj+Qfr
acwwm6kKd1WB4BUA63Bj1Y9k8oYivpvH8rFumwSX1YijO4V6iNuiag6V3f6jFfu6
MVgNp/y5tgQflBDAAKwcTFrA6qRqDMMhtkF5HBa+WGNUnBdEvV0Dqdicjbx2Zkv+
p8NWH+7vmj2GfU3Ak1x7cpYw9l1ph5srkbqXzPZqBAe1fjWQeEI6GWE+u/cr8GQY
tvAFgE/XNOv3TT8M4ri5+CiGhzoL6uQNkxZPJ9t6KGDfE22eAysEJc56bpQSlvCq
5kH+OSIw0GDoyUV/D6GfE0ZpuU4+TErsjsO08VC/62fmNiKYgndHqPSuwhYQcuTc
dfpQFxlQxLW+vts4RFr9zrsMaQBba6CAzbStdC1oNg1qMWbRkhc2MhdB3QvOki81
lnELzg/oR7OJa/LGD5L3mdCEOAIIO5qzil0VR6U0DhUKDyqXxJdg1AeEMYKSr+gN
niXSOsfVyeGlnkRBWUmJ0qPDmo1T/fQBjoa1b9LyV2eLURy5/WEi+4BRrOsiFP1P
TrM4h9GyQ3RSYe1VMAA2V6VIxeCWectbNVnb5GAg8xtLFJyNOgMAJtYqdOWOrHxc
73tGYRaG8Gcf5fLlc3zkZu+Qx75vb0qY5ypGtMKIsR36367laXmy9M9byAVOs1Sc
dAQX/5N4lHZ0gW7AjVha500Tqvc600Gz1qCR/uaOEu1u2Qe4Fwq/q9kFOxIq0A2T
ACEUHjbqwBKXIkjo0M6oydxTIm0/MXwoLwa4W9t7FcCORpuQaDZ3mW+SPgb9Yu6f
OQjmuBwCtrOrQbPTpzgineXb+lp7VVMdTHEkpAua1O6bLhb27UmaGk0efuS4996b
yQ25t6rVtvON42/wHndRjtqQ0IeUVQuV6iHcAzMVZEKaRRAMHHvZ40SRkyLk4x34
lTEWnH+410+G0sqTs1l6neS6/l/KuysPiZKvWVdXep0VfdlY+4teNVwvPj3UXpn5
fb+bOXm5J/CM6KsHB0DK0R06vzWy93fbm6QoylbJCNlXJBpfsFLLX9bNPasD55YI
Nzc8Q6II4dl3I2EdC40HrftuJNbBxwhd2gP1Z6BAYGwsIcimnjOWWVbBJN4gk1Kx
zx+uLAHzukrYR9sd2jVaNCGIJ30Ys6NxxRROGWU6+0wI1QuMd6/yGISpJ7/sTe0B
kWJWVxHtBeXjMVp4pbDlO4Z8nQhqRJW8mSdVWp7j/kQ9zCaJkPf96iP33E/6AVrB
HslPcLEt8/4f6vWJgY51C9yKQFJgwWLxXIHLqlmST+GLCTbnwzl7EqY3eSagkTW5
sTeGYQaL1bXj4RR8mLWWpZKGDhfyKiVpfa7bqNEs8DZCAZ8ACiilgbb8XnZrHOi6
vGWpcISai6oBhjcIc0Cw6uVIe2b19vZKL/4LoPGFMpr336jdNj0itYA60tnu2Y07
VvI79ZQTtML/4fKizsiD8bQpGOHMGX2ygAIbvzxds+txihU7r7YAh3oZ0yJ+ogON
jRCAV8ZrlrPAyQdZ0tz+tCaX5k9kSR/meTFOg0aIpU/fQddEhOq1FBR8oFRkPlfh
nlTeZ60QLnah169ZO+AEaprV88AwQq43r+b5+LVTZXr9rHW1z4spKkIdtfzAYyEk
Qpwh7as7HusnC9OWs/kmVfxKB3tNZEaqrJgPI1Ad/lqs+EwBoYbsaupx7vgske5W
jmwmZgt0K/4ogxx/vvzbI5fLpzWPlCEpTN3j9oHYmpvvbdjSkw41vf/HqdmLKY9c
yA9Zfa7Brfu1fN3nX4OzOg406ifPYyDlfoIYSEsKg3+hW1mIwiCRHJDyKHagCoiA
UkZnIigiVWh47Wnu2DKD2olBA1O23FlS1rpcSNRJ9dlahcGzTMTbzYd5Z054gLKU
aezbLamLSH7uFbH+finETH2GShNqAV/6wklx2xRgC8qAbWWreeiHWIQLN2h3YQgO
xKIyG3qU54Sh10SVV91TT09aff0Fc8E0oABz7xr5vSpagOIJoTIByJwPqJQ5OPlG
Nvc3UUePHbki8eSme1MGdiojYgrF7PAeb1THHaF/wqT8dwCJQmr73LVGT2HIteRZ
JTEOsK+wt+NqogGice3EyjLh9jQyinZpKsXVan6tIzZ6lHw4nokrR5AzZZcmKAqF
Ic8k3EthVL+Tj+Hc4XV0GHyx7t7nH/XY8c+SzfTxPM1PFSTYm1vIgrsuk4i5CX5H
H0Hq/Q+I5V0xynUp1gHR/mPdnGcZAiQjC4Yh5djmRJ4WX8wcnLXny9XaNO2Ch6IH
pXegjEHIO5+Q7SrfEEYTtZLD2K15aNeC3IH3C2lmwRbCo5HQprKL+MJNMxtKoGaI
urLTIrq1/IwQ+jW48XA1A88GbTN2JEYAYiTrrHPXT6EwfIa4FAEAZ0PvAuUvwt18
baLzuPqeTPcOVNmBbedMTAsubMPurqFXWwfceWFcceAPtlLoKpmtbl6zJ61GXHHW
Fn0PMXGYVEvvUmQc+R76qe3+1PBhkKOGhROT6Y1b8mlhf/wXq50JP4OwFCU4QzSK
7YrbC6olLglvnHB1DMQds//kSMsRIYjg6vqBGDPjmaUnpigMIltdYYBBypGkFFf9
CvnLdzFWCfZ8Fd0thtPjnZEsmcXZerTyJkkASVDg4wSF9RAJU+K+Lyvh72meRECS
qpIGPapu6s6n0IOSaKvF4YpQuhfzRDq0QcKHuKhnd11HA8I0Jv8qjFpc8Z2vUGeg
3YY5628d++4m8Jx8Zro4KmDLF1gnHZdA4OV97WfBr+9IvT44xZKvlZNuwauUm7et
OyWin6e0MZs0bvmYXtXhXMv1SO8ThcL9xHuG3VDqFm2KOUUt9yuEM/OeQ2xNyi73
uUWdpJF++fkFpsOTjcZX1QRHTkOuULkVmSFHnccXw4ucvjsiSlPjciTuc765kPJ/
Gk1KC6Cli715XJcImkl3UgbbH1ReWTlCf3klsGlJbr3V3GL/UuPMR0axb7VOoVfW
LN/E7uXPL0OEq3VfS05wvu4j8RUqyRV4Jvthjy9RGmPJeB5BQ2wfngKxghlQyiUS
YNBprhhkO/3sZwBd30PY/RYdoSEeOwzoZwMluNn5sTilrRPg0+MIm9NvyMYwGgId
XX0oEklDIEwc3NcglykOL2+Vj8xFqcQe+2W+IFvnGJQBbpc+KtCyjh+zIOqaMbCj
yA9zlzja6VbPGOxcFtSqkX4iFKKrQYR2EX/hFAXgJ+tjbLN9jztUiBIKwhCgqgPo
djUuOGu8S81G5MJlslbMsMbzqmcftu5sDRSgp/zNRX762kmtiyFmU46TB11Ntr/B
tSoDQy3Qa/0slvDRR1BBx+vEpPgoZLQ4NltMSJvnDeDVx+AF45pcazrcwUljgIhr
B3d4MS1RAtCaRLCMckUkw9yzc1MXSSXhI9D/Au+mInoNic6EuRWEw65gffZa3foo
bur03I9K0J7PfnckqTWSPnznFyIG81vK7C8eIRabaUE6ZbchgbLmjSOEBtTQEbhA
Rnd8PrP2kEbE1Miy1GZrEsepXgM61XaFv46HfWNgDxPHFM59ajjCYCDkB412uGaS
/+pOL+dOIANoo1sH9SITlf92EQ3SQ7mGnagpvizybju4WRHnijUL+PQEtUiOEABX
IbBotb2mk37302TXkzMSUoYPBUgT1xzeaM+xXsITEsI5d+6fULAwu1JEcqFnKQpo
Lclr8hvz3/GKPCU7MDfK5vU7IgPCzSRzs01laxcmQ4VpO9C0oVWZSPytXqJAhBOb
D6sSKQTzmYHaFvcnsDVOhqJoNHNVmthZR1ibhRVeApfRhgeh78BZcUjhLAemx8y2
BNQwpEiJKyz2UU5/zmU+SSZir3iPr1hw6aOAbBHnTHDV5RjILW1EWgiTnaBv6ev1
wBpKO45mVplyDuaw5AR9L2wPVNNXbdsgMSyX5WcfBZ7086bVZ4GcfIsCLKMHL3AD
8VFn9NrymFEmlPVzLdoPOzcSLGfRXGh5DQzC4Z3w6+XdCxY5jvKKgG0l0H8ggsIW
2lPwZdVdS96mTsEl2iySLU0CmNa6BDe6m50QQ8/h0LKA8w2CjIH9RVVJQOBuPR7D
P3lIRTFFvnD8MVsJ9sWPxgUUYBpvspngHrxu5uxAjevxDug9vDacGM2p6O+t6U4r
Vyg3JREM6WMHEZoVK98LYes3OS5X1l6/5/vQXFseD1uIXk2UFT8X8ZDUXlaE0njA
2WfcCchrpa7OuIICPwbU2qrTRBv3mCCStlRrFYnw4+A1fggvs0MPfQ5Darx6yG/Z
Dfke1TEle/iEjJ3mkJkUYri3RF7WvjI8guXYGGcedXDibsl7ptm3F4EXDmecQDhC
qv8q3EP0b+oC4m0AkwEfZtm/b5dIqARrNHLQvNti4uivGDIA7a3LfUq9JxISlKew
Z7RZgVG2GIYgv2R9l7wuH6puKq3/GfK4Jj/sZ2JpEYMXSNAOsxn4N1qmlgLt/XsG
gGQPYxFdc3Ebfo7weTWCwAwTHsXoSuSk2A9sP0zx62CGQefgWo8jueSEViUQ6JKV
zvXW7mRPQvmQL/V8wfrt+LpFHJI7V+imwIQ7jUMn87Eq/fJZRz6/FRhRNIR/D4P+
t86lLEpz2q6Y8NKELmQc/tVF3pkzgZRv6H7k/kHmvq+bYamLgEXbq8jE1QzfcxzW
xyjpmmtOCv+rqONzmRoAlgAZQ5WAzKI/AT1hy2ZgPpMSh1JG6qxXP12oCkpnb12z
M1XWRBdvY+tvgrIERPjlBphKyMIEaYMjFscta9INcKU2gPNxtJXjTUROvjkw6vYy
Q0hu8XcOy8utsTzIMGgWf1keoI4P8rt2zGTBdyR9nN206FQocXQk7tLYtg8Sk0Wc
96hAQWAn0BcO5PwfFc2MVrYAG4WptEBa99qMGYIVefHf5ptVoF7L8sXeOGkewtWq
/lcg/+0tRFKctnbsgB8NlbzgG78v/+pHnxebsMZaFAX1Mt/+3mKK3C1r9Vt+TszT
2maZ333On2ECWES1tPUxYmyrQsLn6babssfcGRai6SYtWLj03ik0hKGWIcP7Yc1E
cmTtkE6UK9bl7Ug774OZT4sbtgKzydimpuWcVbhTDTf7IijxtGoOPI3Y2CPeY3C1
so+yoEvtupQ400s9RSHbAFX1C0YhaZbc/DxjXeX0VNZnp22ypMIUPWMVVT16SQ4X
Aahq91lwDi9G2NQYWMeDYhPW34pUDNaIL3oggBDp1EAjrPRr48QstJpaKwpeXRl1
jK7RxHfakhjeF5blZgtniDtsHo7QJXQ77bZJH0N0ooIb96uq5cbXGK5T1nLFOqxz
oWNkKIhmQO+KnmGJv+4DvV+D0beMKYgbzIrnWjE3l1O41STSv5drhfp6fjB/MMJw
nnvWXdbuO4TZMOhJAFyl5qi6Bx8cOZtGdYcbOuuX5QAo7auucvon5qZXn63xEbOe
AHm52/wTkmhYb3y+wDmIAtVQACXFgDeqlK/8uXcD4lF/GT9+64c/RC/02u2PKxp+
s2DCHao10MoNra5sOnW24EKT8Y53xd8fsFwTyxBP5cXW+B87ThwSZdTXohBeH47x
b80xx3L/hEtQwtCII2mcUIdeLBPIpFlQvgIMtFJDPgspZf5vgbCKrZueUlVAn9Nf
0OYHvKqDj1WbzRdWrVhagkni7iqerqXb0HO/cdQTERafJxxXQvEi+SYa0FpfFtVT
wlVDfRBb10JBuq74ZjF2ZW/FnorYSV/KaPCEtHq3pX+49+Sy6EuztgOCk5hF+K/W
2YYsmbVVKTXUNyFBwCX0Qb2Eyd3Hl2VoPy+23C+7Tv9hmeVhsjSOmuzJkkbPzihY
620/okXVdIqKapHh4pc2pvoDHNgvb0aYEFNaOjn2D91hz+f9uLNye9VYgYQG+e6j
mTn2Km4U3EYEz57yPN1QxrPN8A1Bkz32A9KuHwX0JTlV4Eo9uJHjTM17ASu1xHmR
byX48WgLsEKWI2fUk8fI54Zqu17lzI968vMedz0Kcg6sq2WzdO6e4/+qG/k3rXgH
qIYm1UYHmI3a5EcMnkUMV2ZDkJkZo0wec7ayEWM0cDapTIk+xdvFAjno16vwSVt9
5SdZGzPDk1VCMkHOGTsB1XT2/YWfek6AhDE2meW2TbPbQHXBELqsMWWFTC7dn9N9
mGdNrg1cADp80uSgPWEGmJ51Onx38y4qgNO9pfhBeTVaM78nqXeLZaPqM5Z2SrVA
3AUkVF9ds9MjR1VoQdRwT70agIVb3xwQqW9mN0qthDxjNxbf3ep46ym61T5OpeEa
PMqba4b55tppZB9vl3c/HWr+tYQrC52xaDQKBa0wj/CW6dUHoCkyt8fMFjnPoKPR
aBwZRM89wR98Gt0cxFLJiiop8YRi8t6j7dMsQpgBNV0p147AxwOu7jJgJUwJDLUr
F99SBMWrRoPVhpzkbcebCx/PqviU+pYD44wQOCv/Ih4qY/59Yi1pUi6DO2YRDdtW
tfK9TE4Jj4zmlkXCL1XQmDC9+UTqN9SKO/DjSNhipNCfTczSGPo0ZN4nTJ/btLX6
dsl3tkLb1nGAtQLPsWMdOHgg6lBZNLRDZyU5u7BSwZjQmYK7EhyRIiXB+wrLlMNX
KwU24PxH491uC1NwLIkYTya7+hOw5ZbMoFwnatWo+FD1Cwwv/vGZCCmfOfEJfRt7
3mqfTFV2IFyT9AQTLnPgPycoaf2vNBzULm9r0dPP9H02nh76TXL2GF6AzDG11YaM
yghstOYrCLEu7+KRhUbGRCPDp2ZNP2bQBZlhftzaWh6yT0kFq993KsTcCE0g53w2
/9b6kZ1jLRYz4GIWQxOc3Ob4oPUHDrDciyFIEwLOBB1ie4fX5Sr4G5aNx9xhkui5
evqpXmSdesjSYhcQ9ZQJlTnlcprohynNLlSAV2Ult1a5eV+EOHkMC5qZAsBV5oOH
La3ZXmzybCotWuS2mmzgxSGR1mHny75jPL8Ihr/gVZfu9+8u87E950Jqm54OJzXu
/gnhRGUx3H539s8Vo1AUMw8hFHFFcU9bPKx5ew4S6s0Gl6h8WJDNopZQQhhi5Eqs
X/JBjVxtNFwlZsC2N1H5sLyfzTN8fBBmG98xWCcGoizzUKdlhJF9Zh+wZWWfQ5GK
yXv3XhILe4n2vlxWKKCZx+JHN76nh3rEKUw3vGl5RIEYlpLKAL0QDEwajVLXHTgw
TnwmwCWqwDSPdfmipiE1oZlX9X+te96lAO0y3Wkr/yg2UbIE2ZIjeVmPqg7SnWXl
hpLh+BypBwqvbl3nnP3/bdqTZN++oMnW7MqhZE5F+wXdckghOa8IcFL7RcjNAFxs
m+oFIVVVSaRlQkrdZK/mGRPyX3/P+pneB2pgg7FrITc2aR9kLBHKOytMNOVrcmMm
UvySQ0VWrxtjrAEKGWpnzsMoqL41js36wVJ4VDj3cEhZpH/Z8pqOQ9R2d+PqRJTl
fmaJnWPENItEvhc1Coj++tMZDZf99GDycXKFTDBwReZ6uhYLvc0YzOVQEkSFSLHS
wPfxmEIxBRBUoS8uzUeYKwkGluMw88K5Wpu6ops0ZPlnNqAwvVaxWoCY7fYM7ZXB
FMowQp9qNFvKJSEmOUYK4/rEcaIPkE2I9czS8W5va70uqemoTfnVY41qom95hIp8
fEv4NZVQH9ezelqG1G8X8I7tiq1ojKG9DD4FjeuxpCtx9Dc3ce/Fw/OrngWhpWLl
v4vjHEppj06b9O5hH87uS7Nt0fXEFf0HIM9GftgQFQKjBbVkdXQitdsoo6VWGHMq
L+2ZxVjdNcxfsB1ueSgqHhqI8m4b1f7Vbn9YqOMdwKHpqPcPO+KYeuhKsH/ch4/A
LCQHrQiQvmT9xPW2efb2lDXq04GRjnN5f5thcHh135c5BwLy7rz4yYUdxAMU4yBK
wolIzUSBcj3sl1C8Yj18oQWTUBLT5iSjElEnYd4BjaEuURjnLsb/epoSK/9BkbjC
r24ZQ5hctKyRtfUTSQgrCIoMgU/iO7k/AsADgoIJqkDHbkTq6zVxNb5x8GYBjQeR
c+xHIlE+C3aCvFIPuvZeKSr6EFSRglqQoSC0u5r2qKEh40RzibzQNLEKQ98h1nCM
p09LEhpXW2LobSVq8A0yiZ/2ngRVKK8ITbgS3CBIBGL/+EibtPftfSD/xIW552OL
oswipFXu+q5QZIf2hm5yc0cCKwEEaQ3Hjjh2vlOoXBhqgodrRB4jbaVjjKDL5l2K
2YPX6ypvsFtRiaQf5I/+JO4Fqiq1G8bQRkjF4gTLrWpmprsVE7Si1ivtCNfHb/NS
YoXGnMry1bQz0UZev2TdTDam5zeRRPDQBvo5rSVlcgi4lqQUpX+onULaGrjpy1DL
JIbSAd/X/HBPnU3Xk6+yC2YgvbDy3Vi56bkKdCWEuUpEMy+gE8Fs/wVyL0YTN7P8
2fPYrfbXyxbm+Mmn7ApvJbMbApB3bV7AYMVAysbmRph36JGfa4SRL88mCdlyYo0E
dc1yqRdH3/FNVqipBaBALMqDj37OhaxV84KCV2GPRSkKh8aFgWI9gPMpAHe3R+c3
b224GpqyUw+PH6HsbHXqjWBzAV1HrCQkF/NUROM7LfUeTW4eZJ3/AXgVEC7Xbvxe
nW/0eGn5VDArb7f7nFKg647QNIQPeoURw8P2AjfE9aZbeTDiDlKsUpCpc6xbqIUP
eiaiLU6pdlbSD6F5K8V/iM1OFx0o1Mg3NEnCOtyF6sCTvp8PsNEG4I86SJMDpqkB
n+fNKeHqsiax8e6qpYhxXzwaJ6H6uYAe0GCbdlgyQoAS7J45eMHYK9rdGUyioJDH
51ZqZ57z1VRIHGp4KD+SeV3DhmzMPLKAZXko6Zvt+1fSh/Z4j1kqddbNRgz2k8fK
L8S6vzNjMFfkRW3ehdcy9AvBpZIaO+QXQT+v+PIN6M2fX59emZ2qJODmLter5q6c
BtNpVWlgH92G9pOaUlwznSkMM9/pRe5tTCkswCryr4HwVWHBzF18JranslrdeVO4
7QRFLgCCIMk6wOtvpqZ3nR9g+ndgkj4MWQkaGa6IQPl5LEi//V2ObZf3pdnpyfcY
q6VQ7abf84CSXNA6HpiO+i1rVoVAqaqw+yw9+lYLRJpWS1plixFkmSWnEwKFZPMi
rQGMXf8QigXC8zR2ThOYR72LILbTvW4YBHHfrCAlGhO5xj0zHI5SdmfTUct4fst+
MWZXhVm/KSY5Jwq5BIpR/p+iqDXpFRzL1G1jOYOjmMWGPx3yGhNS0XKSuq5lrSMm
EmRR5vVYCYPKYcimR1TouBS02ELC3jL1JgW3i66g9vVeIG1QDeFHh3P4nb0OWbyc
A/2AqmX0Iw/uJ9wmZ0byjfEb+HLd8bEMYQzH+6rftaVWVxllzWwNtnzU/CGIM5cI
ScubJnOuIm1zxskhimhiJpVphveshikSIc9kCZQTUKdBj8libM1+4zr39dYW0QEJ
TZIXKDSA9ADRgz3kMa+0ehrN2bdBGTnB6+J39Iqj6j/5wcMwOSIHKyRfAS+Nh2eL
QQ0kFdi1hV+M31FW5fz+ALz/VCKs3B+FdfZyR/R7gKzYTt/9xCP32YRw+FhlWaxv
XAk+hCBBbgNRxbUDuY5YwSrPBDi+2lOh2pSFhKxg/K2SD3Pg80VeF8yr0gULQopU
F4ZGVEfdkkWCowDnuHyF6mqyg683uKFzHLYGgS7mksxYsSxySvvZQpHvW+UxIS2V
Xbq4xkpq2lcmKMxLJlLxw/DjUbsfXRLmlTl6CnFKgZFV7AC8xT59+GnTjiQ68saA
iMoPqqUZVjqk2e/fXj/Pys/f+JXPnlYxjd3YjfDVMWY4gS48R1+G1bDGMAXhKrb8
7VYOfvn7RYqf9pJJn4J9nulENRjQ99Hc72LBL4TwH1UWlFL+yvzy4ZzXUTUQCDbk
DRJay/ML7IrpyyJQeGsEKBuZQeD9Ttlg6BEdgD6k3MORano9kbfmdonVbvZXWmVX
7xrdB4dB2Re85ZtxC54Zy1qGMDk8TmL8PaXiTnwNd1nEiP7gyU3wCejcH4RpqPDn
1Itb8sDqZFcU1F6Sv6bRScB0Pilsi9yokFFU49T81CxI5yiCA87NBnsw88kC1Nh7
U5aaO+pTSZwULvW9MmC9ZwCNwBJ65aMMK2zG8swqoKEaCPbQsNs256Gin8Waakb5
UrMSweWi89j2nkC9/bYNClM+HZvgATSWhDjvGqM5s50G72vLMtaKqin15TPVUkd8
Ay13lDUTZYlcLZV0Qv5DvkcweyiE3Mj/zoY6MfofP2xw8cdyqfQbwGNyREEiWIo7
V/zcghtftoelCS9PNYyq7QhatqC4xqoiUuHCpjxcz8ylM1B0x/nxRMB1nsd6Q0vS
50qpBKviSC0gMj8AWL72FucLG9o0KL8nxIzKwszlzUVlmeEY++QYh+daENgfNgC0
/3GsS61vNvcW91hwUiimfbzUo77a0fQJJ2qLiiFU05zHxy9oEO5PIjGeHsN61mPf
9yhHRs5etzR/CP3VkwAwgOuHjHpk70ab8m3+Xoao1qS7crZ4BC7bfJQ93my9vVdS
yW1ytu85uHGi4BOP2vrNqhnOF11q3PEMGca3uqetuMd7gZVbg2c+vmkjLOQ7WDV8
polKF/dXMwbIBWqsZoOFEQS1NM2qHeDkbQt2wQRAP+suUkdP+yfs8fzVCLE4JUtJ
8u3TJzItJwsrB78XdaEmMK8hmge0VbXWTXVtcI3y+13/wDKaaIbdQoUURqbOpi6n
Ie6Xb8jZb44pPtmF5jHO/JZh12AmypXxImy+MAfYv38DQdzQEuB+SQ4MZerVY1P3
VFy6LGui6tIdUhAQnV5FtGdY5Z7z8p5LgP+b1qnZoVeJd1HooTrHNxlWk05tSyha
oYcyQ+DzFlUFDk8GZhfS2RMwEhjXg5B+iQ/lr8GJ8LlJdZGZO95y0F9M9egCuah8
9eQdRCLaBN8NrgTIPQk60jOBNo5ww5DX+OXgdT+M8YArEutlOp1rL2ZAnRaVtkPI
fqeYVMaWneMCjyxpxb26erjFu5fLa3NNv70/JrsEM/J5l31Wc2zaCjf4LsA/aJrM
npdYaAbMSpPZht2m/4v1rV4Hg2YdmUr6i23n8npGi7sjH55XO3GBPnkp0PbXHYD0
upKrpOSPC4F9NrKlzjN0PXc4TAchGhWWIkJG3rPFziAVonbB/TmE9DCdrtgGWkXP
qGlvTnisCQ3WBEv4w1WT4CFtAV08zrYayGhufRXKTYAOM2W9ymniwdmlFMZG+peN
e8Sj92eTAfvB6QIGr3HUTbhjRwtXatFaVmA6tYfG6xPQw/Ef9PfzKlzDKe962N9G
zVTb2zjqokW+i3Dpc7/rbTZeZe2QCSlTAI00fC8269FBKipARzE9gPkciiY6aLzD
2ADXE3VhXpAHZUmlwNW4qkWdmuAhTJzf4tLgZGAgufEsm4RiYbQ70/TfTBE13z85
nyBPNWgGGmZk/LwpBmkz40VGMBlBoqCLf/fIEVfBdLZ8vOHizHpwAh0KL73wYSde
drE+IaXP0xArjoJ3FNV7+fA3HbXJwWkWiP42pR3p57VdPCWT1U8EKelQQNyqwtOT
jCoeVQEoXfgVaQuDB00Eo0BDNKvxxrZSb68qODFmdbLp51jb/DLJMyGJRqGndcBt
JbbTOCREIEtXGm1FLp7J/jWfmMs0DvJsXYO5DZzII5GVLRPqFDRB552QI1pKsdm1
gvB+b5uXnSq1CFmPhFEzRU4DuQY5ttupG0FCJJXYiy7Axr+RiXJixqcxlqJYAkcq
IcNWvKmWi0TJ/RRJ4PKyP1vsOBxVnc86TK/Y3p+4SAMmVz6fzD0tiDF6eyEef4QB
LDERF5mSm/AmoinZwFWwW+5HEMwNyqiyocHouwl5o+ucJOmd9pCsQml506z+NnGb
Qk56FNjC3KqgCODt219eHSyr9fhlJvAT6YH7LF6kIIrttV2vcEkUr1UrDh9Lf9t/
RYBW2Q/YNyhkajg1fUBUYpK8Efzv4fJRcGbQsJ3LkzT4GvuhHHvT+zB3TfHn/FLc
ELm5yTf+hLYoyQ1nQZ5+/CmCJJE1GhR1mvBSHVq7zwy2z7vdUW4gWtpsyNYp/729
T1pebG56I/7YZYq+vVUxuAYFSl6rfZS3sO1VvkoqPVkNVULtuk+RA2o0WsB6seNL
C44zULmc0KGIErvtHsDSEHUCDmEIQxnUcHssouHo/IX16zfwNPEIIk3KVWkezvHq
jKaQFhepY0AH0bE2MbX3BAM5Z1h9vERGJn3OkKpFJ3f0Hs4q7z0dkwNQXhG8jVLl
xxfYoBUDiy8pkgsh37kGTYPVsmsUUio2cxXcqMzYkWyPt91pd1vQECVycME2ETiG
kkGhifuhHiZ1utEvi4fjq1F21VSODN4JCamtYWjfmSCChnn46cN/iV3K6vdSDqF6
QY+BAmwEiX1K8rKmr9gTvgAPH5qKGuGVIncrC3cYPw1dhgWuRyybigHeBN9rEaGm
hOnIYe6w+8ixxsLGQTmHIwguSuKRcA9DvyL9mHbTCsvxNLx00kaiQXT23v04eJnJ
DAkLCeRHOc6jYoUVWwfHKAjCDAILqhN2Xd6ybZiEumvSuqHZ9WMmMUuxkL0e+Dzn
6unpcwNxIk85HoQk9yEsvA2OX5tLHPKpUVJL8SizDtJpWgJAQlBncKLE8lFELlkm
Pvy8g+eoMXQoMvhY3BsbC58ClYfKx0QhQ8/LwER/exDVfxDPnZNsIv5mKSQl4CCR
LVV1bK4+fvusV3RIx2LfFk7DRoAmBceZyUbFxqdMj4+UhokVJcPbXzxKYc+kT0Ei
qZKehujE70bVY+OqYkkyKPBJTQ1Z9lPBYtH8P/5oWD+0wbjDD7kSs2OBYzY02Tt9
PQSMoLanmWBWllSRsoYbXWR19d35BAUyg04o+1r2yGqVHbkC40NFdCb9p8vy+ift
DijmAXfyDFmw+IqEuT/zuZskjQah0s78Nd/6vFS04eE/BX6aRJ5e12s+WJ0QDaBH
ehTSMGAWyuMS9/cbhskXT0/mft+mHY+rZYxtzP26eYBQJENYjw52h4lAAQioKUcC
0SyHl1jOM8OInlIFLqP9fvkWsEgjBa4TqADWpxoAVTE49WNHjdtNMt0pcIV8sz1e
1UhbQ8nclU7L63/VW0aaQk1LfGfkHodg0tD0EvqRVw8KC+Am38SEUu1UMQjHyqhO
7AwyFE2O2HYxeGJQ3fId0apYET1PSaWJhR4KwuA9M7sryQf3MG2tQ2G3QfA0aQCB
dE8rRLi/X7Q7eGp/EQoGAmBjhM+Ey722UX3nVJiMPTW390PFpF6SUKp8yhvn9YES
jJszPNDleh9norZb6MVZBgQSKutgDV4Iz7aL/lRDhOLAY0U6pwA3iQ/j1qJQ9J2+
OZ4lA6xHARQTYnPz0NN5FHtnlHXYg7+66gHF12Hl+XXZcse3lY88LAKxQQNpd3YZ
x9jSGlbeGk0n0VByFKYQ3YePIKluAjyWp/J3r07c+1bIxCAejT2mLRYptSc5eYfQ
JZYf0iJ0d9nImNIxGLbndQt269ACFtQFzrxI/jg3DuOSuQXSYbxs0cQ4ynkYzS+t
Nz7pYEnYAkTmfG5i6sKcNQYI3+VcnzaZg6OewPFkOekNX9Hiig2rtNqZCYAkNmDt
IDvhBue5ClA/BFTSnjOSefxQ0aHVpEZrxBk5BdBHLuNWNRu2iVzA1xDUmVw6uo9O
6ZG5EtjhqC9fIFaq/8uLtIWGUTU30Dv6Y6u+FX/Eewvc3jWm8z1UfKnvB3Q5TuzI
oEB+ktPO0+8H7Ou6S4pd7sJICU7Sg+wJewhVzmJzrH/hJoiqEBi1LkEUYnGUfrk5
BkZJvqBLFGnDJAWNPci1rvsSp4JBx7/Ctcw3sdGqaADuH69HIbXyjXiN4e1YtNlv
mdI9hpmSKTq4tJt5+3jbkkrNd68+PamwmW3uLVAZ6mnSKoNDXAmKTCB95MO2IsGI
JGN4wVKdVULHJpvtsfjA9uvi0JVgOgEZcGAoFCs5KDNbFk3/BoRUhNu+ptjjrs1e
Ua0NI2I4prTSr6Bmb+o4NDPumqR1+e2d4qQD2rKGCCojISmRuTNeTiN1p9qFZvFa
N/mlYTUQ8X2WdgFncMzSiVMYJMV5sRFUTEbiDOE+gZ8mMKfwTL94JiJfhIrx7Fw5
blmqyw+Bh7sWF/uRYgc+IQOuf/ko3OUOucRcXGhSGgEnCl/ABH091wl4Vs7fv7Qu
Ujw7Rzv9KF0JCKEJh5t+tIbOp0EzJGf/qUQHRgQwrP6luYl32OOT9k15CTgzOpIy
rb0xCOt7hECOxApZ6t1ZHhvSvqjbrV1Y4sglX/DnVabCiONuM3FEltTvLvtWPU4u
qMkHI5LG+ruAhaZZns7U4Y460J+bMFiGgG33OCK3X4MBI4DBDyBQqhaUiWVeaCmL
opFMFudPdODSpobtTZNnxQx+iVskPzAdGAHFvMJ8QzzwViTFVZDJRStTO+8fRiG0
69Ugp1Ay1DQlGbyL38xwsoJnTiHM4KJg2FtDAp1/S0kL9D+TwkGE74XPkX18UNi/
ezL8XJWT6gkids2GjYuT3qS1GIyVy9tSiAe4pibs40VJGfg4q/E4ZktXQm/+XIOb
dpjz6jfYthJTbO2PNuKu0BgFiRTFuzDALMDBQS/AX4Pyw5KqbO2CrxPr7ylUccbF
ewjiY2xkt6Bqz6cviojKhXABJhNL/T1HaP8nm1sBrUwPFdNefajkgkGeCWUIzGBJ
8XF7wYp0aNCSv4b3kkUBQHN1n8YG4TW5cvnXArisM0ecqlvJIdyqokYBRqbRaWah
r6hWkrVygT56Th0A4rXiALTapFA8SuE4kYAiY8GDt7YNle8CThhRKIlFWUbFDpv+
xXh/HRRPIffUPug+IboPWT4rPgfyYx9VpHMMQFTMWWpj3882/ENKRWViSqA40J5M
q0QtR8MudYqyyw/tM1fqbgzB2o8PGd5MaP0dMCDMfdgO1dKBobCoIwZTQs71kf4K
28AAmRGoVNV/rAxYcv36S13OS2kCBK+ygDKVLoz6ztk/93Zbv9BVgf+0pNebgYG+
8m84fiEZ6RWfYwX1jCHodcPvTWscnureDEbE+HkFK/56+sAwN0QUmO4M8Zz6NcOa
5LHpzmOQJCclFeSwc/HDe5fr5mbF6a2+faQm8G9cC+aP4nqumA8cWy8hGhRcoqzh
7p6HuxkAGcD2UFETD6OuoyVExOyP6EfZpDFWp+Ug11Hfk9cLG/ZM/7Fxfi8SCl/g
VzmKZH14PqXsAc7qhO0/uXhX/zrnsoufsEInIfn9GiBiNnUojbA+lPcOjHvouV0a
p91q3BDeE6XhAO9tyLKrJ8hVeSKE6IxpjwYVnElDkY3X460Km2WIEdtgOqEA3kcu
LQIMFL24Kbq8ViismnIScUo0MD1/d0qB+u+HqD2oNs1fKkv4e316DY5t3aFc44IL
FGjVB0VVcv+UkqvKrs1nU/wfWDrFdEnf0bTxtNKN0BjIvU+/3PN3C/666Q5q0hs6
uOqfKl+1r4L1jNNczTQyLtWJrGrxuF33u9fOQ7kvdHYkT2axF2BPkKsB5Bi7uRvx
/zHsPCHVPZza4coR+LTmUfLwF5lcWs6kVK7KbnyCxOJYPE8jEGN0LjbWkiFMGMO3
XD2tCjCx1JQvhQfXRfK2MzYjazM/a/uHx1SBirXsD6oAaSC6HvDr6+bZ+7s/DrwN
hSH5ZrbgNScR3fnm/Jbn836orh58nQVZl4ebQRGV0E2DEv2wXdl1cOTU9SsDvpWM
XD/OSiP4hNDhXIW+mVQ2KAOpiPZdyXofLDM2b5R2WparTG+78URzkOIF88EGovuS
Vf/atiFnDOJHOh0X6EGl/0AzobDapWZl0AUhHcztnT1VytILukwpxcHlifaGtpCv
TLi+JssIKkl65vPf/+SZVj6hk3JrngsTz2AMf3uxzYJkof3luBcPTVDXagbmHvrL
WBLcIQbIZMkXjdo0XSuIV9n90+cDUPFeMKksMeTtmPtGODC+v5uDe3Ht/2AfOhVE
77YJ9NBOaKd1NA+TD7/oOizMVpKO45Z6YWg0dGu0KKO4DLymyYuI35v1IJbnBC2a
zyAuuFsvBGrBmtG1aB2Of7dNesWu2ZxrgD3FQt6wnjeD7qEia5yjMf6gnaDcWgMt
0eayIqxl+/gSuj8WyVCBVknWX2uFCv316AlB6VD48t90aUaLugxXpgb9+Ix4KgEX
c54stpg3RaxHv2cV/2nkuuBIbBFoRJiz4YEFziUzgzROgMa06wb2PFCXqXTKNXmF
QDx7sLkNnOZEWjthMg7T9yYwPccxwN4xjCDD0GUB+sPG2OZ2quT58oXDCB9yRmz+
7wvcsG1phfT7hmHP9bsy2NDKWL+5U96vWfrMYrdFlMdQr5Rm0ZJ7OFEivkElvNr2
QINwarA1URQGnBXVq3Ox32DI5XXBv2xlweuH4ZRFrx/X33BnQ4wwTFwIFpyvc9Sh
W3FlyzIhLN9pYMQrXwDNBY65kh2tGrYv5ul5n0INDZ0yfzSnFT8DDUEfXX+df4jQ
mesDQECO+ORwwUSr2VpLutviOtiYUKjDTwu2/rm3zWSWUv3Uceg1Mwcd8KGNYxYr
lWImuXqK4yxFxzvXzDj27DTFxaVIq4UbBgGdjY/zM4iJpFrNqqMTF8HAuXmzeux+
aqp0quUtujqj0gRJjnkqzHrJx6Lbi+qQ2ThQMDTPMHBUky7M4Gc0gHjQ/OYLloBC
1HgyZ4Ob8G5FsPsFwTKzts/nJ3/XKUt4M4sR2ynRwNSy3fXKFwcrsMEFANZVqwI6
bLOOqbfeCTa9xrQi8eoF9kZkdofwwuxv9ZuUCRw0Zxq0Z17/C3cUSw/l7Bvgj2pc
fU9GaPPk2Jmt6gUIiuRUNkI/4Lz/LManLsq8WbehUtyUSkos3qfzXYzM6RJds1Hu
jPecOPLSc0cKsiDNDqUDK9o2vrvKMEDTesnkW7ESys2ywfkSocj2BShhuMG6ONlW
SJjV6L2ffAzl3xZGl+VR3mZ1/JlTwUTVFdhzAum82mkmfhvSFkaDUDC4PZi2Hf57
/xe/lykyIYhYFvSLQa8bYaezi+MdaLkSZ84Uga5Nh/Hx1Ic/yIP47mgE3JcKgeZO
wns38cN647a//KO8dy7kDwz24vjBdlE2zZ0AeEpbS8wgsZPW4433RYIuFimhGWpB
/6y5CID/A7ha2g9vNTweqJm3yPMAJnb1Xsl8BtFXfT5A09wfuVgBgOtE5wbWUGht
OwWAFYD549poUe9jxXHCOE+oEx8W3CvMAZs9py3JPKVNa6WQy8iUwQz292Abl/Br
N6M9NWMsaemjP3fnwV5PuQkd9gdR/QhtAC5LLxZi/1/L3z4rnItzjmgKj3Co23hP
A1m7SLBY36Jat6Bmvi/XMPOuUMWymF3zeIEgd4euuGtdzYkzPftNXiX1+IILJj5c
7LocjuSeqsEgwczaPdMld0CSgDRKEE7qj/gkoWO8zy7KhJ5D8Aw80eBnIPlDnkCN
gQu0h0wYaCXcqJD+SZOWBxhjGEwUc5plR6v17dIrRkQ=
`pragma protect end_protected
