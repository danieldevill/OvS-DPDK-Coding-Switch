// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:04 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ItPPo5BqEwfWZQwYk58D6iaUQYnN9Wbn/hQOHaClLzpk8EPk0vMW3NKAG+aBH262
1CQfkvFXmPd/VHw8qWKVFMXOXTpvi1LXR/dqgYHz13oRw6pTM/LBCmVceHzOJSNb
xKccZ5CXhpM/tDJbD3RCHmw5108RpVr5Ev6bqm8syGM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3216)
vdgd6sAYNAuJforiyKAYv4MUQd1GLoM/4ZTj3Eqh/Mke7PyEKIRD7Vs6Y8jPFvFo
OsCJGp9AV1X0KswpMRDROE/4IcLJU89RDv6NI5CIlQVHSkMuSHq7RJJ0Ro8rM7QQ
+Ykq5jmhB8XUlrwpdDK26ON2KbUs8jMs0tph0QSmyrKmTPqGDFlZNqFztYEFtBMx
BRUnNWtLQvqcviiXzyH5y42cNivfdH7re0Q/NMj0onBw8if/Yd9Wk/WTtg5RlZt3
FpgQf2BNyWIreMre/dMrdopxo2P6rNh9FGC4xB8N4Zvsw+QwuPladKg0/gNsEmX9
fUxhdr/3BPkUUZ/g+ZvlGSGx0vP+MjxVeGDre6r6CKouGA4FhKFRUkVmMeZDkKuT
pLXJeTuLf+FVdWSNztceWgYZGzkH2MyBHKaVqLJHaYIkeznthD9/6JFDnGRmhOt7
l1BY/qVcGgAfr44epIIOsobckweyJH+hj6qqCaHF+FjjOpz8S/F6JdYTGj1f3VDZ
GkjK4XdfuabJOjQV4PmYmcJfaW5lKbTheulD6Akkz8oTwizErKGpf8qUM0sqdcfc
043MVfuDdYSP1qY2xkRAidKzUFyovPHCBoE6Yhd0OlSLUsAcG5Q8bucf2L4KJsAr
tfwIRHDeWg5io/eCJ2X6ME3qZMbX5lTNe4T7Bi0eZ5rJE0rklLdTVPA32d0274Xv
34rHkpGkf0DS/Q8/ExHTZ0Jbug9cQGQUeuRmqfavffki63tlnSw3RL4l+gW2BFS9
d6/1jF9t4ufI7lODlqmTszEopyyyxKc2JjZF7ZJnthDKEGBuSp+evXBA71/JAxaM
i1Jr1F+VR4JnoFxCnrpYr7fX7kWHt28XQSfUCN1TMGWgwqcx3c7LpmuoIJbLMG5W
AuOsLJa8I8m62PvssKM0nANRWnHOeegEkAcg2slkm4AauQE1z9VnU31t2MyfOkFo
by6xymiyvj7/Fd6MdtCIMI7ydIJsf7B2edHSWIOn7yh8DvkkXhODqE5mQkDa3e2b
lD9j6Ysbnl7NVxFakbR5EMlBqTGkk38ZvO/5k5ScJ85ok8U1f/e4Ylkv2DZTRO5v
Qx1XjzxK4t+ymhBnYcpH8Q8DInWoXtHSu5zVmhptdJ0HD3Ml0MXeviOqlcggsh6g
G4ofk/sTbUjNkIoHB8koAfyYp5YF74ffOHMhZqacQanN0c6VhR1v3LL1S/DGZVL2
wEvcIcP+QlzeN+S341qFht9yUmA30bM19TxI0FMwXoMA3rrwiMeJrTwsHWpYWj6p
emFko3BzOdsPY+7UMF1+/OlObrbMOV5IzwTcnN8Su9bl3poOAK2eRES+vjufQtw/
URFSZC7HeIU0apF6kEGYvaqiV18fZyg19HAlaYy4z8frLJHXDAdx41TG49lcpIYO
8xhhqvzQJgndFD2juCZ39gaXioYxw/mk5GT8CLoJGMgO/YMv8We6UfnfXlvpLFzk
R5vDKq6Appa/TsEJ0KqzMV7HhO8jvKDVeFmDJChSqNQw4aqEIq3KyKWL7AC0B4yF
qOE0YV1YcfowfXN+qNZ2PTGmLqL69vofi7QcZpfp9ibAM4EcL/6XYl5TUnLyFpRH
EXFor1SPiG+gk6Jqjkenyofur96CK5Vtbury+2jw/W8oTRmRnd7DLBuGEw03yKnD
rE4zWgo4lGNITax7+2xfLyqv5q9lx2TXRuhvXEwER5NnDnzs2obU579jFxzIvTKy
BGkZ9dzGItjFF5rNu4xqoSjIo7Uf+xiPRUtgIaklCXsSHk8lm+jIqK9RYLajJwKQ
L9vyUI3T/kAKrhTIDM7W3ifTO46CAHcb4IMK+K2u538QsmMrJ0z1Jo0VL+45MIZp
9yqMLUWYbl0/E+iLMvlXpaFkF4dNMZdrWnZZB9ffpISkeG+3HZ0DBNb8Pu5SDim9
zTxKH+2KOGvSPHLBjb+HRn5EwgimwdBEsiRrc1v6t3cHEWhEPLMT6AjjeUWM129N
bB8TaxJDlhsTTeH2CQZt98i/kFbgfcOMqK96AIafuF5JSN9svHmYFJLCgEKYz68n
x5e5J6s8AinZ646OszousUR0bAsA2YPEI8W3Dsiwl6e03/Izs/KOx5PXt1CreGSf
ceBNAvabn4R0n7FaKV9R9+pjweCad8TcJMIZUHjHhYJU3cNtcXtPSXDr4iyHAr9K
cz+02DejWXDELfOWQHvc9WtImc3Gnt8g+D5mlEMxvpq+JgIuaMqawWY7GEWWu1nt
OUb3hxqQxq4/9DQxyMuiTZSqrl1afgZwpwHksc93dJYU82Nk/Iv8YW2snu+zCxl4
oB4X0gY780LR59mLnAj9FfNHxupltU7TZcWmSQmy7AbLoB1BbwYRuxQfetxhGljO
0xZaklaHJHQvCULzaz2YGez7Mrnv+kSUib3KD8owfWrGrlLRo0pTd21+Sv9rydeX
T9UQQ/jqIf32hOEUdQmfHIdj57dFShpi2SxPTrrhr339cC4RhKBzxr990eORU31n
3EwQ4PwPi5jlO/NTDoeen8hwfK/PmYDEXpkfzaw2izji6gCm1IKW6XHvjRRnKuZH
2awpcNTTypXBfffD9OYZo7937E8BU4GuNW7u/Kq6uC7wMU26K2HTnenpOQlvkvQt
Zpapqi+sbHER9fcEF8DuJmCN/hSzvgz1ENougLOf/B2+eaf1BxsYYizCsW6d7xJq
P4pdQDP4dg613oCtmQMBTuXaNFqRIgEdCI3w6FDu7KfHFRWDSdT0FygxUQKkwKsV
eEsa6hnBrl9+AORaBmYRtXIZc6eS5QXs7I//w4HTQQLUXfYD3BQEcT1JiHqH+EOo
PdXNub+kyswm8VsrNRZQ7xZDj5QcjgY1pB3sMI2LDv7bnkfkD3JuZfvFCTjmEIyX
1tdzi/7KPwh1/mijUOQNqHF7SkBUbnwcm5H+bNAm48fmfq9PaDdVfzPW+F6yIIhf
xADaZuX7qyPOBK0RNlRgbX1e2Mf1It8X6BVbs3pj3qOM2MpJT0XAVxI2m7umK4++
HDHShsJVk9jMDhFRKryVU23OZCYc8cPh5auRE9Q4ENMqW+dVTi2AzxtAffZGnjSG
3mgbok9OjKDSMqRwkv64VCjiv+paXdjNK0xgM7QQqUKCSLbYCw8/iFbgbBxxudnG
snFRFNcmTK5AahvTGOBtsbJp3wEeoZxZis6muzM3JQVjrNyaHBAJtZdd85UDFQxf
h4RU/YXr6/oDH019KyWXlvrTHh3bObu2gTN7yggPUvhpz+6DlDJ4cEupeVtajifo
Gp+e98eM069kGqqk5WBGSnjh5oM/okcds7xjuZcaR2dBRhzLMRqf4eOvCqk1rfcQ
GXr8nsLntVVcQ1FRsl2ldn2/eemDhvuBosp1ynswU8KlWRAl1u1Az9NGb6lYNNK0
FvEVrW19/c/j79mozbzHPMIAyln15C9ONwm7RcJJY8RvPM1XSfubPIJDXUrh1iMC
iNq9QGxqLt6Vmsc7AD1Dgwwv4PPvIVRY/LYbsUya6TKIiz7nafiRzMQuSfyo2j4b
cd88dkgd4arA7V1ADat/jdupvaOdaGY54F+ot5BGCmvzjmBLXO+ddxSzKTGxdBC+
/UcXnYs6AKXiKa36bj0OxpS0Us+hdvtKYxpIftyf80uoLWAZMW9Myaug135OBYB+
OxpnKO8/8kZg/O0LnxQTXv+Md5/9kJFK1i8lOY9KsBvVYTn4UTLZ80bG66NNPVpT
rB6cbt5R0CovIiJ+u9RqVwFDrFUsNbv09zDBlZs9E+Zzyown/9HR2A3DC2SBfOsB
bOVt8BBxGp+ey2ROQZ6sbNxZ/mCPeBkcZb2uN4XlMsf9WCDluNP9IjpF6l+OPkdS
8xx6IUZ50lEIuUZrQhCP9L78ilvoT3qCEnJ/jyd22zzZd1Buhin41eXbHv0WE3M3
2dybohjIlQ3KmCzFOdNEjElSV5r19W+sTdl93CJzug9ePBDd4wNv1LyGfLpBInGf
4MmjECOsFfi+Cukn6e4GWoRHceztqC6GEHFgjCe5jC/vxKFavjLvtm9J55kDZX6z
B3YyoPgKD+9d0QNA5OMuD9rezgl4IhxGDErirwWel0Z/waHGA2+aJfECrZ2vb8T3
notI1mKvs1+FEjnxx1eOA2DGzyfDsWH9NmzC53KMhIijgNVWXhiEFLyWc9SqLawq
biqccyDbX50b3nulaNSvQoeHKdntLU3GAf15yU/mTUarTfjYzol+Rjx0yvFtyg/u
jfziCO/EHw0B8V0dpalTwaoXBDYg8gKbZ1P8I8I5nQ2r0o2jiu4qfTxFcgyuz3FA
`pragma protect end_protected
