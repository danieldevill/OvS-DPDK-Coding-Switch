// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:34:50 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WucOx7SZWTCefqBJl0rLAEHLpYBG9VpVMn3T1TlIy/DSRbFpqdmawBsvsFlcFxvx
XdVdQoL0eVOQOtw9zYV+FFEMdSLXuc56bn8PmvDB1QYsRkCNBUCTOJyX/EG5FI0H
JS4qqK8d5BG0VC4dAbAAf3XdrMO5S2cAIjJ3XKnhJJY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 41376)
bfZ7dWNLQxNH+UjOZKwRXnZ2rsqX6R0X7jv78mf25b1pkb6dLargK0dJDKq+qm4B
H4SNccT18MWYcBXlP9ubLWxXtViyOVfAFqqXgcJZhurLwN29Rc3iGab3uQBoITcF
7aO0WO/BZWwD/CXmviGHL3lVTxAyjYrYPTqpSoKBYVSBKKFeyFkk7BDaeW69Pg1B
ull3OgEwmDjdJ6YDrE0yCPCWsh/pD6kbdw8DrO9B/3MaGMtgSGyY/vOc5B6Thii4
ynI6SYJUignydDv5iXPIgfh9E7uP9kSFl0h4rqLOp1uUX1RGrMTszPou1TeRKBaT
FKjV5D/9w3gQ6PNZBbzDSQgf8R4aRslsU4YCJ2O9dLsMoLbBrtd/4uI0KZRBXI6M
vjWv6VCfBT3ICUO3GGclJKe2hYU5hO82rorXwDyZb6Lf4zoNc1ZtZ7Pl8SihsT9r
9sXulEBi8+E3LJhH5f3ZOss8MFph6AY/r5IshvkwdqrmZv/VhlRNqXre/4+fuApp
mtGVR1BJHHPFG+WKZbHmp764sj+SqE9aMzz1lF4ZSzszb4sr9VONk3641S664CCb
cPXCXTLiatkW45MYanG1xcU4/a+0HA/CizvpQsxY6kb/PGOMDHUfOzrD4bVozvyy
MeoYBiEs8pBYGmVyR+5HzNA3ZJdkYT3kYf+yk5yfsI+oJamsoLGbVW1u61sxIguo
2snI+FRTlq0ULkIG5td3niqtZI7S1VipcnDpJGsRai2jmhLSQzPj5DAKS7psmSc2
+WrKA/DctWaZAoDJSSXce453qOIqamCi63T2gaVVNU+iRkix+hSb7dHXRZDb5WyW
BngAdtN8uwQT95GzPQCDlhs3H7uNZG5NUEgzLZALzT1ujUpYtQwqSWXXPWumVsPS
53UOEqJke236bGMlKc3Trl4c6EdOLGkfRiSfVwomsYt1gUF9YnQs34wARi5tCysb
/2zat46V2Fst+H92HFba83DDvuYxNqpdQoheXx6NdW9XIeKfcBzoxSvE7NOd/ZWq
929YZto5l5G0Eqx5S7AWFuieYLtBGbU/riSCBjnGM4igwwK+Ozk/b/qHBofyNFNM
4Je/s2NoitrC505WmCJXM/F0DfSIZ8znqGmabPe5xnWDjnGGFGMe6u1Ktbx2v90e
RuAAcn1kK71HrYwTxUb1hdHYEiKoyKjquHjSegHOUcTPGJmP70HbEQ89a+K/8CCP
Q7ltrsTuOM8gmO4iz+vwpt9W1iTy3xjbaQzjaDYUjT5CLYQCi7ZogH2ggSs6QyV+
OlXXT3ygPJz80mbjc8VVF54YEOabvTbRkpwhLlIDPx+jHxjhtyUOo5Mp2PJmn/3p
jUx6hHdcr/JkC5VUunh7MoprySxN7o6LCujYiJyRp0lh2DY2a4rA7myHQARBrdQE
YmzVVc4bySYp9C9jahiY8++aEd65h7m2iv8DBG7QPmjOoIgZF/l7QpZ4hlVaxYHn
GS1EyzfGMyW2WlxPKM2KFB1NrUA39ZEMXYV9vvvxXB/3lv+vAFhmGGlL/4D8/+CS
gXVV54D2UUlXf9cB7dPuaPSHLAw/GIWVC2HY+/fyFw7MX7OYfarJnw+EUufmIDSc
R0KjbAPfTyEunRuj2pbFi00gIx6/6Zuxst4qva0hg+wtSRbFpiGO9nuMpUllvCAY
CSL89AqkxjV99T7PSURZ/P+K37dx2ReglDP0JoRxQ8Ua9mY80IDHk0Mt3xAx8sK9
KKB3IYWPZJEAG/fFl/T1x0vyT/mlswV8FVkHjeVtjHNgovt45itVOVEy9fjo29nO
0uYooYU9dDTduV3D670wiy+xqu0ilS2YZADTTRcpR59WPWWFKLCTUuawrOGaCZhO
7Q8Pfp6uB0c9NsL7Z5HcVS8uhY8otzIRnbof/EBBZ7IZ4q1+AAR2tjRdpwzhhjCh
OvwmSu5LJN82v672DuqD9KhDdCXfgma3NT7If1nJJ+Yp6Al9FBHb6oVmGA3T7aFs
WzIdYfcDP4NYs5hSAEh1FFK+ntoBdW16EvmQD4gJOBkD3c53JsmYQpQoLGS4kq2D
6YSMkgK2+rNdoTrFpQkiUVsO77dtm4krcod4S/EKQqydnGMEYhJZw8c03svBzl6Y
tfYKl4fuUNYbxas1VgPKsilia0kt/e5vcEKopYrpHIUFl9fu6glaU2t4qVVOk41t
5D63sifa/xZLHRV0giTYJfZvo0LHTb6hkJDdimDbEx6ogPmqT0onHEBbVcahUTig
g/PPF5o/LCc6dMtShw9CWfVpjecUwOW2rLi4YWjVApHri1c4ovIgHeLRa23wtjFT
5uS41Nqdu7xB+XWBvwN+AbWizHZAK8w6KMmxXDNwv+WHacRdBWvJLKj0UdV2FAxN
hty7n3bydPhi7LRY2wX98bscNuJ4Ii8fHHhyQbEu+FQoqkpNQalE/fU+I9ZyrhZS
W9u8VLk+JEuM29OtCvhE9lix8+TioreqNVV2J1zApFZnK2ng7fA20RFkWofXvdFC
GQv2MgbKANJ3cvNj1ChPeTfojXeKzJY/lWE8IhkB0yPOyzjPrSt1cMMBC1k0EQ+8
BYJ1DZhBAOgsJLj3vYJo93M4a8RUrBksY5Y1gOme8k+1kxyq4F26l8M1nkNZyUoN
y+GdvcAsN3r2SX6pgK6HvOi7DWsTBCEaMk4nv0zdU24ursMGa5f7wuSE4JNwSvoZ
o1p6+MgTAb8ZcBGYMyGQlUzNa/PJOsCzhp8dyyUkj15G6YK/xGyUjtYNGfwAFGGq
E+bjY+46uRqcZ6KuLFZLmY0BRPeygwVxELo73/At+Vjg3kf+KSxOrdt5YYAsIRG+
zxZZoX4ESjXARposIYpF+rprlUcpGZluASpRgzgHp6s7RWxAtf02DNghcvlWFDYU
y78GV2q9zqozz/pYJUq7DExCCQnz7NMBgLY0pa2WpuzF0Rz/Wbs/4YRNxI3QWSaq
YY2ASs1s4tqor7D8VFULpka2fjaN9CaCE/pFQPHn757Y8CICVjpq7Scs6c6oyjp9
VVOfmBoJDYAqUIMfAFsluy0NcBzHIsdlFKRoi8PjokCjnjFYqpoWXzJtNK8B0Ky3
hsC8V96c1Msof3iSQccfNzQDqZTmh7yxP1TEsHsRTPjqa73/W+KMZAH/NJWEazh9
zj5o7SH3v0TGs07+SWCl3vMXpg1wSh0BV/f+7acksyCeh/Yfq9oiAUV8bqg8RGDK
mXRSSfOIL7PE7f3WDmwNlp0DGns3daDSAtzERiatFs938XX1x191azQuK+ZxwHfR
mCt4EsemSaCFWZBSWSmQdIrvn1wt8kYvnpbK0jsIScBhAUhJc+g4CuvJGA3ecE20
ULck5mR94yGN37AYfX+1lBMGN5h3xCy3za6Xn5QImrGlah86DMOFb+adbbA/0jn2
oAdO3B6tiLVhOC+2jmaSH+85aJ4n8yvsXaA95nOI0TLQq0Fxh/Mrz1puHD84AOAl
cy4wxUnbVGQaphxWmOmKpam8W2+/88ooQKlS5nKF75SZNmCaPXAOeKmW3R9Mzd/1
P8V4VL7t3Nx52xk5i4kVgAcSdoqQbYhZuKwSrCV+XN+FslIwTogD546lqguRBA2g
iTNN/bYEnLrl68bJESzEBIWSIAdhAcmqjLWe80Z9AaeVyB+ux5B9t8TU53WEjmKA
dMVTj1t8M20lDZK9A4xbjwGdIFvKkiSLubyCx7LZGmvu0Xy4NuWbqVX7F7EjwStv
e42hB6nB8rLEOw4CxoNNsZ1gEAkw7Da+NotxBPnIQJoLcoQcteVfAY5GSLTQg3eV
mBbUzr/NHvYtTfL1OHQR2KCQygep3u4aWnTnM/PCUuKlMU/+EDq5YKb456KvpDm2
JutW5xVHy8PSweD/pKG6OZ+omrIrFLGsngRKzALXSY+sepaag90hdNwlnTBHJdmK
R580n2NCjHpjeHOkzsNeydusSdZjCNkjDXHQtgfY807Vx2o2bNAVAZ2vH4XaBrbh
A/HA1tbRZtuX6dTgI9l7kNgb3rfaicEk9mhapMBKUe0WKwv2crxkAjmXqc6x8IyI
HGUtJs/SXdGaafZl4yzWnK64HyWajLlkIU1gmirKlovQOAz4g2DLrA2oqYR+akIb
Ewdaz3UpZo/PsCxeHapP2NKz5FLWaSW9i7JH0TA/Sd9T/dZUt8nVk0w2Rhi0wLC+
6Puj1z/GjZcaHqUTfuuthCMeicCZEPc/pCnTcLU9g1z5UBqkt9EnViOS+gUpna7l
X4QLbffNHJD+GHk7VfdtOHGPgxqiW/AqLRy6XMCbxowOBx9Envme6mn5gzGOfzpf
WJKynumFK/iCjx7vb9hraU0gLtQaqAFwKeFH2OpMSb4WTYvRFe2aj49nROZzG3ha
BL+wPSnwqz1RZ/FhiqVAnb56mKPihw8kEusoIVKZWR3yUwaB0XENpb7yszKG9egq
SnqIXzXWbwSEC5W/F90AO8NO3Vq1Gb2Rmqk1SEiF6BWeZZgYkfCWUGKqTqfATUBb
Aa+FBckQNCR3/I8j8XrqX6Zlnx1kEL10BQhXEbapQMMxwxNGGhrqK32+3+1jEOls
d+/BAXreARUGggwGbB3JcAAuXm72Bss2+2E8+aaJpAsZ0r4YRpKy1cAOQbXe9Cad
IfFzWHCNWmwED1w4uJ+MxzEytavx/79JqgFKH3QpEby/gA4rpFLOj6M3W/zJIl1T
K6IGwSavnGdt6dW3vzoEZDLcZdPa6bV8dimzDUuniQlzUz1HzSlzQsHcz06mOAgH
211aF1WLktv1lNAyaoyc0Zo2dxbl1+P/bLNOh7SzTQEzMqecea64vyNMt1c4JAIC
rlUoQrY9Dkhz7oBJ6FdmI9cFMtk4Oh+tzVKvNSwkkQDEL8BENagfPA3ONzxfBSGQ
OOsq/6lOs9xUZV+sIR4U2WdI6LVjrScwtfyjaSPnWFdzyRQc79Hxx4dxbEoW+rXw
jyp+Oqd1KAno6gEFJ6p0k1GcUoGVBawP/TKWEPUH1ukc+Y8dbqr9f1DG7FWH/581
Fdnvx+m8NOpZFgZpV4YGlevZIXamSue24pMoxQBylhaM3BKZ2JTlusJcUM9qKobF
4F6w2PKBOchNM9ZVll50ptDnpYW5U+SqnEk4nPtohVFixGmUAWOicCmQjtP5S0rY
922km5egxnsgkKz05N7nEVPtUvQ/gjhbJpdE/JW9gcJvPSlKmmMqc49ZvpqigqTd
eAYcKqL8PFaygjqFQ5yRnHPw2OdGdpV1wh9yUWs6cnaDgS7Som2m7D8yW2BonlPU
1eKSS7J+OH+FYpmfT0pTlFsNjxi9EL09mkS/Rqb2oIZ4N5NeW2OfwhjLflEiJMsS
p9kN7DEQr4mN+NOkWZKxw5uI6jn31eQYSDfcSua7Ry2YO82PypTaigr9FR3NfmlS
B6cAADAeseY0U5Sf0M//p34omTB6j9Xm8gZoKd1yxnAaifMT9/+2kjtPN5eWePEs
ixyfzj9TnvMH40DpaYPvEkivXGV6uU7W4jYk7OzZv1LFmn0eIJaYB/CY8p9wPod+
0lFby1BQ6CGENFblL2YnNCvUrllEjIA0wcAoggltG6D3Ooqa4IcVJsyEa1o+v/rz
N83/T9z2dJUvieRmkFElvbL91Y+2XeQ3++6glIgSUQZkG6XNf90ssV3J3bRmRkTF
qykz9Q5dSEq0sbLiNmQtlpx9FSVDLyiuCH30+3ZdSMifHRZJDlVEgKWqzVmSicQ1
Q7dlcFllWbg+eSuwQdiyq1XzORrCR8uHwtc+TkyRnwHHILl7eQt/oGknSt9kXgqv
ZbPdnQX6VHachqROS+J7oUx6q/iobquDiB0evrjvU8fXjxw9Mz/qtNFlpgn28VlE
aR2iFV0imsbTr6O3yPRj5tG3vCrHSByiDb8h+lS9q/95B4JA3oRDWxkHlt7DYEDe
fZx8UulK9YLu2zDV2Gl6ARmOJU0o/vaGqesWmrdeWKI8rDEngK9pqhiNwqD3FZES
ywKRUMxaXbYPBrhb/6HJWWHFgh152BaA1g1b02qmI+oRjdcCbQmSU3u2CKqK/TNR
2gUpw0MQNH/cFWfEvtDJ705vcE157k/8FAxxU4u7QJ5hgqboSQSa4crJrPCvd0KI
+7ekXRp2ytrKvnqJE3Uqc4jYKSdvBmsteQdYhcfsbeU5i71mwCln6LQ6aCPIJiI/
PdSV8ScdxjkBEW/sFue16+nOsF6l8PTlHYw9JxKtEaV+fuV5pUOpIqXSJXLp1ToT
Ch6UzY56HCJRjat73q5ySueTi4Qv+lGpK1GCpLSS/WW9MlDlRDEUSyQbwrvynX0O
EhAdWeCEM2WB4Z5tctPTJfhhxaf+Xy4wsvk6MuLRoVvWO/Xd72wK0GevPAbvBcWm
rktghtKvDxfELYyU7uNlHI9aDbuGRuiCVDEKi/QenmwzKK7Rif6dCy90/G9tdoXj
tgTsd3jkTrFJ7nuByu441/FjqL5CZ9rZcv/iRsVCRgqLAkvQ7qOEF9JTdypd8Csg
4R9l1DyVrIohIvQ2/VVThe4ch6LjpBAUwJxhZSn1r1YB/Toi7Qxm65wyElRLoVJq
VBzHbn33YVoq2k6PBF0hBGSVP5nYKh83cNmoHzyUIKTKTCmg/N+tIuq/ZLcsDu0O
8tQKl+4ThBhe7yyNy5ol/68MOkh4XvaVAJu/nC3x13fnGjgp0xJrE0VNGUzZ4I08
aHx6r6zWZr7k4twTfo6Kuxs6d4PdVXw9fziyWzveEoGwDeU6ysP07pykmWlK7Sql
+6oKdYFmeiq1sTyQYwXLNpGXE6q+MPHufFEi4v5S3cn2bkwFH0ah0CSKc6KhHh1+
T8qO4Dk9682aIIcQl9kSc8iPPxRb/p73PCxe3yZQNbm0+im1nid8pExeW16j1Qnz
zqloA2RDvTGbAbXJovaTByc5N12IMi8N3qfEkxOaNaeTO1p17EjgHb2IfCw08Zp5
yZPisLVy22aLy2TGFv+IECbw3ckAhGYp1jov5LMnIdfWURPDuXKzoopakolvH1AA
LI45EF1eyucFVfmXbtsHcb+r6YVqHBQSSiMdkrdQF+2OdKBOrW5JbK0NXfDinGFA
XR6ghx4yZEwMT9dhPi+ic5ANnZAcuBvUauk3hAhKV1vAGETjgsFw7VnF6mJntTYd
3Mi3l03fon58kE+n/RyqeKHpazpIVHvA8v3pRQQ5NSSwoOkkfB7IsuBOUg0eRsCE
hbvdgS7AmjIpeCKr30MLu94knkgamMOvj5Zb57HZCyfuI6KQTeFXCxdzv8fbXYQD
SrBA4Ys6GOJnQ0IryawATAThXK8UBy19BtV2LM1urabmTmA0gfI23gOEyjL2RTUB
6JsIDFJw38uve4mN6RxjHoZC74R5l67GzGL8Om8bIlyyIlclr6Gz1sWxWHXvFzd+
/JEmtOGHDu7u+22J+hUPE9OO6l8jX9hBYulMgdqo9J4J4xqt8RlzvISpUHw6tmVo
joYgvMTn8BUDf+vEJGD0sBpMhE7g5u7FbTBIeyfBToVnJWkymYADzzL/JNmXFqLz
P17ifzVvcR2XnirArkVAqxPKCp8eFJru43/sWYS3moLOUpRROFP+zjyAnlSqkagT
UXxZlJcoUm1sD/edkDHZeIDI1I3nhx8BvNWOn4WYBDObvGPF7EARgoA+kJRarEMF
yGqIjd+L0A1z/TlJd7Lmwhs66an1Eo1M+gtkiJa/Jxb+IqNbeMs6BmeEOY8vSPLw
jdqXI4L3yZ0ymFs62uIo3bxSEx+OUEj3XZoITy7wI3NE/SUwIrfSKQSB7ap+uf0T
NQxEoWL2bAsGwABH7qj8+7DC3is8vO1ABXjLUZVwtaAPg7SVVr0cjrInT9oOa4VM
ZezmA+V0VRWtxuR8M8grpqxc5Jo324U4d8BhLXec3XElrETve4pYuAu9kteeJqpN
fcyUweu+xIXJtyY2F/31/qqUvTJ8n57HsZ8ee9Nshj3Em621+4POi381Fepp8s4z
uavfYMlX3AFqmpAZtkBqwEV3LNv8r9GsJVEbv8asZ38ohCY2CaX8gyw+5Bjq+gWN
GhgdhiUY2Ik89C+lztBLD/8cAedd2OAn1qX2OCzI09DZV5iKz+HUYwvJVfbbPsjz
ejG4B0VSlYHCzuWfZjJdE95NRl1Dqqv+QjzwdbqujLTaiO6DvZGN+eLJXndbLqat
nNdssCDApj61SSYOH1iAJGJZLd5N7apLknZfSAgzkSoSp7ZlGvvG+an7/ghIsI0k
AisytEqVYkFLDVSLC58FLIvXu+4xWgFDFq8JPwRugyxHSuXjeZpo9GAXTPQHZs4R
H1uRMbqawMKvuRD8GsxWMW68i2LwosNH7h7HVgovCA1QApxWx0GKO7uf9qoyYoBx
+kNCy1cqbZ3Jvd9Fi/89MKdC5NUS5MfW1eA/mKA5o1uSRUQswY9nuIvLVnjS534H
qgyrjNsSCUM2SuvygHCv/NWcjtFLwwkYNPau3LNjsLkoQIOQCMeW9uY1/4tUIHcM
JAKmXiRbTR0H4zeAAWjDd/SNuFnGQFphMKW5dckuLQKHObNfgj1W9yLlDUn4gRp6
z2ZjOBiSjrzwAfyPNPv2eqZvBBByDg89uJl52Du47rnUOhW+Xr0k72xZGeqmBh36
ehTfmmqcMTufvvVP/OY16jGxfjPHXULkloji1KbH6p8xeUUVFn16LIWCSjkE4SKn
GE1BXsaaE3K0+cg0w/1Vx4z6QuXYA16xJdYqbK/ywP3ZajTu/GXijfIgSBBCUA7r
5aRaVbCdPobtnh0T6ThcCzQL9Zbx/XbF31XSG8NKCy7uL8hRB+jlbUbhGELhwEPJ
p0Vpff/m1vCWstU+dePfaHGoK5LyR1yAuHvZGBOs+CMhZCZ1NLGDXDF5o/fLAYtX
kukzw/hk/oEVVSVdKvx4YMROO5wBkYFG0UIMFIVqvCEnkN1PJeCUNP0+uJXsWTSW
0zcF36ZW4QnmAB5igr5VYxLq43unoJXSlrj+LSDXtgZF91f4PrT1CHXcOr+wub2e
0tCGyt/Mi1q9DI2fDCJHlcwKgWY89IAfVZLk26sQTt6h8Q/CekHbw0aBWoJCafoy
tAOSGsBHQvn8sWY1DdC5JrsmTfAISXwxOcGDdlEqiivQUOatlbC0E0In4IWXjYx9
64MGZBjdKuDDOPc/ZX3S1XWYAIjMioqjg/UclWVm4cBt1sIb3d+sI3scqAzUZZ2O
q5qYltdmK6As0Kwy9hM1l3oqc/6dNg88lrsBP0dOvjoMtBTpztEwNHxjJ3Ymdwfk
tpKe5pFSUFb3yVwXBMmwjbbEaMCPiT5OVZ5BOEhK5nV1L82Yjf8j2rt5YcMEWWmM
u4b5r3TbR1Ct9ZWWJl3SMOPK3oili9LAV6TTiFOfiliPW303uGANs0MUcUTLBIGO
1hEbWLG0cMqVhp70pPKs3Dh5Dfme85iGGG4cP6wDZur1xowSxdD2SrYojPeU3BzA
mS8CoQaX4A3+UDjxJsjHeUH7fW8DgUiskshltVqMdC2dBHqYlxCB56k0IaXu86hA
5h7s6Q6jcqI0SOgjyDfiOOGK5I6PdYUrxMsYgw5mZIkMUWo3QTfYgvMukWqa/Pnl
ePpjUcfMUVNgipxojFHMgHXk+XjlNhyjaJhmsQ+kHs+2MZNAa3vc3p/4ERlnklJL
KGQRm9QZfrWtAKbXQ2OreVLNTEK2anLk97U/y6iV+Ng7y5LLdqVbJLBjYO3AIB17
tX27IANx8ks3okWVDwMeAGJrHZzLINtLlWmw+qwtwizcASFRXIE88e8goo5PA66z
UPAAFLXIBRuEiOWpC6/2HjI9wC0hqVfD05+Uk4heD+gJtzoV7upNCkzrfmrE3GoX
qatKufPbgUW9prOKEIarGuCSYvUpiWqXUfDkoor/0fp5J20AW+kJ+OvN/t5cdNeW
1uEBQZZdl/NpHu02OLf8Z/tB5G9HLDkEDZ1fK/77Oqf91gjBB8GgrXax6AsmxVfb
KjAxf8HHknA4sk30GVtk+rPJAyy1TDccpB0d6LIm2aPQ0pQ2cXIavDpbtD4e9i+Q
ZrKiTmUPB2Z4fZO9VV2eLP994oJ3ScY/aKR453KVLae6/DwGg5qwVomWz1L0Vclp
spmEZv0jnPlI37pvRE/yWxIct+upZ6Y0yIipmRfNN/9+rtZmLzWKLc1NUQh60pCe
OEHQc5GnWUrliCp20LBusgZ3cy5DqnrHTMUvRwkZIGwzcRoAdORm1K1rHQ0VLA4b
uq+2K45JuOTLlnei3w5BDcWHmG44UKD4SYNEUWtguohVuDlsRpWTet+jDzN6nPj6
GVebIJItHzNBdB2jXKnUbTgV79jK1clXq5m3bqlE9dHSy2X2bHfyC1aPX7sTdTym
zGyQ6pQTtOqts16qit65bH4K7a2bMpmMn/6yI3uzKoamMxFuFlxML3gLuVD5UFWv
eFp3ALZnJ7zNczosvZ3cYzMw5aKpVH+lu55HZ29+Q9mTSOoz4erhZ5SBBIkeXJoC
hbIGFrDEU3g2iLt+C08aVGUSUWsNdiTxDulE/Bd1B8/Kf5Mp3bHOKvdWVnS+5mzr
/zEE5J/uP0eYhKDM8VuIsG68xNDWvLAHFLzeCmvCeCUakALh3UqhadviqWd7hyX2
TeRpuoDqqd9n/VWKEXcBUbKobWuZEROQA+eo6DXQpRsNWt/1cth8XL2jZ5oQnb4B
g76o12Dhnu6Z9OIpuIVDMMf0lXRNzdoxGqTvb5K2cEcAzyyOvkkeDDS60cD2rlHQ
bjvCEOCzS20/ERybl7XDJ4I0KR37z81P/AZkSQM2Hgl0uiKAZ8VsxyHOpKiQo5NR
U4ot9JDcAV7R9Ms6NQvbRT9UgNgz1WZuLPo+SSbWjSgthVUP0TRkJcx5sAyYJ8uL
0xYxAviz0enoD9S3Csl1i1HpufSuTJiJBxTQ1Z1tuSk59odpg2ilTrVB/7ocOgUn
cWSYGLBZIBQ8uUQvwnYUxMncT05Cf4S4f5CZuzVBRuqoGuHvBi348V3SuGYrA2RN
EH9Vt8PW1sIa6x3kAdT/qJnF1MYQPN78OpsRhUUVnRAJP1Ffoc+/wWlvEiJ9+nHd
Ynzfpb98IuDM/Yv4nvlWgksSKYnsjDEpFSuEOwaQt6jy8TN3FUF3gf3XxrxWaElp
D7YwuptrvgdSk2ibVgQwKJV0opLWIHv9A6uUku3Is3AfeCeBKaeLl90xAUFK751/
ps4QqWxSvZ/5QzRWaxgUal/PRVCvcUmCwJiTANhVPqB23/MB6OpBUmSmlZzOJHgg
KDcD6Bpg/dA/YoNlVG3Z0/r+h3rHe3e2760UZ+bFHom5zuPYZdDBpPagj6cNz2YS
mSjsvuo1HbhR0zo71AIdsnfKowo10Eq+OOjoDieKqWtseQcMqzw6Vbv9tQ0geiq3
e/zX2yJqLs0mzE8J6g8Q3yzLuKv/RQwPXeHalNoSOo9G2Sa6FqwZ0iyq47AAFF6R
HU75CGF77qe/ZzPdtLv3qkOuVqGgUQ3lSKNMoYZsu5BefUlukFVpANw7CuL5QB8a
EZ9Mwl04LvkknHc9I2neE9vP30Fw1uYYfmE6xeKl1osPLxhE30Ckv41pDOB7GfkY
IYNMRYuVxo1A+HQhrkdBG9mrh552K+WRYch1KPeJCc1w4cfwN8W2dsne/itEO4uP
7MK/Q7qfP75DrJfcCqx9LXoJHK+vq8t5FnM1k5n8mna9bucmaB6/890q3yLQ8+kj
WkgJH6yJaOjluuUc7zVjT8oBSsW7Cw/BnCEmp9D5RyFeGzWKILoBImAxa4YgqjS3
26LcPfno7I+cF3gE7QsqO4FklaSHa15cMuSEe8H7i+GYZSzgMweHTHsgdpXaLjur
FeBbT/4lJyFjd+Q+5NmjMYLmF0z+vP/G8DXBAyPDuLEt9P+uA5dkFTNP+L1J4Ytc
jhk6tXOlSAsAP3XGzc+8iyo0qG+OoelJ/2Z8NqlZVPfxZye/wZX1j2v25ZgMtyOw
+Jn7sqfpKX1KUDLljBeDI5X0NZbTPymamyMx+2McVb/yjYdKl/oTmbR3x2n7mvX3
88F1fOEvMi9YlLCVaJVxJ4gvH0s0KKRmKCAlTZTFgcBpYDbk9lEUjGCfG5h7Uidi
aHLhnleGPtYFFU+a2NNQQmhMeCNiIFSFSIZ86VAg5d/0SnBeZSxEL/kY0FCHor97
cGcBFz3YSV4cdCTqjo8afA6+l0pgEg8PanaOpH5AwzwQtAsjnIdBzxaac/w/nVMA
Id75msFuAjxPu2/8hvvSU++5jm8tQi8PNU84vu+JU3GYo3oelHHp4z+N8g8C2rTn
7pwtEauC/9T736vuKYEg6KogUoet6VIYw2jnd/u9jRM4oZz6B4AnElCLc84BEd+N
Nw6zPqLZkBjt9lB/DO/8Ewt8YMdznNxIr96kWC9k8G4uulGQ+55Rg80V+FlCsb4E
yk2btIUycbYW+itUWkEKb1Bv7PTC6DBJehmHAt6GZ1zJcLP7eR4fwEhpYAcCJP4H
8j64gpxBTwWK1I4FCWr6Go5bEg9wKXt6+sTCophLfKCIBBJm/EAT7Yz5TjfbDpQY
LPimyWT2bCNBWnumuOqMB/x6wtxLdUXtTzcPOIrrQmA1kmN0Q0iruUm28UHex2xh
Pjz0Ip/7/LAB81TOz6/dxdlk2AHdvJuvhwV5mFSj2JjYtGWjn6pBPjtSpSUioFSN
3ADcVJUB7sPuDb+GaeQ81raTcICiNfaxNYUaT2HZaARx++uTFYvKsYlEwRqz1sHE
oJKmN6OYdejdvyLQwboKSFrke/WnGwzNFchKenmO6iVrJBZZJdeA726cxCC5vxML
IF/dw40lWtyF3muGkh6+vihBP4epH7geHNmgoUTctS5N7T1A+C00/Kzwp1JZXNAi
MxxPnXBNadR2ucin4uhru0wPRZWEfIl0rJHvB3ujTfJf5Apd21JjGHbl+mSlV9MC
tHYIZXhUz7Uzp7L7oPYOyVWuSk8fia9rk24XcQeExRIZ8iKQwQNazJ4s5hgLC1Nv
OPo7KVsRBMile0N+lrMxtwpnxvG5xt54MUcKIVUOyIcxHdZz2tpEC7DOJ0PKfofa
39BdKc9bdFcARmcTBMTqNmy5jHmnJmdjJitX7WQL+okRA4Yedh6sY+AAynWZ8U+U
60YajVjEfN61RsgOx5PUy7nPkNKCP/rw+c4lkIDbE5vUj3DLfXmn51n21W/BmSI7
F2tnveHBl0QTs+B10gVUMFh0wGSIGEsC4AGPTNmJG6JOC0Gw+xMddfZSrS57IGpK
fV7ZZWSmXxOmGnJxGfJsPvW1XkrhrFQ07Tg9ViriMc3XC6Ln8tzJWVGy7I6ehWjK
SFU6bqkpzsNwgcZroT03Tz84NJEua9Du6gF69mQsuQ++d0LFi6JwmPrpGIIziVCR
KMx8NmX9uybdwB+u4CgEG4uuwbGiMFvjwUPuZU1NIV6/3bSxoCisBLn7uu5kXPJI
VQeqRxN9Z6GXqfJJW/TypTts9xv7CA/TTSSjhjllbf9cbvi3703aTEbcm2HEU5XB
C0FcSTlrEB0iiY+t/c1XwmI56QaBq9UJRpxf8i5hp1YtjhWUm+04P2RxYsKHx39v
FRTnF/UvLJf2vpgaraeWqgAZCQsTF7Vk1pxhZAGwqjBsLS4ydbv049m+3bkghEPF
JaFTCMiXyegjwTviyGGRPoJVHxlrvcoeIFdEoTEo3q1xKEcQZcQt+nFb/6vH6Bvu
YCyoCkn/83VqeUp7ECCS0KhGLpILDF+XfnpRvX08AeYyJkkDDsmYFHDdUtX/2a/r
PW2+pu3UoUsjSKlRNGW72SkRKb8r5cnBP/9v3S5takAvQuMVfFwrhd5coQ+XXgKd
4NVOnQCkzo/uEJbu7uj5jOCVEdQKIhumzyL4jSjuAVjB1SlW2CuswLK9O+/mBwlz
wbGQ/F1lx00VchnN1RKYcudOlBn1qQLBHP/UCJNRTUHLiHyGOusAYWUk6G69DP8L
fXqB/ei96rptt3D8rbX/wHCjOWX9J1HDj/9YE2IdR8rW+Lpg9KR6M4XAO1dGwLZ7
9MouhImpt/+DB6xicwGhnoHJxWhA0vEcpKC0NKX+xElzwX6ihl84k3bu6GIdjbgh
TzD6McPitEh9rEyhuONaVWrfhaSbfrNMPjNRJy6TZeDZRr7fPG9Y0//54dFxUUOU
XDEJoOJp1JbXAM105XxEw4GkPUb+boi44I3zKmoFtLWB5kYy3nsd2FSqg+QppLaE
ptADYHK/1pxQ4E3vJLxsm+9Itg0pbLIytZp+6JNoCNQzoiiW4Xvas+xYzIMZGeZS
hfAjT3lA8UrzOgKRbIcZossTYRIzkz3LIGbqcDna3kIY1hqxQogTHKU7pIUo8eEL
E1Zt9YyPcb8H4v3Y/AIYhVMeOHnUzRiTwWvNBLczOYWCqjPXR2UI6A56CurLVy4X
js16tk34kTfPrJOEs2Diu4jdjccD3kjN7uQ/ojpLJiSyDiFwuTzt/j466ARwPGug
ZInIo7voOOf+8qY+LPWGH0QAA6kSpda3Muc1dqZVcm8wO7zofK/J2FA9rXRMso6q
Y6HsL/5seyFH3jRYAtNaLwmELWkydYXfs9stfyi4iAKdoa1f1SmyXaaHepPAR/Ah
zuQA6LCU9bKs13YVs5nZlUPhL6B4/RJu4Z5G9JXvFAnKW6u080f/xjezm8hTKK2Z
VzD0u61Uuz2hB5sMOCXLP0wR+gwkSTtPhGoO2VdTYBMK56xfJcyQPO5IyENCbCX2
vwZ3zZPCVNC/SXauf0Xryp0UiPe5gRK2P3a2xr/kxCpk+XzMru3ATvH6f8ALb0nj
2M+7zteiwO+vflruBuQpVZJMyz/6rEJQzKxc7EK747GHnb+jUv+kdE8q5JtVaXpx
JC3fhVKhVYz61iMn7JNj65FqQqucLDlqwkTxWXvLfsWo6iI38OsTuU0CqXqzNILT
yu6QoJqDW+eZwiZLghe7qRidqM7MQ2bpFKQMTOIRDZEYGuqAF192SyN/hvHplZ1p
Dp/V1IaZstLW6u+ADAmAuqbuCr+xF1d/429NxIEHIV4fde43z7WbjtbYU6HiUoWr
ISIzBKJGDIo7tz8EpC6/KH1NvsyzxZrEIeSPcdHhCM+7kkF0WvRm4hZXlnnTc5Nh
n+jg6wTXHFI45f6nQB4+FfwULR5XUxmi8Dg1uTsEHY7vsVoj8BInXvbzXW2WfHyL
638QycgJx4KUSFdpZWwB8sbmGtl2YmByWBR2cz75guobdxOeOBXeSoOHNhwB/6W3
yX3JolBf6B1TFbNJfxGKEkgPVt5fxBGw9n0DN8ohj861UINylysoYDot0RzAwCEp
IRiv6vZHYmmfij7lGFrp+QcPJjt0Q0sh8Y8Z/HCHRiMdajb6Hywco1Gru5J1pGxY
+prsA0aMOmqiteqpVNGFjtUeNYvneExwAi3MhyglATuSxGKDnnUBagAe3Q8SUBhB
5GpbFczcK7fdVGGZZ5iO3umpHfKQb9pR7CfD7udLsHn71dDPuI7LER7FeESOCu+r
vRNT2uxqoAdZ5K+MuB/f3CCyvaSl3l/inmkHkPjuQDxob6G0AnNBJHQOYN3cfFn2
ATQUGsKx7GMYShuYeBwEBTSQSa9ocxpPIr5uGOeNQwP54lIaQj6tWKTwlsSdYqiF
s1rgMiB5cwnGE+x7Aqnhoruc8b+TTsrac/rvFFV7wcdEE9NdyFez92KRY/QEZD6y
TV6tchQNVFjOS4z79OlCd6eYHsRQ/VwLiZPObloq6oPvK7lQic+NHknNJV/TI1yK
+40zHS+i2KfUIGeylx4HB/8ArpyFmL+T6ps+bBmfWPBMljLL8XsCrHDAx1Ybo8gV
FxUVFnVDYqEt7L1j4GP8fLb9htUtIt27iO7lMCDu/HaBu2NqoUcqaThkhfcescla
iyN32OG5fCWdzmwrzdORzgJw5B4kkM4KguG130ISUgT01BgDh5KYPe6Lv7ZnTcGq
esbDFiHvpYLFnkvuaAJwK3FhCQcdai8ONSP5tGgP1sYaEPzTHU0eDoF1Dy16B8Jj
Q5ZTfgnhKJ5VvyeOx+L6JdMD6uaFh2yE3KWvZCHHIvvivNc9hTkToMc79P7v2+QF
S6IgfmSWO4FOowstfnbBie0uaVW5i+XtcLF4plitoICMHY8Yz8JuEfNQtsydTC6h
zRhQCYu/6+WBHMD+JZyE1c2VHsvVqBoO8LNJmZNRyQ9N918u1T0pDCSWGUXDMMSk
+uRer1bvsNo/6ex2KUbvcVFSHPzh2Y7eb4b3nVZgQ2ZkFuf7RHCWq2xmf+vAyu6D
Xpbb+N0BjuIZw3WfuAJo7SEym+bssJd0O3bhz3HIa5zCWdX8wr/pNmm/rvY9xSdP
7zfCyz+Oty+ZGcQ+sLXE97Pqq2xmC/+hzIDYxcDXTTRX2zdgEdH7eBtvKQYP3/n6
LccSC0LYn2ao9bgARfNSpxTrAvl3qYAAGT/fHXZ4tzXGC2JWOJmKowSMwQFaloiI
2w7L5IprrQyCNYswqVSE0mvSLOB+/iSexPDBvo6TllJaDEK6QfhJoXZl1e0baBTS
jAl5TZ7VfeOpySEct+GKpo/0iBcQQmO+DtCSa2BwQ5TNYig2lkYlCcyPv/xVmd97
dhqY9XLudjF88ip/BthT4iWe+ge8QpxnxpViR5Tx+Yt8QOHEwdSjhDAfV4Zz6Vaj
m5ZDPRjWCIWZ/A6+QY/ywX10aNfA9hb6S53pceZpg4N9joBNyQ4lGYzHZ+uxt438
rpZ7DhqHTsbH0gCBzGgP9fLYuARcWSrladguNqFnDTmpRdqZnkdM1+FMvW9yQl0k
ctPjBJxWLJkM9VRldT8ZnjPPyqNePdhEMgKNhasOJwmSNkDU3Gd74u9qW9WLr5oL
aj7Br8ItgKuGmq+LTC+4XIW1IuigAmAtMyTAzbdmRKVuo7j6IXdVW/69se2p8yUF
jfkKClFu3Ai6j7jWsxvL94xQQ5+6Aru0jAcpJSSeeZOfmP5cprIPYB/ZcHY4smWr
yCdFgKlW9AJHAVDh8l/Z4ZUQmsdGsPh10EhI1YJQy6ZUWP4DAiHQ1LW4uHYEr54C
qi0uWWKugAeFYE6JG6oHctbSC+XwL78YDVgdH1RQ599m78h20Vrk/Mkpd3T3yYpg
938hwWzKMf1xYS2ZKpV/1nB/4r4tRlvn2/MhbXRDsu/DKDM7OcRl7T5GfC2G51nX
iZ+ifg9nmJVXjFyKrUDjxGJIJT4UdGUWV1vh3I7yFTMgH6idcSFvePjHyZzAsUre
C8VmEtStS0yQU+WBE8S1cOp6rzh5ZCrh/kYES9lh0ES9/8anS26PUgUb43ishGN/
d/MpUpSlB7PbTY2QP3ZP7AzwZYyejj2vuvC/hDhOrGyXFSbuPRyk5iNN2GMn5Xrz
oeK6LeHrlMdRw5cMO9770QhFH51zCUmd+aoYZeVybanAwaRvN1pjMGaqO/qujtGY
3r/bMliy/QqiOyxRJ5oIIdP5At6D8VLk4cD/YxHOAd7KsPlkI2GIVj2xWXf3tZks
bDVW16cMfTuMuLxfMUEDOzPSQmb3xwEd+0t/LFp1/264yJJ7ofIL1GtC/+AVa+CS
0BVEtkHCjLQboVrBX8qzG2o3nU97J38pvwDjUrDsbwFlm1Lhoc4v4dyW/ge6fV+l
KFo7fLVycRQy2ra07U+qGLfk1d8bRMIfZSHIQ5SJR6gv36C5EKySFGLe35crTei3
6LKrQmbgbSMHtYZWa77r+4rstG2aTxosmxL9i0DGDdREqf4YZsltT5XMbFpNOfgY
bvldbjnNbuDDhCIHJupqr/rzbnT204wZak1QT7nn2cih0NAVTHwjvt9EI2UYGlLb
kaIsSd8MYxfz+GTAIG6sGUhAiSknk9gx63OHKL65bnahtDepuzeXvAhs0tOOSFwX
bLHSyfrkkLsmCXV7s/zld2DqSQnuxMyvU7QYH29c0r+y+V4xhKSYxiSmuxOwSNDS
m75mYogCbWPiEVZdtIVFsfLcc46hg0qKsBZG1bpZkrPCUY3yLqJjMrwNW2wNlL0y
I092UOeTx88IiRN3Mwa7xeFy5mT0xUZFSkFFKnl3DUmtwFsBMJz9iL0Hj/jil5G6
LQ2w1NCt6A0JoCS0L/FC30dvc3EloVvqQTYIIePLV/dTNvCUrisxDj4rhVLRz+XI
wzV525B0GD3cOD+fTHKcttR/dwJWL5nPclMowxPp7wpexLCsuLwDjdOdvmrvz8MA
qHkybWSVyReh2VHaQuXoow6PuOz/cxHpSZUORZAqCuGSwKHAHvb8OCfIry/DNSDt
FshlVBbwlB89vvhvE/ZDnMDgX3+M9IX6GeA5ws6DMEmzy7zQkv6STcysr+x6k+uu
ZtoZZSKU5ENBFkxUp2Q9IzowLqpvRfEX5T9V9cc30I+Le8uirVBMoHbGQztTLmRz
N2XPs1gzyx8vQwTJ1FvU6WmEKV/cHGFH7jcfciOV7Fsxjel/c+bfnlhGzfUapHJi
LWnuBNmPseHX/+QWXC0cfmb4AATLSWg9hVi8uuk8HCEkjjfb13MUb4q5c3TAklJl
ScF+wFMO0vyU1A3p/V07snGAdweOKKfYrS0irBN1+5UfTuc0ns+pECHMsI9lZALW
EXVR/6v7jZaZtWYLKLC2seN8Q6fEnvzLEjkWW5wRHb/PVWdhgEwEu2iAzrQFkLiF
GadJ0mVr44uW97wPxiDKVtheEJeBiTTPGHbc5eUYgw5TaPDjRV3JhWND3EVoGLXx
K+eAwF/C3IrXGp1ViLjncBxzOeqLl9ZzzUU8rbtCy/foYex2AAhr27ROeVxDJweY
3ZjG3jQp/+wEfezu10MJ0Dxd28yv6HXSIeGuK958rGJhc5fuvZ3OTd7NnB3wkhV7
1qbGDQD0HWbgH9eVCoRcESn9lb9Patnpy+Ckn9sVNSkGUPE0BWh8PJtwiauxJUrR
jqzRiiWlA58rPUrCAiKif3I3ZN+ILtYTuIKmTNyLTYY/syEeY5KhfvEy780yd3WF
zwSw3qejz49b7TDbzsLRLsFZPXT6qLYLby2EOwv3sXpRZXi0w83dLxsNF9wJQ7Ok
xcMfdKusnFEVrPEpdzdGlG1OH0X7mzLLZPjHq4a9D57mNjIbEI4r0mNqt8DHoaMz
0w8wJGwZxlKtz1g3vp5VYip8wo/E6jAgKZ96UYjzBdF8uo9Rz2zBMYDTTw269qBO
0lxyMQ/TVZ+qBf4knSM1sXtceCDplLl80FnlclyE2x7d/Z72Gfkduv6VlhCzjxWt
xHGARDHhC/7SURtWi+8ZNwi1x/3KW0/2wfnWWICM2uEwcZg8aN5Qw4FJIMXj6f8d
F++hT7HBh2KMZZgNzh6kcULyNHhd4ss6Lv27ttky7Bk+2PguG7dqFfuTwrZlswuY
FEKyNM9e6k0OUFpfMtYnPtwWPbkkXydI43P0gTiwvSPDUpqqk8l6XKm1X/GBiEvy
npvdbzne5lFW3zyevTLq7vHSRzPn6kB0Ffpq2scgNh7/zshlbmU86N6o66t2B9oG
Vv7uur1jarel4wTHIVP084LAFmptwqt6q6hg6XQeSaVHsygCX761N6RsbI2Z1jM9
ABNDeH0AJkUCVL5iuN7u5ZL3sCsj9PDTxTr07lhM2QbzlYUPmjO//vqkwHFbByo3
WIHBtLy1KXnu9zRDEzhK4rPfnHuTU94HFX6aGkdEIgHxK81dO561OS4YJKFZsho/
s/1FrCl2Xwf9NHdzYUtkk2ZP3b1BsMbSujD5h5tVtTdhJ/KnKlllmKraL6j+DrAN
UnM1QsJzDuav2naIgAqC7Bv9nLJyrV/n02jJweGQ/Fn/f0YsCKbK866boN8PHRBA
eLCeJGBIgTdd/YEgJVW0BvtBEtiDxu5WIYAnsF+Gabf7mLVdSHdz3ODeFEPsi2Jw
5aXP52Pq7HQYrSNQSmYEdZP+2ImgB2Wb2tRFns97QOqWuOmZ04VQA7mNfTSN0Yy1
VLDmV/EYwl8qYvhIjBbJzb+0xllijgPemjLgr6U7ip4iJtGEl86biumDX9eflbvT
zcmDoC90YtPx4XuB+pBkgOlqUbcxI7hQ+sGiSWh+anDOU2+edYcAjMBAR/a4ylR6
azQHH8+a49jYI3u2D2JeHDEZiPfJdKq60ffIPpGmENnzIGkHDHQWhakmIDPXaieM
K3DFa4mBhZqfUd5Q4LIV4hAHVWJZz7ZqptZJ0nNl/ioUWXF+QU+8/GKW7TUNgRDY
yMDgDH0B0KKTw+ehL1/Oy/ffM8mUXezTDCxzuyFbLpNyfEiLy33fsbJEj9u8lB93
PhJaRF7SX1IOjXluF73Ao90bH2xyt4Qvg3R9KUhN0Ek15KM9P5OlWfc9FVf1SAyg
mZ/5gTUGcNi4h5R/J+JAPzrG2Gdgg/gWHtxWqRerYObLkv2XSuR5+hZNDyqbqo8A
Wv8p9BTHxntB0WzT/sEgG15gg5vYoMGuly4LfKVDkeFZ3rPgK/AMO0lXIPYq6gRN
/YSX8ywHZXBHWkMMGBlZz/Dpdmz+k8ZY9YAvpVkpibfkJOV4ysGc0IAzLAysajwq
aUq8CezjApkH4+YhiP6j92rFTMlh+kInDjZ0y6WaauWRPfrWfiruD/1iCnKLTbRN
tBDiXWFUCUsRNiOZKHvHx8IRrwOKMtGQSExhOjDVr1B1fvdk4EWWluCsrSts73CU
W+JQrJaiY3pRIMmtO2U7coq//qR/zdQY1EHguJu+6Q+ZZ10jbj3LkHqnKwfOTJCs
a14AJQMvjlxIbxmA0f+kA18Jixn06yb8FfPVe8Pkb3Y16wpwVJX0AdxiCjOkwJOz
zuKJP2ZSrsorSSWKa/Gu/+MHcga1PDAiiivJtiCBIuzhE6ClcE0CEnw/vuGYrZ8u
8+L5LLwxX1uJBEmZ1+5a4UWjELQZ5c+2ECqZ4naxjNepZgCzsEC7jh39BxAT2COv
xon3T4z8KGlSWivMXHNUHrlN17c0GNp3/qqwP8ar6iKZepkyU5zSCjEYm9hXbz1R
yqx+QmrBZuTJiq16OEhXUZvwIv5Iqy24IWGzYLjafkeXOHB99j4qsmu1erlzgrZn
KAXCLuDPJubDmODpkxhQRqJ4mAtrzq0nTQZzBACytzUhadjpPVGBq461hxFkfn5c
mcM355hml89zNJ3S+LiqGwK+wlqhSq7vEbE+3o8MQNigxX9vHZBmLQZpptgtyBc/
nAi6n1OB4hOaoXtDlrq3LE1mNtoXiZIRs3ao8YGLF5MitZFU13i4ZdoGbYz5gUGY
A4jxf5DnQkrJ5Z06HBLHWThzTsOFV/2TeYQN2blhnbxXLK+TWovY5unq3vnLZgm8
pU7d4Q+HOq36MV/BdJSHEoQmNWTDZhUZxvKF5K77/6IYzLE3aRIlEP5I0I+8HPyx
V/VThyeymxOC6uEenFw65pwFymDLI+X19p2aaf/GTkXpusXcE5LrSKRDn3IIzs1F
kAH7+NwmJjVnhfmCphHsAAp8qafzrseYay9ayJXKk7rt9zTpuHZuRdbd1i8izrhU
PKjLKM/2rhNYzvPAmMTALT3u/NO0oOKV91s3ctBtd/4DGVwhD6oR+SaDSiTaqOov
ow57MpM+ekLOeiSsysr9TJiyTw3xMLbWT9SR5HUj7rFpSqjCTYdJkSkq7AXAoH/3
I6qTWfiaYa2zI8aT38YLpFcYo1oFBLxNIM14S3LSVhXUneElui+nvSOayUZ55KTR
PFEvwtcgYqnRlt3C0petewzSZe1qe5+q8bkhdgIRi9gxXc0lj3I2hEP38D26Extb
djsGthT9RGtJvYyMw5AXPViwE6V63trv9BvE+aGTprJZl0CasObvcFc9CZXVlJRV
Px9gHbQcR29FlKQf28lztGNSziAMAw/0MugpZQLcdYsMewzX3/caIXj5Fz/26SA1
tKUWDm/6ImpVpfeWGHqzcJoxRrIsWNviqsdTRVkOPpnY9LhSRkHL73xlYqN2MHx9
7/NPH+nhva2W/5orYyPIe2Xwd4izBY8jfDVeii/OWpSjd832gSY2fq1Z4sy9UC/6
dRJLYIBVO+cDkF1BpzNHxVHSE2peHYGphGi3xzKrc6W0Xvom/bDq1KN7+yJ0plhQ
uCChqa6GdMcKyMz573hW9RrEjon7ULJqvIHaGHKHUktTYwnZAVkLaEIPiKmTFzeo
X5AUG4x6eWDsuHrpfa6rdEOPxWB7LilWZzKZDJ+6rD+djDzahBVQCyPVB9U3FSLI
Qq50zJuj9C9HN+N3xyL2Wl/uKXS/8qT7jCss+Gu86BcG7T20PGnEnuPchmFkJIdk
ctBiRqKLhgxfH/VialJebFyP4gJbHUUIdXPvo1bI96WcUaz9x/soTJMkQLCCDEi7
7uZaiV1Y8bApGw2CaYKQdIfJn5CdM7htirzukgzB3J4SdOw3kS5yUB727GSUXGkq
LPZXd/ycnilzJdPXxNfbnULxrbePp9TfgRp4/P7AyKqx3Ec7tWTE9Q9qFRTC3C9J
c8SGnAgZ8tHKV5Nr4uQxw+AA+qVvajHLV3ftWEuS3sNwuTagE9OxiOcIz8gW5PAK
CtL6HFC0cJ/DBt1Vefb39OMv7wTLXSpGcYipgNZxK8gk1RaMROFOTTMGMOMrA+37
CzvDpPrTxA7aYjOU0MR+HIiJPMxc5LfASbxi9SKYOTtiGND2s/OJa5AyCgVd+++0
QJygFFAKGv7doaUT77PlfV8kBz8/hMSrao682ceUQ90/SPxvsUKntq4X9FJ8l0Vz
pelM5cr31iUvI6SZ+ktXYHHa01GFLa0E7j9tSSVG6FrM5ujsMD7obGZ8FPYJnQXS
P0twnK6otyRkuSPqIFwEBlznwu230BupkfT1o8akqvL9D9CaU4LKsqPUuNc2pr02
6LgphWW3Yvp430LMkkYE7DUc8UNv1H3jPIYbJOGNc6qjw1FM2Dxg43oO+HN37lAG
iRgfTDtKfpNySJ3vwTjeT1BiFAJNXQaWyu0npBm+vaQekTlseqwi3bY+b27z/Cgr
TzpMGdUGQbMgXn+8swb0HNCDYfkuakJ4P7usV+4g9ubqWJd+g1NWT4gq/BsjDPFQ
DPE4lFy9GmZil0SvtLdLk+HYDM7kezFyvpVKHIEQrYabhyJljl4lbnsqFZ6hRXyi
klQsaoI7DSWefjE689OPHcthvrd3PoW2eRzTJUyvY6w/m9kB/s30FGJX0GrglbZ/
MaVXJwWJ5JOsrI0BLJy3Vd/JZq4UqA/gHs3mPVUxygQVytbRElHf8z4ULEZUb3lA
9uvdiEV/AUtnydZfEmJG5WG+UyWmPCWQ3hk2ML13HYZelfRlI68JWUQK69q5Soky
EwCtVjJI/vX9Dr+mKwe2n66cZV/j3gyM59cCqzIj3z7bksjaWY6DFHnYRAOfsFvS
7D2HfuiF/FqswQFcAp4YuI0w7fn9bgCfs4sGRUd7kZa/PmQIECo0zrOLfpvV7V6e
Tt1iCg1MnXk8epunE3J4IvFwjp3sUuSi6c8QBOYCzZER2OStgaJsYIPmgpsgoTZ5
SZAZsxx2gHvuTSGKbXxZVLUoPWhHqlcSRX3bu43/ZH7w8zdxbcSgpM1pqbnuB9gx
e9H1kR9cUpBswn/FPIRNVK4OUFTlt5mXzpk+wBoMQK/Z+fxzRoSP+5JUUdcHGffc
OsfOB0/uQ8W+Ro8gGi8gDbLN6RwgvTx2HTy/KX3f3fBsLXKBIXx4GLvXUGqmVoHa
9V1+tQU1m5ZcIF8UggEpHp8MQPmhx5bKdzFuHZn8Z+BilDW9wUfBKRnEg0uWXrZI
J/tvq+qagrou+ZhvFY6EsDJK5QnKRlSpk8THDwdKHyz6kJ3cPHJHpl7/PE/GIQHn
Q6j2a/Hq3Dj3z1xXHQSzboy0iJem/EdBpHYfFhkZv1Em/3+ch2AY21lM7NY9i3oH
lt7o5JO8jvhrGxacJe/ByLJBzyHTmhR5b3FuN1Yxm/sXC/uEugeVwSNzZtUN9Ez/
d/Jl8Q/4d3Im+KLUT3IDakkMGlE6xt0aqTNOE69Mhm564jPSFKuAxsKiAWrBsrm5
mGQUhnrgTVyOqVlTbLakwzqFXXCA9vLRtdrFL4lKPrvQEmq5hL9EmlDGed1KHMu7
BGUUhSPjLVfoEE1vsq9TD9BEz+dLVkQdkQ8A9o+nso7yw2nYMtC/y0Vt0CwbU7AS
IdVfpLyWc4tWeCHuLqDN4v1nXPoqHGnre2ZozdfwbBKAQpTyhGOcIC8ENkB1TnUy
0W0FvaVgBJm5O3N30TaETwPY4lgsNnDBVu3vuK1E6Sfy2dtok/0v4GIOy71bo7Xu
aXsGZj6K90DLQ2rqDJRNcD7/NwlcM7gAwUc17cXmDdy1utVOJBaqSl2Ou7gm/axl
q8l4Zd4a7LsJG2KKBTHuC5enIhrqL2Li42x3PcvMGB2oZKh083a87ua8mpKNYxJY
7mSlTtskwwrfKzle3j/dHCNaTXDlA/oVXjamoys7bgc7ajI2xOUsSf7wN7VnQlt7
wYZ4leFgC+zmFTzDPPPGkYa5vLsdY48RB9MIY9dLN4Gniq/cUJ7t9htXfoIlSnW9
YmBwMZpriaGlVuL+iKeyl9xQg9XLe03mKvI6NdQswSTb6dxBeCvgZN99C/dvc5GG
3gTCz9mk4XA4JMF4dXdNRE8rE4efkaYUPyxk+28DDEeN7fb0G6QCw4yp5ChD1rG4
m4bLSik7NHs0pqADEZCbfrJFSye5PgpLExeCkiekt7/U4byUcwwN/V2Lj5plQeA0
twpXPEwJJ8oUlOcn2Sm9CfYwqCEtyE5ShA4qaFf+EBk0YqznpSC37VqZedb1S3ee
iyKkTzeBWq7fnqfNt4H6C8nzD4Hb/u0+J7nyVMDCprLLuNMKB863exIsFy6r8NKZ
6p4fraX45RtNS0IY96khYybH6CRQIHtQvdbRZ2jaAlshKS+QOe2rQXPLukBizfF8
6X0lH/j9wfaMF2tC9h+dSt1o1SuVEWviefGCRLaV0rlbnnxfx+9oB4wQShMRoxaS
lK51r3UDbZ18tcXIUl9jya24wAoM9pbvWjs9IcZcx+a0ktf0Sr+D8qs9aFU2BV0q
Lj7I7VJNN4DRNIOke9iLeLKaS2NCpeGU7PANgWayMb1RTyDWVA75sMaREMVD7GQE
S5g8Ip18Doti6nEYvcwuUGGMz1zezNZwSYZ3vTK0LPBtR9mLNLJ7nFa/uppUTvA/
ItdIhlv7jWQofaMzJh+PRVe/14t55Lnf8Or6fKD+pyDCnJJl5qXNH7w0MNcEinRX
nOfVGlO9GApfgOoL3TGqr+mxz2+eWkk60YA0C+bJdyAhKiWOwSvuzIg9U+ZqeCUD
TYNql6goSqIUDJKosCmNjQTXEO7v577uu3sUG2L7xO+9Ockmj7B6GkPyv4CsHrk0
TqtPyccU9O5Mq5ykPpsKuS3ZFtRT41tOgm7LBbmFUqBkVsLMzGP0vddXU8g0cM+E
klDFJTmmW12cQAQP5mZPiQlbdNpZEkFSgeE5S50Vlw0UlxTrrZ4iECEx2f95oXKk
kdYer0G8qtpLo5MSK9G2BNZazR6xLKpHM+Y674AWnIdDGUK5mBVx8Qq9DhNmGsSR
ZbIR3c1nBPcXgxGoeJZUAKNfTu2+tlSbTeLNvR2t11tDRKPEeQqQd2bvOdLv93KZ
G0CeYIvBrTjPuUYVZg0Jlcca8R6FXdt3jZyM6llcEEyOgPilSu/W3F3zM5IjDGNR
JUBSUul/tAhvUva9tOJpMhUC3XXt2mz34AJTOQrDiR/l6Oy8f4SqTfGPX7xGpGlm
ImV5CJ5Ra+i5KxK3WGy6/dLC1PVt6lccC0LXXdYIMUHDULtVGdWNHMmx0VT5P3Il
BSGhgs2D4teel6zIybKOHUcdB0qPGUbNS3dgvJNtfLL2jKZoEFzLqn2NojV33QNZ
dJwSBGM1e9SJ4Pj4LwPXQlT9D2xEXzmX4SoW4XfQawyExn0nmgM7+R2hxHB6g0Lo
YG4qX9NLsSWZpUyUReN8Rc1ivIC1eh8SZmKZkDynLVKAuyY2k8XnGUwi4ZV3tyPZ
1gIvRXX/cCXjZxmMbMuu/LXMe6kA69p1Px8sdKipUVFZ9YJSq+ucLqzKyd4yzWNW
/5bw4wLzUup2F2nVg5FBOFhSV7oM3oE+visURT36mKMZvehpxOkQkSFu83s3yK9l
+53RPENRjjgk9JFz816VVsmdJzOYMccXSG4Gznt44KIaBBmyUfXxMjsYkJMRJw4W
k4YmqTjxaYurgoKvjGSJf7lFzBkAetBH55piExgaTv6/IgQ+MBh6IuCAOQc2IIFb
15KSMD1uR+pXW5SjZzboJElO1znhRvUuqTIWSMFnEBIHWkqVeCaUCMtQ54eQDLU8
kkewgm0LfG1atXURgqId9Ewf6098Cbiw/9VOn82oMW4rB7bSigZPVmnoUV4xVqxG
TvVybab1B27TilUUhc5BEWWv9lA71T98RR8Jihp3agIDArqV/3uQQ8WG6jc8VCYx
H7dp96jESDtAX7RcHS+sakfEfJ/V8DKCS9Y2JIG8SwNVlRKEBZhyTJkJ4pCdL/TT
F7vkdDKsBFi042rod2bKX8yyBHO7wYzYWG3d3fs7D7x/tIkmuRKLohEDTz9BoBQo
azTjy2J8MWlhYKSS+car+uq91SdKs5+7VdILDbussEmmpC4T3DcsOxlfwOmd9nMA
snKXpmtdvH+O3wnXgApJZrC34d1+Udm2olcyVR6mIoOWZ+0CPPaD8xyj7gobcjho
5c0H7G/a/hu9vtzakwHjaPYoncgICgH/nZycWIx0qDSyRMuvidEtEu277JwLjzEw
RcgfXGOW0z4I78xll+UWfntBF9QntmAt/ipIGXqeLXoDM5EGpcRpUm5NJxq+AoK6
0jKw35TvTKNThAcK6zne8FFUpYMqxEMbFzfTg20uZNtW1iJnSGJ17K7dSAaItiB+
HyovMMTj8RgFXhqqox2+qd0YejXMs1zagdaoN4EmALDyKE/NugMJ9YwgVV3m+DOb
aJcDhts7eet0Ln7PVwU7M5SyHAlkdO/68sZnAvi9Kw5tpEPOn/I/T97IBeECi3cF
OFXQaNDtc+78fWLD8ySiS1l3GvESHUcPFy/FdNJCk2oLVZViVVe+kBNCQd9Vwjqp
i9KtQ419Osyt4YX/NdYh+9OuOtJqfN4PCUUsnZFGtYPaTmUcXLYCMb3u29DAJboc
dh9UQNPaY3fxHbQaONopCuxcdSjnb1sfx9RO9IJfunLEjttaxswYEd/c6hd/l33/
4H+CHvCrma4eSq4SvUxSHOiEFws4ymdP7Z2HN7gqesllsBaDSMQbUrMY5BUFQ1ko
FYhBn30qHofz0TCdne6+0qwYjojSwkgPN5choT/qHfHmjOK8M+HAox4W7wHkAcKN
GVQgrMYFreQeYPvD37FkVl7wc3HzGxOpuWNMGq6BFfdnFJVIVRSSNW3jZm0aOpg0
h/Dg4tNAAzOKsmu8wi61aZYrqdaavXs5Kz4Mkg7dibKApjT38UzSC5HTj1hgoIM0
46lzgOjFgvzibyYOgDca6qibcKcUwSMD/PHUhlZqsxg+vqCAqy1+N/V4CiLdxOly
qlBlClPz2p78ehUVQUvFPWC/JAQSDOMfADz2k0unAbZygdaM8TQ7R1r/bkW/+vFZ
uZ+wUkWL04wpQ7x+FPRORLvs+sUanb0toFFpyLkvWMACxZcUyqvzyG2kzfphah7r
v9G7zPhoI2Iy9x+XNxdV35klFOGa6YRpCt1oZLulnNTOw+7vvXWLXRPWmbQ2/f1d
WUm4X6XIn9/l2tskbU0Z+qkJWt906edc2hBXzliQVez17JskfuQb95NjJY5/wDtN
8R06ajNomLR21DHVQY4uc8f9Eha9yAjPzW05HvwGj5wFs03Hz/yhh5F7jO+9xdMQ
aQeykSQFPGLWsZKAsRb0y6GVGs3b84sxx9Za4336huRHelHQmdUA2OoNtFRrJXL4
C1LH11Cz68Js2wCztbboqQmf3CXToROTEf7jXjzBej+DnbWwmh7kowYBys/SvWPi
/1owpEu4k0XOfVpe305lqRO/BP9yzYLKk6oDp4rOHGrtumsvhH+SST+0I+7MlJwy
9cmSJkTpKAlSDjPV9yciDFzDawSB9kdjTZVZMi1b+q05HjEN+DY9C5QyLYqNy5fh
ioDPRq4lsbN/qT3Q9GPzb1wnDl1KaXEqYXHGZAfMjLYqQlcrlTVuvR8mu/iKcuWy
qq/7zrmejWwkqTwpFb0MQrj95bD23iqpWo3jYjt6M6Odt62BL9gdi4PlCICf9hES
9EnAg2qSuBD9QRWO+6KMmYpUtikonpybpzBnaA/WFzxSRGeCgS75c3DoqYK4uZDW
o+QU8L8PbpRPiKhHJid+3RLGCgIq2YNTEF+j49aZmgAPCiLMdGpw519G/eqNXkmI
isaDks329ZedJ+u8QoJV+24ACZzFp5lfACXKKENWSwHR3afU4EJcakQ4xQ23/zHN
jRpD2uXZpQDxOuejTY8E2NtQeM0+fq9EnsVHZMfEpF/1CvTTlYbNLCW4KHi202P1
faTyLnLBbKKk7Zj8eYxZ1wNn6CPHWHCXE23rx2vWMAndXDETS0V4JgqWTNsHyD7D
cMI+JxD49pAqBUYlS43Bh8jpavKA2IlTVzFyTI1FZIDSnFi20uO74iDf042t7biz
vxRTLDGpDGjonHT1Glrr3vRpnBc4yCaNaE60Y8Ewl1ZGN+ywFPeTxspS7vNpcsIQ
BWnrAabwcZ5TuFWuQ0LMaFEZjnDmWaJWYVeGr3gEsjp74bPhBqHJfUn630ErIE1I
OWvgbfXliD29eiE5NGdkgzo/FlAJLJ8cT7b6CmWAGxtaYxBn3d0ETXQa+WEzNAOF
n8m5E93k2NMfB9nQJ/Mgt8Ie0P0fQyPmF5fjZywN5t2ahNNJNk/vIBK3qICGCChd
hmpQTbrzxu7/blgwWR4BIc1NBZckXw3iOdHpE6qe8gmVBljX0VVVOrgw0tcQxeH/
DhBgPXpw8ltMAmdWAt8JElzHAjAQjX/rwdxNqzhtJTD0khz1fN59g8i7Qxz5tdkv
cI9wn/1lPJpFAgfNLecZLjeh4sJPcZOVrsNwcgCSzIzcK539Ux/5ekkMoSw4hT+r
jOqTX59CoYm8St01HEwwnwhZC0MM7CAveA07Wy+EmE/yQ9i9EB99sWACMuKlxgX2
eJfiWI098rjlAv4IQGx8NS03430BhQxkKLZ8su5ZB1BmLDhAJ3odFAtGvTGKtS2N
AOQ9WO+LGsvdz5v/mFV2O2hGgE2d5IRLiG8Won2sTwq3DrQdWJhFcXEbtYsr6XJ4
h0bdTmyZ1hLTykY8bBiHQsKvSWxxlrb/Jaq7XW1+Vr70XuYJaWjueSh46PGKWIq/
yyOoQAB5ECNfTN6l1yk+/czh86m2f2z6jRDaHzcQbHliQ+/5tfCAocmT2oyzZth1
6NCa+VK/qhFKWJOeQJtMVvzLuIzhkzKFBm2+mhSOlA+Ej7N6GeQYbq0RYo1hx7ks
0KSvYrqkZY/Y/CHzIFNW1GQWfhCPcpiIXMxWabuwrkivQ3+0vMdYC+0CI75KfxlV
IbmPB48pWk7fptzUIme+y5vs5cBmrn6LoA/VgTQo27mapTV8Ua6mGUBPFN7zanBE
EMT3Ln3lgWxLILx68lS3ySsTJ1O5BMOnxc5Xzb5bn8SjRa0nOvEYkpdZAahFdGIR
kYupxcfI0rU7VgjWJwb6BEULp4DSml0f9g8kYE/+QjVqtxqyOAwJfAWdFGw1oPCP
AHiKpaVYUScVdyRZEZ1n2xewBED5z5pZQeadZtUcVtoe3kPSlrCgH064W/qX0iaW
MBgFFlVwCbEMNKlUKsk7PIoC9iHXKpdTHrTTBN5wsO5sL4l4Glh862LCxXEpAUhT
Z3yljqntd2k72poJMQx/Q9kZ1enNQdbJiXYRE4nIdU+fbnEU0/g9Lb4Qsqi7IvuQ
jCoVtHozRgLss7KmDlH8X2olklk46vF/pT7HzhhvIu/5zBGvN9sIOoXeSUwnouBr
J9LmdF0XU6KgKIyzuBk3QicjlzMU0E2aE4VrNRCJV5AEHXSHMHqbPUFqkpaqox00
XmtGd8Iw3TgbXOeJiH5PcSvB8V8fBPHXDRHM7uKTmIUCM0xnklEcrnIbHzCg0Dsh
KfVFyBjqvBmipXoEcCPOF88HgLgSxuJ2eNXP82XlTXYATOTyTKxL9wRMD1z0LBQP
d07tLMFdJLXwKrwxoqnfPwgqFw5QFjSAzTnQaAd9+0eHvK3XXF7kGGea371vOzEO
nQzC314cuyFbZqttpfXjfkj0baWRlP8RS720djxO6ERCAKC/OaTYtsK1rRY4fprb
SjC4MJbj9WY5ptPgxeb3ugRJwSQsUIMRfgojalokFuAPGVc+eL+b80ek3tgc76v2
JgYRi7+TpBlnfxN5qvN3jqdPtZnN/r14y9/EMdH9rEyuWi5a1VtgAV20GhnHRRar
EGYn5c4Br3yAwE4XnbVTVeI5dUxn4+8nP7x8CqF7l9AYv/9oj4jwRtzgPz5GrlMu
XZzonuaDBRDy/Y0MNlzUvM00gOW7D+Zr38Yscp8/Wv4C9zjjaHYz66458F7g9D3X
geaH32YI5USNAb4nRJtzwWUhcAuA3/XjnxjsnrX3Vdq2TnPAmJwqJtMV0ZvUnK7R
5RECezaSZeKD6tuXAHiVEEnXyUnavDofjAWmTZx25t22d2mYd0yuciu0u27ZGO+g
VI6SM2HBkn8TqcnbUi4p60ll95f1q0geRK2I5hCSQeLqHqUHhwBGnueE3jZuSP0D
oXrnEQ23nBplOZlxwQy/O7hjHLFoG9yPCgFG675WTa0x3/YvdyJ8fXd1rmjj/nBf
dAia7mfXBzi1izzRYCZSWCe+kyw5Kk0FrFgvNX46TLgeBwn6Hzefku7a9D2/Xm9k
hATMXCt3A2/5L0FSKbCfEIexYwvtRMsNPVWNBHlAtW8fPigWfsm03UQnr9T/Oyum
/e601eGgO+8mtIGPsj663IZXy9ERy5PaRky1zIu+436Bx1wkkr3Mnp6uuRCjaumQ
U9kdzU1jkLOu0PyNMkRgh+PwGe6h9x0+7N68c5FGQQaLF49efDWOlnWQUkz4gsJL
sBY/K7voytZYrk1yCUXhSJrkHwxpu02bDsCvNSRkcH0LB59GGSgKykE2MiudB8rN
m5ZEAGY2EtpjBVN8Ek8qUx78XmpKYzWp5uRCuKxe7+UNev+u21UNP41fl4BTe7bv
xHnvaX4ms0tuXzpg9EbDouKVzt1+yj7UjhZK9hXWVUhnPHwQwZJDRDpE5vWHhAhu
7PTKchzbXXAlWf4cl3pqvHAvrndPypi1f46Jqd1FonnKVJBt/+sJ+8UvI/CNzGHN
XKtNeepieAm3ekFE7ouY30I1xQFm/W17Ny3/10nCJ98sSxSNiBx7qtSCaW2hhj6+
Vq/h+24eNIQmi9d3GSvg6ibtFOA9hDMxAqJrz4G/gIEijyAUSrZWDwdUYIKNQit0
FpYdozuQS6cKqk4xlA70rRpRsPGJB4WRm1wkKOK5kSI0s/YSTeJRbQ4w8FdNAvo/
mwxexB206h/nMeRzjpFSw+KByf9zguQ2olZwox8QUUIUU99hH9azvWADyAV279pD
M7qCvOM6aRZJCCv3q3aAhloi6VkOA/7XCdT4AGO9O6bPYa94W+9XuIA9o+3bNdYX
dz8xCWbPEKKflC9Jmx3DdlxjaVgzLQ4y+v9edZl1buEWJV/9ocDqin+a6T2nDsIz
dhvzMf8V849SPp4WfhMd3ijhUVswPXLEQ4JPaqArbKzTkzD6bdG8J9Kv803/pVdg
hYlhI7Mk4muZfTDlH/xC2O8FrmM+Pjlq8TPn3SgvXceOOYs0Ykb4lKiPZDOD4DSc
3aGEvkR7E83Krb51MzmYgXFnd6BPMCdhsI4pakRB1i5Tn6xp+pN/iJ+qxEM48Fl/
jHJLnyg3DbcZb900xSEpi1/MTO4kH6L89hGpbRZEk4UnOpQj866/YmGKr9jr+gX+
2yp/k0hLfcSiI08Q1K5Ye2XbW0ltEKf+iafCqXNrJdCIoG7FBS2fi9cf/HXB2WW1
PErUpzYt+XIPZcvAV8MfsBxCUp3Z0cDMrsVNoLZKbUPdrQfpIekIIalVSiifJPbn
1f0sI+1Ur10qymwgDCZsjpsoi5K6GZB5yeRGLz0lpmnsqdPN0q9BSQafRnYzSZk2
UZ3Cug+E8nztG/NYNEss0mtLv8bX4CwP5BRO2IU66ectzvttDakdBhg7VQKzoaB6
FpjYsRQ6VujhpuFcRSEiWtJ4TQx8BcxRWhbISva3eX+Jg7TpXtkENsfQM2e97qBs
VP3BTXosdunO6pLfQ8MQdQ0HRh9FiuSGwY6sgP6DjFJELZJ88We5VL4Z2fR21IZg
raTw7YE1HgJBRpajTbDVRBYwQkXGdD/Ymu9cOqQzmAmLr8rKjISl7foi66SLWhBl
0xNSEKWg91AoD6FK7DWjanF/C1NANsd1kovqrx4eJjcLeJ6Tf9Sen7hHpbfbR3M2
7ttuOlvkUvxs1+lGpeD3rHC2eFPjcdg7mKDx35Cn4UFDbCTMhS/O7wu+yV0kecO4
pzh+5zu+92BCP2qEkRTxSoz9zWFj/PqLq/JxGwwsPJKXdk6+aBKFrNJAiet9bpIK
KeR5tSKb7YCSfGtkS7fwsNtEdcft1FSEf8s+vSNs3u5FcYd2eT/TTghnjGhM8lWh
zpazzK3Asql4wWGNZvHhsBGPccyrzd5MGUAYo8zq0URhDpdzC6PAJFrEPWhnJuCC
LF+vk4YUGRuoxlhyK6eO9Z1iJvyB+kqSwUyVXFv9yngt5MlxBiZ0+97R2Mhfr8sC
t/m/6LJG+VOMsifj+szW3HDRcQ/yGXj+vlMcVV6wotU2ye7IiJjklJ06Di9aJJF5
51wfAhEpfnTyTg6hDG+e3rjqEEJj+SSXzTksKonbuKRH2jU16o8zA5/w+0Pce/zx
v4XFoIiogiBeTcozgCgllvhF6anRDLnL9/yd6TpURpWk02A+dlmYvRQJO+MTSyy/
olzND010srmf6f7AjA0i0dck5om3krLbAtJA7UTUumXbXRKwq9V3NrcAtMrISXpH
YH8L0pGidTNFCCluhj0+i/9TZM0cA4RXDYQ2aXlCHi0uWRmvXlaRuNDzL2gwKHrP
aIvNuLtwM8YKf2G3jkdLmGzSOx4teg3xi1CRGZqsDjxr8l47pkoI4XzBLvr1bqsx
1Z1ReciXJ3A6WZRGw7ceanhZVpKgkuJgbI6tzoeU9rzm7vyhtyL4DRfnXEw2Po4s
wAhX0HVRYqBcnSkbihILMPf1ClZzlbug53BmC2oS3QypcTRiEaLeGkMVgPkrme7r
mCxvoOpq2tfMdbwjpdmBvfMBnIdKIYZAujQVfurr3BQZWmudCown4vpXH3W76uVr
WQJPW7lfnMX86z4/LagVfZ1HA5Cg/XXDlhwCdW/g88CEhzDxwh2bnAoY6A0YF5JN
0mE6Wnzb7oVUOsZgkgNzcjAdyzqS4HdLIHq1VMk7zksWqJczU/yKBpvceDfFIRoG
6ZuHPWsr4puvbCfZhFxbC467QJckZFpBtcxvjWAAqoAuGvQihyzk/oiyd1W1zIVw
i8+S2y4DhbQTye0CW892xZbNlOBUrRl+RPKH1NYIfRt5QthSEUj4qZGkDjqWgXJN
fdlUJLMikNUuI3PWl3o6D84AuEhP+qWv9Eow95xP3HJ4EOveRVEa8IsukqxjtHDn
LIG7WCfWvE3+Hc01ic8kix+Wrrnd9gOffLDgKmInElAVuALb9RpN9jMaKECZHYEJ
Q7eeOyOlpeDaTNadmLYCfH3eXfri7Djhp9vuZ1N7URafAmRFb6qCs+jJ0jbz/qx0
+j9hY1sxYs+F3AY7tx0Os7O/xayLBrILlp3m5FmYK0Zo1t2Q87KAMlDW+k7u30lB
8vP5QTp1Ih/kUNpngMWOLjqBInLuIkkkpZpU05kZFoY1BzgLExkyn+mkXTTVGf/Q
kv+4vTUu+HKSArj9yHqq4cRR/T5C1nVMPv0sPGSvAzPCcbYEgA9oJEOimelBpmaG
jXxnSqZGcrCu2wzJK1fA6Ea3Uy0bBxHO/7x8zEFB7CaGFjdCFed+C0Uq/KW83HS/
eHlsbLasm43DqjJjvbEzmt1+hTpT8XQubR24syIaAY+NDJj1rik1RYkkhnyqf2zV
0FuDbxVHXtvIrp0WGi6bm0IHSo2nx7xCahrBLG9soalpFDq9rm3G/6QnqectHLsO
/wlL0YZKa51qexRztxGXHK0hgh1oS3fM28zCdUqwWGwOUfUXzBY1lVCA54GIRubz
uVbtmU7RL/6Iouza2wUbT/k6EWoix89NqtLXvudBDfN88tG/8n0X/JUtC8f1T40P
fkqmshcT5jIZQQ0Ugdashz8zDnxecW6+Jr/tQh3oK5WU6kRF+3+KZf69fr0DJVzI
NWkKdWZs+kXCkZiDSlSIXlEzvOV9g+EWGoXTV4DeIdUDV8XNquUMu1LAbDLvv9kM
Mh3EsIiCCHoFtEbug97q0mwxhr4MpXezTH6C6O83tdqcaFxyjRfygWqOJKheUsfw
A6kebO5T74vSPOxKZESMC1hwLsetJLe3ZoQ7Z2i7Ag6HnkzShY1wbduVVxtHtVDP
Ka5xjAeOfT4SS/EhC2/1MWHYHApOsPJfAy4IcLdPtq+XY6FOBfgAu22dQKK6wmid
Oox7wqgmmP0vri+lEUYLdTMNLCB7fFMLC4r2v6CGo75ZwGmoebsT+WgyLqaYHt0D
kW9bTt/d0B5w1wnMdsZKh/K7AzIMBeVpkTL/8Hf0vr5ytacdiJ2S3mkzRbAgjMfa
tKauk5aMQ02z8d5DfSP+vkEFCFztgQfgLBkG4cyRepVWwg0uU0JI1B7SMH2ISh5u
WsIpCNHffyVdk52zYRVPOjUE5L/n/bvLaaVpf8KAQWR8P0SFkxch/OX4g3oUNPMq
3ciH11b9726nx8bEauzUrWvw/OWou0GnoG0PXz9xWn2T+XRlZRCZzL/LxHkzXLmM
dOGc/Som7SyzcT7F+BpslYj1SmRC38u9SflfmlPmGK0Ox7Z6wbgaN4q9j38Yg57P
/SigWi2wp0KpiQMr0SiknkHWCVdwn8Gr89vbrVfAjBXt/LZdgeqQFbrOO/jLjHc4
3NCrVhqZihnvJnTyBjCubDW0xqShKRZcRw0XpPwGgLVD/XrxGgBfWhZEZt1S4rJV
H4hRxRebadU3WvLmgFwMSkt186ARBfJQJNbrIMORiQ6SNgWLbrKCvsp6WputOdMj
32tMHbwQC0JVYHSoSAW7Yqo1+rwqy+ltKTL+WzPrRNjorQF8qjc9CE9e8S0rdxyV
qx5hQ7fgByR23pVa6x1vEnWF7NKR4ohLSmS2pNMFTl3KyCTwQuWQ/hwCZeMD4uN2
Gs6hbY3/ixRBTpPiXNgi7UrBY3hh9ixJqhXY/z9/dAU+cquUY5epPGlpQMJdfTOh
FXG1JgJ0eR6N4DyHynhs5+q5imYZENdAor/q4UjeCNAuDxYvzzXO53iP62afJeWz
Lv/1hovV10j4/AH3A2Von6wS1AIpoce1/kyYTMEm/hxLhOO/9tpEpkITAzsNkqM5
FqTHd2r2q4qVuYGf8CUAaw6dG/luXoPvYSes39OczKtD2nQfTUL3o8axaelvm8w8
/7KXtOdj/+kOd5bjHeqkIlAGLPTDABtu5g0umNZrDkHkOLGsqP3NC26ScKiErie4
j5SVl9/GzKUv2nsOmYrGtCqXRtNrdFMse4pMJIIyHuqpvDiDR7Ly+aKdlqchhUQB
yAtFYsgD8RCFiuGYMt6LSFIi9AQEDFFuqsaowul7i1K3t7yEb227n5BdHrqTU1T9
fi9GfwmKUEyqOHvDqPCSch7P/DPu0evYt4TQJsXMe3WW/plRLndMyhgFd9ecKtL0
4Cve7l0bY86hkhCdwNNgEfvWTEow6Dz1Nqu5VHrR8fs2fKOSWdEl+WSqNpLyD3ok
SGs6FwCDhVeQjjQKBWMKeputHNnk342hpiWHqYBf1Gd+qek3Cp/EMVGDmvlj/447
ps3uMrT1O4T97U/whuxYpYZ3B+MJCQ+p/Pu1v5jRCClGcHC3vYen6eJEFAEwRzq6
U4Ko1HhO3/vQM97AoKdMXkiuJqflp8byl30cbdxI16YlqFlNJQbYC3YbQkxBr5M7
a7e4AKDFvFBunSNWXtBn2W4T1go+RoY6cqwgUH3jp8DuiH7xYMP2et1iQ4CDBAEm
hy2lhHjkMVGYvQjuFloRJTTf8A2HR0ON5b//dvQxaFBJHXyXs7HvlQb2Gnwv/Gzr
KQlz0vdTZ00o2OwSSVEWpVvLqLeu/r8qz+q71N0aOEL2nBlmGjEhKZq3KjInvuP6
vEzaj4VOCfhPwed4SmnWMpY7U/hVHhfWYCe89+o52VbvLMpvNTM3b09Imd9PxWbi
47zHKsv+XsOCQqp9aijGdcS17kT91WAeb40XjfH4xdPoXuabL4i4LIf9JfXMsVNh
k6fQxS4MzKPDP5PrzL2czvCzNTxjPxF7h4etMx8I5KQaLvDK7yYKycIYB4eZBkvr
tIdamdSB94MBDxGtOZY89Oaxw8X1jisia99aWCnnHTa3cdyrskg37F7DY5IQnoCO
rAYKIkgZMkdeFZP4LUA2YmtNIFGfFRqeiaRP72i6YE9+CNq3lKwh2RIFdaJbgdMg
dsIa9U9jHMH4R239uoU+gow9CIy+Tpl0xNYRo3VP5KIzlXcWwEqbgC+IJof/N4uX
Lky3aWenwWehiWsI44XayqYOUbDmtweJjEl28ueSai8x/oFliXlTG4JlK+YGv9AE
GNfk1BFQ7DW6ePfQ5u95YRGry59EXkD2/n/oPqhiP8HnodP+nAJ0idY38xUSdH3A
OkZUP1pQDkhGeakvC9MKBcwKMDVupgiCL91VWA0/DwdVLhIAbb43TRvaac4DkS7k
2ZzZKep6IEIjfHClSx6/gt3aJ0/xi8tQtz5v1HjfB+tl83sbmwFmBZEcSMoKmflf
zFfeB4noEa1LmCZCOgTOzdf50gAfgmVKCb8sE3qaj2i6egd0mp7WhONCHZbp1N4I
+9mQfAtsU8ehlAqSX9Sys91iGfAwfSv5T7LKdsZdy72Br+JWdWPsyB2jd9vhA6cL
7gt9ESqe6ayRRgz0HVLl1m3CdfL8wRT6bS+v9RIT6fvUmPjlAKA++oaVODKoQGTI
iRimZ44uYsgCxaZc3p+dSZ7DoIEqE39PMoi3fRxzO55OaRgPwD8ZC5kBG/1cZZwv
AbdZP7Zevgi6Ia4MqrLFljKEzAf6f1ObUonq6BOCfVzJd0L4/VBO5ILVJqWh3OML
thlj+fICXTJMhOK+qMbTwxaG+ErtI5sTkCD7UPPpWauQfgdddCmrToB0BuM39jMD
YQXC4ooVJIqwVVljAzbmIVIC1GjSDM6tKYCBGDZX0l0vQKI4bY340RGVHIvq//el
3fnApLiNp5BKuQSURgLFb7LblmH5mUtKFqZS3RKUdnDGylokHf0fWVDuIBBVPf8g
dE1IZ5e1Au6hAX6TkckJeS8N3EsoQ/UU5Mp5MVF09uBCn69PX8ANbrqXUs+yCVRI
sfJlj4+AW4wAJxck/+lDA7OxYMD+HpEp7qakhjutdCOHuGXIKmT+rKNSsf/xvJp+
jUmWkOxFKoFSEFNguyDsY/Va9qDnbHjPxuWb7N1fB+ug16nqdJl3W0BNyqAJDIFc
0Rlhnil15ML6eFjBaOYLvmowBx3A2EE9w8zJ7/gG9Gf+ELa4bHu1sYZVv2pSGQLS
yRpjWtUtQX3+/uQlsoziTw25b1DZ4mbHnDdsQtDRph8eFqMX2iaqwR91Dc7deylZ
HfXo+0baRoUWFMtWOkMFC8cXR6zbME+tDooWPzz9katO5FsIxUfjnXPsReLcW10x
l5afsoGYJ+NhjhCqLWvS3RpVTk//XZuZk5Uh3eehtzxd0j/Ypgjr0CXU957iWPHM
WH6rZvM+YYPchTHYME7CoLrHcAaG96oguFLR7cCpIvplt6lCZqhxVFX0uiwRL9nx
MsPWhUpDszz5eWD3PFTd4NlVnEN4tTulTzZzwfSfPqfbLjBK9Fqnk1wUDly90Tt2
2NX78HEDZXxFVMM7ayFPch5KL7yvF0JhzIh9En0YfHrI2TSZloGPMad49tBU3yyI
9BQ7BHkPezfY9a8hPoc2PPbqbnF6aqOta+W3273jNbNmB7Mvps0dWh2o4IPoWvuq
JnJaThrrkcID/ea2ZGq0Y/XydPYplJLSrLC0G17gc34NPoMTnTJRnfKyVoCNgOz2
1bW8Z6eNUI66O85Q7xymHCfd52xShCO6lPCl6wf0ATZ637jtwGp00UiUKx6wBR12
WqbFwJbqjtSh5U0lTHasqt5qFErpTFhjQra82VvsSTujUqL4HSDGKfmzPloTbGnY
feb43kaSgpKp8Bia6Lt4D0KvSc/yA/zb3uGqivsplpdsXsYx/IjbWI9jBE61R7QO
BEPYkQu9Qr6ZYcUFk9QGXmu8IcYLjvnEwx27YHzwR6EftJdbydRMGqlvG1GnFUOa
7AIZ85KJLZWQm8WUUeLy4/lhYF02XUwc7EwHiCb+jkmoALJEdIR970/sOtbDa5/v
cfj16PMMDn8atk5iYaLzxlhxXq6oKCbzRXZ3zGyt1cLERVUZIU5zz3qwpZ+F2h2l
pSAkEkRLep0XX4eKKLON2m6cAfYa4qZ+EoHwycfDmB3VfKjjsUHSVvbQ0IcbszEn
LJBYhI8IXd8c896jTyPCE7mlZUb5QFF3GthJKOAx4S4b1Yeh1kt2lDWHrSn3S6DT
IdQlbcFEVXDnGw66/KBnLFMNCiaROS8FgvDr26vFrypcNAf2k87XxD6z1IVzlURo
kxoC2kEBgJ+6cgcL8QK7ynvW6y4ED/FREpMJ4mQdFx/7YvaunLqfpqlH+z521RiI
K7z1A4zsgMMaMwZ25sRqATn0s6ctHG9KWgWSmGNBt8ocd1cmHpzcdY5Vqs/+d4Ma
vjg2qzmX1urFlS1AeAdC8jurh4SE0UpYeHvqm0QhbYE0ATtSxnMg6iwwBSETgAHi
IQ7810YNe539rQTSolbAlIU2r0LFfaHSzdYJgH7Y4aPmN+sIk1Awu7poqAp9ZP7i
Sm03hT15k9myQ0C5pfej47SoNADw+2uvYHhrD88IktL1aDcp+7VJSQHpX8Irb3se
5iJ2ynawoXpGp8e45jJTrp8SH+lkGaCjiTWiQRNGvTC7IjlrTakuLYvl84NKwvit
yKC+R00R0L3gllfQLh7GlPCzCieJTkjVJXTD6b3FrayXEjLkCNw5X9dtl8z98aGp
ra/I2LleEVJAGsek5pIxO43CCnAU0hOZ9qIr5hMRMDT5nDW/DsVny4WkA+oRmYSL
VAA9uc+0pE+fD1OQSNFjiMpD/pSJ9Aiu84/qSLzLmLupCeqsOKDSYZ1YONbIsHVC
+NvYR2Dz5ULb9FABzexAKI4yZ4IepVbURTgj9cRL9AfqFsxBauyyfnZNeshE/hav
NWRzal/olq/5h2MCN8PDbRB4piBZ1VmVw77GhmGz9btscslCOeKvvrIsMJlfdxFH
Ag897t0/rR4drww3J/+cHIagbNEiOtt5A6PZhSM2GBTdBMvlMItpPoajwb4jhpjw
aFS3CApKCdSBDa25pwgO6Pu7c2Gd77dA4AJIXLGV/ErKPtSj44MJS0a/Krp6y7Sa
xDH0KNFmP4XVd1S2sgHcHxTlCrQj1/dmpILr0zk9mdig88t5QF0m9qcmYVnuxQUB
ZvOuOYVpu0i52zEX90EkgvXdl7KaYM6g9TDTvw0/qP4Af3QT+2wlDVJRuyOvJ2gC
BVeDkEz+26MyelTIjuzS/K4EOppoM+KxHy06sxLCtlIiDTbZk6N6tyA+RDyn3mwT
BBQYlfIf0eElieU8ui72t2VYoTkJ5bnMN8O0fxsxgDVzZVHGRjzSOQremP7Vk1M3
QbPvxWtx9UgFjDJjTgzkmX04MiZO4ltGfkigsFFoqdnAnRxrLa724rFJ/53HO56F
5IPQTTB5XEwiXrNLZrtj9uRoxerGbP/7Xs+liR63Rb8E6OxnKjoO27qTSyNxqq5u
zEQ2KomqL4isiYU7ODRTKwE1d1g47iLe1GNOZ9957YNES+2aQ/wOvPS1oKeMoPSx
EWRP3euQFgrTeOvtlmwvuUCpxMXfsiwaUEaI5hoLvnNG3/lh6l4ivr9OfJnSUdRy
hu88gwG8rpjsgNCyUL1Ck3k0ABgYoq57M1JSQXt6l2f4snDkx31llzlrMvUrKUO/
T8g5YVEU5YwM/LEsMP55o3wXqFmWh6FiEwEVUAcL/7oXY3dacrE+M07KhpQore4+
qiTB/3HfpI6ygQmxT/O2ECUvyS4n+zDae4kKNZLMPmOPeB917hPCoBytd4+qmPTf
btDd1UxFRQnteWVh0/p83wIumLcB23HR11D5jyHziutbxepB2nL4AMC1rJsm7MEc
dnEYpWmlzbM2tUyCSeYOwha9dZQl2lbewIoGZJ0j1D++q5dc28SBlKJ7SCTDpDob
c4G5u1vlBjzARzvJMTBYF4vL8y+LlGhINlKvhSC0ef/Dbir4yZkF9ICtGKEFbUca
solgRBabEC6tiXHucfxG3TERXfI6CAYegI7+JsDIAThgF3wMeHOotAhGgVGNkNyr
aLGEoHzuUUnkVXw2H7wvaE/7XhrqAf5uCVbHTVttye/m+SpyUigplfL+CnPDipyT
INJQUkkotFzB5Taoe+VEx+BBEMOBVQ61O2v4/fPhXM2xmgBNIETlHRdKkJW7eYgL
Obpvi2MnPwJHRd9UwMxnLvvHQn83FndNx3EcUo4qXL7VSdV3qzVDjV3YONXcZItC
lqVgN4s2o65ejiylwquiRerSnWiM7z/bI0n8H2TKIiryR7F1IUQFuqVbqN1ps04l
5u+nXaKKWhaAvRZ0r2JBGF5aWO4Pq1SkztbXrMekdjT+XNgDGMnfWx32xgsgz2aC
N/WkxHpTSoT6YpvV5VS1yCzQJPjylZdsLQGAbddqhp0tispgxcOoikidF96Odmw2
OA+Yu/CN6KTHe6+XtNpR5ALTa9CHqXhakL7xLi8QuL55p56ml6wfUJTyJp6qaEGW
Pl5/aTMIJR6zRqOZDR8ptRuwpPtEubtt07eWQe4XPpkkX2DaSavnTIzrtTb4woo+
HO71gOTsEbFEYyRn5jmLcNk6c1ltYEZQX1kNMbD02Uf4VGtkRcHDUxwtVYwwXzBn
b/9ea1ad5Saie6inANT18CetIb4nnmcbV368ML9DQIIB6UxlfXXwdtnrABO7W8RH
ftBtZErV9eXAyNHfWFFBLg3MxMYC0IYHPbyn9G9sXSAEe8mj9j40lGoTCpgl+UmU
jm/sxas4MvqNpM4NWorUl/7wEta+eRGuOSOlF1gIZIAAkAng6WXdN2fiPdjeZnVa
QrEd2Ylhr0pBNUrcu1NO0OVWrtWCtj5YZbIPbb83QKIk+p5nl3pcpi6jMVLBXZ3q
gw3mZWSDxzzsTVClLxxiCLEoJlkpybOnj7mou4oG5D4a18inpuQGDf7q4wtJxfqK
fJPMj2bAtOJ6mC5bH0JgwWWY4urjRnow5dz5jINsa2znOYLVBQ7ZNy/kDX14hh2e
K+rjCxyf+h2zgqwn8g2cLY0E5SQl8Dn3uGA0eluBr/p95cYZHeYKTbV7w9kP5c4t
F/bq3MG0FeHbkCsptHn+OSJRFZ/eWmsjVNCpUNP+QrFXYnJS77oAUihEyvFcPVyu
/cfYr7JkMEb9EVk24B9/zDqJ/Vwg9+2TsKX36xRZtAnR4enzI+S7b0nU1/BiXNso
h3NdJEKVMGxZgFbg846y4HqVhuuvfA+6PzCFoeeg8N29fsJGUF9yQ/ewJhtVOLKp
3U/bEGiIgvXd+a0bhbGb/+n3beZ+kW31+KlBpoMDV72HBegTkMFOuVC0HN9m+yU1
erIur4O/7BbB1uYyU70tgp/j0r+5nM5OE/s4b6/S2hkwXgZtgC/PX/cWgRy8/Jv2
59uYOhvyz2ZdwGres6xH10glZNmqAVZntbTr5i1SVUXMLCnLf19wFJ1HXTRhMLid
sTZLq+Ek4NrVrFI4MyRaCl8FLEhGMnWZ+6EOcQnkZ27ihcvSHzziUhcMJh28MGeJ
DfozTXMkk8KzPd49Rbtr9WD3SiDsCVCqEDSNIx+K9jSAy+1TNvmNSpKyGFuPJW3L
F+UYrU9m08s2tkn/gUR1Da15XJQeoc9tLDNPJo+AnmSpivKUXCIoP9KOC1HkFeZa
aq/pcfDfF7AFa5HtnwCS7TeTdYBWQYZ+/Y0uknOlV5UmaFUkoWeRgUyHnVef1+/T
b7Jrigzk4UxFhz6PbyqRrWj+W5OFjQXBCoPg8DV2UhXWNzwb0TrIue1UQAL8FTHX
gL1JwABiNyjdIzkwxgUn5QJP8sP9zQbKOuuKmitRNpswCADVmk3nrnen+LNvoIbU
73OBUdL9DwmI+ZGzgt9yI7lWjLNH+QkDCRfU1xUSpkX0U/gfH3ksd5veFqxz18WY
7kUwX2F0Y0HVb/MxSlSGp3klqrVoa8RaDAm4jnT0+9SAOPI+7CDK8OrcxIstx/0R
SiajW0U/0499J1+v9lP2XB+E3p0rc9Cb2UtKfVZbhs1z7x4XtQerDuVRa2qbEP2m
e9fg6VYhMWv768FpueqqhoVISAKTHteglr6bwRMfD1QUOO4RZHylkfzbSwWMX19/
APSyEcIUjKEkHSmvPGqJV2a/bDr5gWEVbJ44CzEM8aRp4yFEKmsm7HyHovwnC8zY
uVdenVt8vIHirPf8YxiMl2CsOU8DB3mvjUb099LgcvALnFbWMMem1OnzUOu0oNo7
b3BdT5gqtL2SAjf9KBDgZhYAiMFoqk5Yloh80kxpCklMwmXXHk5JxirpdPFfg9bO
J5uyhrI/VWPi5n8tFgVjMe5Nxz26byrrRIXxypuAzidPE0Tp2f2AdpSohUKnBMCw
QyWsfmcPVp5BwxpB4UfOse+AgfIJe7htt9tYY366T+W2T/FAIjeWgQ4W7w5ziky6
S5Ud1+g2A+QapS4vudf+EyP2l7Hp2C6UTRw8ntyFXR15clxMXQyhdwpDioG4c3Q3
GQBohzcBgWla9m1FPTYEzMTzw6Fbmt5w5dmdaaKec2NVbm7N8d58ZXhADY66nGio
9S+NUCim1U7gpim1HqyOj/uq/hhTeyB/LAv1msMZrUaSeeh0el/nEQ+h5yUgfdGD
5+af6w2m2N1njEtJe9cJh8V5wIV/pGqPgN+nUA8PSxfg7csYM/04zGhoX1e49gNP
Z8ytjohhR4FiNtdT2RnVsWl/XqQJtdXRPlimOtsgKXucKZeOo2Er7NgQFJo4oKzk
JK70SUdxLhEer9y2pFAeWBYkdYe70om0rFADBJ/ulu+PUzYpyurDa1deGbqSW5r7
CgKx3ZCJvGM7/Y9ITCtAt2VyQaTgwoLcVucxil2gpvbU4ENfGsqt8ATXEk0MC2Ap
bI5bBTqqvPLpw6iv9ak1rrmq1kkKDUII1SRMsX+/i8WjoidyJmMaAbLJoCEL2aVP
4Sb5NWZ/fm7ezlS8qZe9LAmbYi7t04kpp0Do9teO78ENOEoj9jg1DTM+Y38l+p41
mXhSzc9rjb0xE4/IhSDLGRXJF8ViHZfn9c5J20CtOG8BVs4l9IRkpfSi44a5t2IJ
Bh2YimpCZyhq3KZVaPrN/9hA5Zup82+5Pn5lsC4LzaZOfa7AS+/zRzAfEygqCY9/
NgrXxaE/63UREKHyy6EjlpNuqKDXjtiaTCZlsgGP5zMfCcstbUurafj06JMoVTVC
2cZma1CS5ajY/sx60wR62JRc/8qDMKAcuHj7pjhg4gkUWJX0KsgaBwYEWytIAZ9I
23Ftc9+MUZ1CBSMKsuQBtkOuHpcqmURAsxry06RpiqXp3CidcRDZ+e2UCdEHIZU/
u6o3gm7MBSIAMM8Se30eBtnWuaANn0nBioNmTzV47SPdSK8vVTYyJUE2eNyD8+XM
R9NYnHeSMASbb7CYNGkDD9ZJk0tirzGKteGhm4eAOcx1EWNIyDawReVnywyQF+fo
BVeAnKuOPNQCSmBKjt5CePAOtyKTTs+oCsf/tz6g7bPrOw8d2qDvG5QMKDT+GGQb
GVpcVxLJS8gg1Kq3wcxQkJ4aSYiX/yfQvjuUh4WlW3c9rxO/rsFAUXs1ePUtIOzF
Yy2AXPyR2NMkWS+MaPIgHhrIFoU/fXOYiwMGHqiD0pJj/bc9YJQl0S4O+Muoyxxu
rRl4+HthbdQzdbO5tDVuwa+j41rgVG2YP47zXQQjcek/fIqzIkMa+vYeV/6a1mN/
RqqiRKgkF5KQ1wJR5BAoyBMs0+RNQA4ugOygRHz34lDeFS0psTPoVaNSx8pVBD9Y
SGzTX1+mV3hexPHd34bZcSs7EieE8tJAGXu0GeLJW5RJMd0YsFKrCoCAjoNxXkfc
dIY4Gce0+/LOzz0xtMfI7+7PbpqKYzuWstkvrY5Ay5ZhM0Pm+yb5jngprrs/Fydj
pOmVPLtNDyEmjOAA+86vxJluCvssKHHuIGGlZwyj7FDizIIPfd0RZE4d0stipM7W
ccbV7OVcN/wU1ea6WlO33ICQlN4m8ZS8P6DWvscO3ssZzqiIQbbQeMSHEOeQcZeF
+182OSWVhDVBItfhzQxA75ASzpHE/f8ctCA9Q06EyoN49e6zv4BXkFS4hoPV/zWw
FdVJrcFUCiw6bBia80cHNDpIdrpHt8/psff00Fb1PxZOHJnUAkK5ZAkTaY3PWoC0
a8hdKKncuWKfJzKB2NA6BkuEAQAwH8vfon02ogUlU1viP9uIit604IBhMhFN7NKg
j9fzniI9pgzIyYFu0iXfls1bdOR4qI0+WlPsDUw//LfGOsBeCtlec+X28tIuiE4N
aetKEUb8mAHCg0Lywvpc/DVabXSuJ1L8a9+7pqk4cLnMqkZP5QDEZRFUaDx8NlCs
Qb5IwbFlvrjjunyMl+uK7gK/D4QppCzZF7PlX0Z3MDI2s0XaLogrJcc5gAQyM+ZJ
Tikh2/HA4AGaXK0mvdx3qfSxBnIqPa3V13OYrgmKkkRjrZwphS0nHslVuxyfuyMJ
j0GH3Img3i0tyKOuwplJ6dqDy302OVUubMXyaOTMh5Myqy2u+SNSYX+EpAo0wc0s
i248RsryOw1GRVoiZgiKFT10s9DnEjqgE/XY5D8Fz5T5DZb68JxgFflx4/Un7+Hw
VXIgtNRh8JZSOVtmWoc4ZoxsbL6QDYH37XrXMh6ZLk/5kVPkT7UfNtAwVEgMtQXz
PZ43k+63VP24qe5rc59WfP/0NCSMh0/kdBgz1AEMRu3CLGOQmCT8Hpa09nNo7vfg
YvqiHRoK7Ng2xU9zUUc4Djq03O89FjFiZs7goAhYU1kWu8uvMWSD3+qaRhDsKiR2
XPhIwfoICFbLNus9KtnWV1VCtsvy89rLeMJ5ywrAEN32PLdOo4W5fRrV4xIy+4A9
/ZzATNrE1e3ZdkBjob4xsPNISc+4sRXOHwyD1B0H1CGYmkUPfQGmqNf5WgVTpYCB
Eqsu0gsKQtUtaGSyot1Vf92a4GqTeC4vr7v6qaB5/T19YgwHo3fWaof9sTa6us5L
pKLfERA60bG3hLV0L/HAK5IRT8zKEH7p+p0x9HSaOEVFt6OZ0nK+uzH90WnTHXWr
nBrVmn2bNjlZMXoQ1b8bx2W8QChKB7uyvXlKrjLnDa/nGrWwpqPsEAY6BuT1BdpT
ltUa73xzIJa8qf93vyvHTmUrOeIZzoEzY+XCaekhXWNMQbY7PPNBjt43vPQ3Eri6
NwzWXQSo7gGwcjEaMyDBk/YiU2lkVHi/2y+UkJ6kIYJ8bm8TQc4Mnpx3bwv3BZZp
FosuxSE7TzJUFLtHojlxWzSqZ3Q0GNKS1YZx0RrukRJUBAVZXp+zDThnN5S2vuCC
7WYGJs3su2mEmwn/DvSmP0e6Gd9diqxSk58IPujf+BpAE/pq/ILqM6/0xmz+Q4bp
Pns8uBwlJ1oqPSzapswfxjMETchy9M4FnCNOXPrNIHElg1S2/xUQQRlGXCXS7RIc
m6H4IJ5tSfcT/gSFZj4p025LRBGqSksykmMHCIOyLjZUqEfCXWlyzSGbdPh9/oWk
Fmny2gsFf074Z+L4eadB4kC0RkDwQeAnBrR+GgKZSSpaJJCUWjnz09JCq2Z0Xsq+
aiQGhEyztPkrfLwSgVPwTXzlsrlXFkky3p/X+DYiVXuTM5OkhKRrVxi5SQDCmLkd
V0FLn+kGGlsVOmf33aey0GiX9SDfiS21VgE1Y7xDgRcg2aECa9+aKcb5LRnnV1b2
eah5EywruNkhf2Ve9IWdQKqnlR7g/StqV+LelId0jOK0ij7x4vc+n5ESaHyrArnu
shugbz370KF4FksCURz5QxDX4kWQbDvUNryO8CBvXAWpOUv+lx60re8jBaUe4ZiL
Fy8osVjknievt3wdJiAt71gkokzDdH6K/NV57XUBMCNc9lzohbKUFvrbRhLGvVI4
1hi9AhFHbMjLaXEMurlvTE7a9zjSV4R07j+X6ZgjAZ5thmrAwhFWFdQeDoRd16Ur
Pn+ocdWxPNnUZH9RYtOzH1Gd9TsD8b8mUtF5P/QTyMnTrC4pqv0afrAu3WjSsX3i
33+D7UjiPK6ct1mYbniuAPqA0V0YtEAy19PJNL1grYbPtoYXjjpwPBh1LwsF+PeU
wNEd5r1T7vWJof3ACeibj7DLFUcep6H/4hpzsiikVaA6F6+jzywg6lRfHP0W8tRN
ZO3R3qjZQeFsdIbm+hX42LI2CpRH1ysSan7job894XS+GTMumkdEg/xMxrMpBObI
10NtvjlJqi3oJ7PjKypv6eWSMV+jv3wb+P5yMnpGFFmyCct55uLgTZyQp6z52I7I
PeZz1wJLD0qtPFEG8GOgAbXYMiQNCV1YgPY1EbojkSKhp3WCMjKDmitKABe8+S/Y
E9yEN9EgrUZTg7Oev2dvKV04l11eqIWt1pe44fTE+Xe63XTXXGFftSjxPcWl5OUx
joFHkS0nvPqzIpqgWeK7OQnxhRyM50VzhCAxH2P2aL2dtq9xJV3+aXLCokebxCpx
tzjNxdQZjUXSjocPANIIRR38SW0gcTwfFI3ZZP1I/k8uEgmu4uVo4VOlSxF4LXB+
/3DJIGPbmBDVrp8EAfQrJ+3HOqRX31OzXDIbIBkM4mMNWaRec2q6ImQlX+tUFhKr
DKAij9zo0lpPcyxgom1374aq2bNIC3HXujYADQy0MuWYNKxFRCH7MRQ/QiUozQXF
K8b49ue+bd5j7R4GNmrLuQtygdNYo659Kz1tcg9AUGrpwqD78IPtAcFgxCgJc4rp
gHOt5NZQPXm1R2LbYWApAILFa5cAOsrcWfn/7f7zhcdV4CJtrxRNQ5Qetq1UQqlJ
KoG/rMlzkFH0WvWED0rSj70tLVI5L3K9rUlhhD34RmNWl67uVVGCWrVEHwM+L7jc
y+jGKAPcGjRFYIJddvPoI9Q99BjitzOneX7k7XijLi4igY8tBnABhddykPFLo1JM
vyqVwmViMORXD8jucPzKVjNcw2E8l2BK7LhKh9xYJ/5s7dI2oigR6jqxsQ06lYc/
IYTanmr8fGHr0O3FZVqmbm91u87ADsVy/fT+aEk2GwWGVA0ouTCV2S0JEY9SfMwD
ASMzyCT7YFx3TPzDuWKGGeiLm6nVbHbNXwFwpU94cXKZIhi691mDS7ULmjryEpRP
Qg01U+PKNv26f4g5vID7NpBT7i8qI9Qq6KBEeCsWHd2+tiopz4x2tYQ2zNZM3ks+
g9Y24fR2SIjcSYNGIyJy3dtpEptyC6xUh32PBrAJ6+dlxzE4OGPuR/j2pFwGDnxD
On65sCmvVA/DGv9EinWGkKe1SAYhQlSCzukuY2FsQ3yBuBQAEqSfCnaNXMHwDtzz
tZBkhXZdo0gKvH4cGWDNKG7BnmHhOyPQHCLQhpd/xK8kU0ZSRuNIpd9VT6dleooj
NxpExs29jBYitfweCy8LhMmkKgatui/ZiIbCJNM5LBEhlgUYIu0r7qQb9h9nyR9B
V+1eYP+k786RwpMAZ93TKSD3x/Yx2b3jJxu6C6RipYH9q33WihmLM6aY0ftpK+fl
u/tgBcOUKpq6RFMxvsZ7TjK19mvJNEYgL7XRmqnMApx+7IobeEBIObQFsl4JwTrC
Qq6IMjDmDqFdqCiXkQKouDUF5aZi/2xBOeezl+jgD4Uxkj4SPRqwW5v+y7uIkVcF
87Nh9JQ/l9Phf/cQZkcgZwOhP5oDgjTBORbEGimorqMOgz4xgLB+/cla4OGaoxZE
X+sHGyAcqj23dh6lLkCJMAfOpjjwJaxK9MoNabE9kPUwBrFKvchoHwZdjq7b+N5C
Fvd1c7PLANviAid6wU4E+rP08OPDIch/X3+XX4YSFr0EZJv50ScFimiLbgCMvpH6
ZcKZ//54FKWmu+KHkfbcxYXnacPmJFXq/JHbgBETvhsf/IqgTRB8rE2ZzZUutHzx
dNdu3xRdIitfLNeCBfDJwx0kDKbk+NP7rK4h73qWFSn44LsBSkHLL0CFkrsaOW7h
3C+rLBPC9MS9N/ROHA8Q0ulnATobtrg9JZvt2zkMMjjknielg2w6tcFPFKlAjgx2
OyKOQghqP1/K6HnBWgn5vcZRs9BB0p1//jkmS72R1cRMVqkD6iIW8NQwX2HuGVVh
FXGBcuwIePNQODsmVFVlnoQg3J5Kb6pVR/ZxSmGIZ+/NvRN8VtQSmWt1Pbr0hbXR
fX2peqOrApNH+Oh6NG6lg4LfW0lD0YFOiNMFuimAdMbuokw8c39xLd3To0YZmFkF
+Ezg7SzGHss+gnRppPKBsrc7YGxlNq4XUFbv/gr0BdeGwWhGkGTfhpilywWO0/8C
pFsQJdV0F4IwdJ35RM/G1lsQCwOfJH4iQeay5dQTCdzxGcctJkIdYgHTERje99un
xhX3oqvwlbn+eZOUhUpreasB246IbHpmUC5atKJmqmmzaelH8hGnBnjsAcCVjEwU
ec4vmoo40UiXGEQWjnEznC+jrhlO7/KLxxjZnuMYX5oajhTFt5COSHJTazCfXVyp
KWWXFyyhi3wSVds5dIvF0usCjnmzGMQTuXCawiqNeGvRZUhrEs7cD/LLoZGvrsoM
JB89TdNn7dvL2z1niAH/LPCipq57KnKTUp6Tgt8Dr7MCvPoKIWyw+af3JzAnDDbw
vUl8CsYPKhDVpnFj1Wb4drdekfrB0IPluaYJju5ds/NAClUPxK1Ya6V7hKgPZSTe
/BvlsCK2llcnhOL08DmTlxqEKOTXb4JAkU3Hh/6uRTEua1MeJnMMolt2ce5/tSIj
5YBsNyWJQ0jo/sZy168kJGE9mGsM/DEj3GU0MJ2ogLb5pwQtv+wsnURYg9Cfh9Oo
lCVfhy3b7jlQaciZhBBM6mDInEsogFvdw0p3CKMzOne79GAQGEK/FCQdig5S1wG9
rTUSB1lbxptHvO9qlDP1CscTs8HF6eDSoPxr1OrqdSCJ0Qyj15D/kdpoEm5hRt9h
gI4EEGLeZ7AyZCbJgIeXZyag5f4rXh20X/ziR1d5GmSvoppvrYmn7dwmdj2bvtjV
2cdjzCcb2y91jOQzYUBCMZTLdU7+hO00XtqQZbHjFh8yD60OOkbiT8Fp70TB/wqx
aYixpp136SvDsvYqdHi6m4agiFIzjuNgYA9HwXXG1mGeYjp73qpoUJ1H3bVn6b8V
ZY8WWEfAu7cd2M2xE4xD0lQ9aDO1NfLD622PE4uLW2BqJphu9xHFCjEzUVtZ20SL
W6E5B81edaUe4z+D2PnrVIXmypy8q/Zde5AmObjbtBS36NcMAQ/UKPd/tIYY+2u0
oGpCYZxK4vYauY95wbpaM8iEJPEFemD5oublbEDSqm2yXKVHJdALMhtf3EeYfofo
KRgjZxTNnjgsO/QtEPgCd3gCkLYK8kw5XtSoBToqqaAMYjfHR8t4hUhPFE52DfWZ
F5AVooOrxfn82reb/UNqSi8DpJM6vuq298vicbO3HBHi7U4pZ70r5cmj+wZ6vksy
fMsDnNXF+GGhOhWnk9Os9jLHo+WKucL5pQf0rIyH0Fx4pyQzv3UlsUnDcRiN9Lsu
M4uUIWc3zgLnHDiP0qReujXIooxAmf1gMIHRLfRoXtaxYP6RqErUEDw5Vu2zdR11
QfQRHSVZSfCxdg3sVxfBOI61wJjAGJOZ4QxoCFLd3VLC18ptqt9Bj1zLydf/Z22+
Q8p6fQHLnLbuEARAB9sXQAiTOLuHW5q2fJjqpIyGc4L3sMU8gDJ9fhMYKzShMIjs
zQn6MfRwtYj+kDCW2K04MTBz3TjYen81Vtzhp+3pFBFz8kF8BBx+ZD4slPUqxZ3P
Egvd9+qyJagzoxEvD1snx5AatVdoXVduTB+R+wb2ykLKodocbA+qW1zi6fZX5uLT
y1fb0UAFHwY9ueddRMNIAF2FwEHuULAkJNGSpabc/p61m88BDRDZ12swicvjKTK+
3gdwwwG/S1ULgf38h7HMVQTNogd1VKXkfw0ng2AlOLE3RoPX8OBZgLf2acr9NhEI
OslJv3JWbtpOZ3qxtBTOMcLkoXR4IhFPtr11Yb6A8Wkl89WDVULF4HfVfNUBlq7i
8FxJDtwE0RTCQk2zUUrZYdMpelO8IIuD0AkZCsn5P8gVU7sXuK7EHZJjWDvZXCBA
PLSxtCDKnSW41sPvXb0V7iaaek0vklgI2JjvKCi520YdBj9EdQmxxywaSemAL3Bn
IVnXROAhXnthNhE2dLKUXchR1TKTr9NHnNpimjqY9Rz+Dl5SraTWYpRDhcZ9W12V
TFa32U6FquA++d54bplEjM04nvFPuSEoh0HgGbuvI1tgd9q9nkdPgVNqRDJyIpjw
ebUdXe14UxaKBn7Rj9WBi8nFFztQ0lULRmBt12Qns1rQuqUs2wjYy9gu5GO5yUM9
2qGAH7NITMAnijIvBnRa5wGrUN0zVwL+lhe96vdmhwawY0uAKW8w2ogYIQt8fWzE
V9m42XItEy5Mrkcb1SEphyBCb4dc6lKAqBnG4W+qBIAo2uX/2OsnSDZC+MNjFlVO
o23yt4ANIDRxwDvV/qpAZdgPNxbBxjgrtVXdmu0pGs9+Vo66YBBZnyQZH72PtH+e
fmWBYFrCPZu3Mrmx7Pm9WV8WJMNDe4xsGbC8MUAq1lbXP9I2ViUwdAYtZc/XQwRZ
yQ2WhAZfHlJWy2hucSAP74IaoVlHnnf1oJfIGywIQJOHrdVApVdXBZJccYzfF6Bp
5Y84pYxyRHLlUqu1oKmgagZNsbznDueUXtMINznDTEn3/ZodrIzVsHfNjxzZ9eYC
jkI91+LaJZ+mrygYgIa5dCh1BBhKQQhQ50p4+vDS8YP+EDHOOLbWqCvcbe5D0n2G
5ZgeINCH8g2rTCULH9vkEBlfdlFL5ma6krHLEa+xIxYxFSZbHYBz/ih04tm8P4/E
InUO51Nx0hmVE3WbBTjEBFzNIjOL77e7LKUwV3Cp17PyiV1FW6V5gES8QEFLTp2o
FDirLJdUr0lv3cSL+DtHjBIKkH+xQTyZVawtS3pQK5s2gqiNhicFL483mM7Hzbxx
g/bCTQkqqn0tqe74p/VFUI+ay0MhHY96Ll4wfD+WV16bIZcQSHcUz9fF+m2/E67o
cmVlFA/S3qiPviobD37LFuhbMsHZp/8xLCDEhjnHRctyEQ139cepkOMQw3sFPzcf
BXwssx0lawQVox5uRUlGBeQ/2OgB59zOhhtXMHI8L4zYfz1sN1IwVY0m03IxqGf4
oUEDg1WAPe7bhxK2rXEkHuJRr/f6NaaOn89J/D9dswsF1Cq8edwNNKfUNdHNHOWM
wY/kdSFdqtrqSziWPiVtbELvHU1LbAG7UPlX8RJPGjbo/tdErHLYt3PTOvk0VRM5
HX0DNGPPrUb6ezatMHxn27Q/e3TAY40y2VHzrmhwWOkJi90RGVpPDYpHR4gWQ4HM
RuJOEDG1T/UkaXL0xlW+vYKdB8+iXavmY3m7nGyovKGgV0ulmvVpa6eno1rxHjzU
BvkxNK9I7P+f7bYzoXCrWVjY5Eq1I/IUNWLJWcx5qMt9x01blscVpJdABMG5f7IS
WkNCXrgcqS6saEkopEHj9s++nFfESx75K5Icv8o/1ZuwJMk87d+XaUkXoRwmin3G
Cyi+K7aJ9BR15/j44Fctr3QoHifJZy7+5ODE3/9O2pbKPDSBae1Jlk/7qfbG/vLS
H0IuiDH1Ppg02KPFS/YeSvGy2qk0RlpD4bL0pYMIL5vPOsv6u4J68ABAXDF9JUpL
3KZeZg9IYy4z1hcEsPCKyXO7TA+ajMyKeJ654fUZZUWVFEk4qZIAgUm4RGoucGNa
39Pnye3hX3btwOQiO/Yawc6rUmlY9mKHJTvJuOad7MJ1NRP57xDDvl7W7jfT3kfo
7E/DgK0FvMm+0W9Xq6aNLBCPVaDINylTIVF3xSfeYHZvNQmQOplG2tNXC+h7QsFt
HQ1d4Kh604G28qtCp2S844/KgIkGepB2PxiKTH2N2eFub5TJJRashXQMlZuCuHox
QRklTRKK6I03oTiXb1N0rwN6H5cbbyEXgRXZ9+WjzO3IbW1zW0h+37oPto5jucfw
XuR7/G8IOAhdscafQiH1Chc++ysGjKAXib9NnPrSYBHfxqTVmuP/eHnjI2ayePF4
oigZ14mzfn1kcueG1poRFHYwgOW2DJhHCZwYR31aPg2lEMAFVciVLbnNmGLSVLD/
llS5/R0NeE+n7Fp3fCC9z/pHcj1JGV4UrqII+Fcd3D+D/UI6TgzQSE7amzo/tGQ3
/W9b0T8f/E8YvVpNwga1h7lRv0GU9NtCxPj0WvnxXTb4jrYd67NcAIsG++AB1+YM
TEXYx1VimhcqMFKp9pfQPI5Bc0zH0Wx+Z7ui8aJpJgFAuPV8aGR9orQz8RG8MaCf
BxS48/hAwPpSymjV0QETivLjpWXUL+Q0y7PHfzLR0wQ/8sONDJlKSwvrbA3/0djh
z1wxKGQM9R/dsVtu+Ah/TtQVDLzaOGfXPKH/2F9xYCUoH2rtBzh9kP19YL44QoAC
Vz9KoOBmi90OTBhmCZYJzmjz5bkAfqXtlGZ/rkoasUw0Fs/7LWunxu8JWNj3nPil
MvNTl42Pr9yyQvAY3E9mszv4qPJonsVplMSXtRZS/YGJCVgpFPpdUnwUC9sT4V2N
N/LWumbz95KZcnwXt8VycHzjwVVs3O/2YWCHuMJ8cGtpsV6jVrZ9Rx+9KQa/tI05
0M74RozBV026fAfhcAb9X/pZ9CVWJ1+jlHDB+JCr3JrWAzJgGryS8JLl7EyCLnsH
T696jHQr9M4RcSJaznDSgiqgiVysFm4fG88MQ+LoR7C9aD9z/LTawKVfMyoNss36
riw5/tloTW59/pgw5X/kmOBHj/le0eRtStc/Ygei0DzwXAAC5x0q/MKkLn7gWNDT
2ux4hB6iohsn++lmKRobaNP89J5E6VXG9Y7kKDuySAhfEFTpNyUKFghGYDTMs/ZW
F13wnEXhv3IcJa/QqvErQKUwfM1Mo3yw//omCejNHsWFZTXPSpuMUvYKoz85vvUC
vQzoCTgllzbCaN6HuuG6OWAmJ0FeQ9nnrpqgJHIDumHlgD9TqUmeNqd4Of/NPqDt
MjVh98o1PzC4nPgPawN7tlNbCVJ8lTC3/mLRz00k3odmQ1Qm5hBZ5Ey7LT4Zbn+Z
L4dGy1PgI+gRCrjpSDzHQboTNTT1H+g1F+hsW3x15fIuICwTY83usYHg5d8n69s7
en9UXh0dvFsOIR+pA0R8YguA1KH3VpHFtP/coKfAjWN59bWlYbTNHo4wZcNx/PcG
65Ee/VIzRvqkyfOpwAAj6+mrd6pfk2yuYrFOLBmbcK9Ss9azaANeKjLHRVvuM/a8
egGMjHdpAacUbPM9PnFY/8S6DCcdvaaMzlglOE9D0ccsKLyCgoKTfUyOIb+e4P2L
6gJddbZF5UcHNqsckzpv6y6OSunefcFerhg5c/mW/5/WEZcuZTyf8tvVt/vaXwOc
qCovtBghkMphCLqVr+tOjf5Eha9hzsLBH9VN8e+KqDVyGJVLKEmX9UzOt5DQQnpc
EMMgjkC+Ov/mvlst2DK4VKjqx0d5Xh67kRGFROAlhniG3vHjg0h+V0tJuxatwdlR
v1HuBqlAWaR2RxaqxHmvG3OYxbZJdPmOJEnmZq8TNpq5vfeSk+Kkp23qFjr6Jmid
FzOyK/Yz8P+sAapev8aI9ehteHTa3EcEAcvMPIjZFklywQ5sfIH2UypDiEYnx5KO
TVlv7MhwEXZARjkYwAf14tnqSLsOYqA0eJCb2Hywz7xNu7XvIjLyha0Rc1VcBGrh
PlQYtLms8ep3z5/yRqIIs4Pt6j+za7xYTcsFGVdRsCsZcqLc3FdudXQwhg7RsLs/
7fVr+gE9piDSTBEoS3+6kV+YInjGFv/yZO42rBgLK2/OiFAnyU4WrbbcRNgEX3Ni
DfsW6N7GbKQnmKEspUMrHWhD+CWnMPMO9i1muU6q7mNy/GYi3lfnGyo95c+XkZ28
oMCHQgCgZw4IwPwGfwk8BOqwzJ8rDbyrKRzcz3VK/kcuypkm5VYLFbKAf9ByGBpj
H4bzVdjOmeTPICqKu4rYuefR+fFOcIO8ZSuYTLFHjJ7TpEzPCnLuzK0/ZhBhU+zo
b5fKiLfF8fWF8hg+RoyUWo6uvJ+3/Pm1TtM6hrW3wIzlLsHOZjQ4AzTeKOqDX7IW
E87uCq0UBfrRy5uxtxel9+HLdJY4loFj6FsS6TuMl+b+/tzPzfKS5+Ny8V4sXcOW
0v9XVoOH9k7pnfAXjqKGJX+EB2o3EFUId/5vrBa0kF/b1dX033evtvdRr2bflA0l
Itcx/jglJb3FB0glzUb31WGe/yJT46mDLY0rpRc/NnkzloJvdb4iWqHaJEaJSI58
8bIwm2QioL624XNhNSk+Spp7caQ7elBxL9KPqoMxmjPOq+e9ghRUUiP3UYytLIIF
EBZAt+QDUvpXWU975xxhE/RnW1xUJ5BrVI2XaJmk2NfKkIvasVvqBkMubQ8kssxQ
bcj0RXtS52/7x7SA/SRSKcQO1hhbNAs45AEXOtD5QrDb9emMRfhZ6urFLQltmfDl
+lixjvWydtHJs2XnGRIyDyKGlUrxplsppuAYu9hEE5/8kA3waNiGQOFCY6YkJ78S
hWdSW3VUHlcPvJ4UygHfaCvSfCiIU2knER7YZ1bpYBuioQOod5hvw8DMmKTcn4MU
5qACdKdCUtOY6pAqIHnLU7BUghGYMeLqsuVwgzDd1EStyWQxM+urZNZy/hDf0XIk
mpp0ekHzEFfytYPTxFOQSvi6L3Mz4n6dRFiAlbgS5zpb6sV4FRslLka8zis5NWZ0
eab9Ku+BxsYFnuw+sHnNeOrJncV62ipUfWhLsnD+HXZFvUqHsyvCl5y9AQnTd8sy
`pragma protect end_protected
