// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FWsKTL8XZgEcjTS0HsydjD0FdXX/z2t0uOKiwCVmOgrdeK1glCsSa+QSJ6JkYKxa
4tue1pc5p33TzgOL30Z9KyiLe88LH7cHtSbseGKVqxjUTQE7C0JgBBO1z5oBXDgX
b1NdbyvcMiSRCnQ4OLGEAhhumY3jmuocdGLqSiE5/QI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21680)
uOyVffbvQmXi4hGpN/CKm4sS1xmWvCZDgl1LpKKiuR4q4IaPnJkV/zvNrH3N7QKN
d5iouKmJR1Wk+8jvTmyJOkwdp21FNWycb6NWhw+nHBiXmJeN+x9atm89qJNNucla
fUht6ueyDP5hmOhudY1vL9nTiBp4Wh52S106bkwQFc/lMdtucPcgD3boWCz+TA/u
oVPrUdtUgMzPagZ1E3yZobFpi6Vc5SsKQjSYCidbAxC/Mrca0aqAJUPLLqMdsvIt
ltZ0mGQbOIMuYI94PRzEprU1bEOV3ZpTXeY41DuEAxHrrXO3IzFM4qoW1MUGuGeN
JbUi9Wan4SQQ0i8DFiWqBDOcNkdaPcqTxtsn+2xl5dqWf7kZxuwfZwNDj2Qc/IUr
vh2ipMb8Rwjm+nWJ8l34ZfsXNVQaP91XGDmpDyDbxSZJq6WjMrzJUv3JkYcoGLmd
wTd7Z3/2S/URQ+gBqzrXklq9tE7PejFxRG8WcmxoTfP9cAsW4l7/DbL7IGhBXWj0
5+4JxEFukHdvoyewLydVy6lboaTkDJ7V6jj5Q2DPP8zx0rpMvMsMa+2ORA6cBPpE
AB7UCpQ/VXK4JYgxa7UwU1rmq+zTwhjeo0FXydmubYGFKw8crgh1WFAjt5pdN+LU
FePCptJf1ssxdzSo6e/UprjYrAXsWgHcuIod+GQ+YJKpAqm8el6g+RRSxVvrIb3y
XYm1uVhJ0bdP6vQp8l/GyeX7hgNB6hwLWkYSsh4YESzv8qQoFG7KyvLYSHYEoKAO
o3fxiAcVnuZchE66I9wh6mMYGWHb6d0iS6/hdDo6HWAgtNmHyDdqqu0Lmje0VSXV
i1SGcw6ncEXvebXQszsg9BIEAFrmtZZUcg7y2HVz4Rq77gn0KNJaepzJshAT7Djo
UmcL423JuF6/cIbwUacjagDuL7+Hg08HbSfYTHTXfZyPNB2/Oc6lIQ/wWIHCmhCv
FbkS8l3ZsT/LBAeEtOchx2GlaBwpC0Z5h6yHr5ZHIA7AFLIrH78clvcvf4blguzZ
0/eY1WrVV21D4iewHVLPGvVTpaki94tUsizCqw//T4PvJK+/SiHxe+wtV5bhIT4M
ft0daOc6vzjmcWMOs1Z/BB8SE6OcVbYIElIHfvlB+oeoDZrJLl3A4mEQ5VcIUQa2
3k2NUnHHBjO+mwynh6MVw1XpbnXd6+j0HKy8922QAC/xHVYa8PHwuCtl3Ba7GrsS
ZJ6e8t0jhR+XbwDH/8AOhVGHytY9RiZPyNMYK3pd7dXWi44e6Tnx7DbaHnFs1fF1
GX4zOky5slzUl2XvcdBI/yoshQx9hxd9RsAn6JKQO9SdY7pnx7sOaYEBawaIF1Hk
qtuKvNWgDe6LsmyEhodmr8wc57DKGaeqQLpuBqlV4iAJatPA6fx1VrwfmG9Yvhtj
0tjWXM+lKg2+Z15E9ql+K8mRg4dzGMGqYug+hL+j0JOmUCucmdoDSWocfe/T1w1G
NX4Kk6WzutQjeGJE9/cM/QRqKK8pb+vqD2+r/XR1EqX0p6Y/3gjhhdVySSmMztqp
w35xxuCbNWwfkE8PeSRnYo4gRGJL8IzbHmrmXkzqB3nE3VlB9g09zNk1XcsFwWv2
0FUurenIqBGXVzdg3XEB6EzTT1uC91IrKS2y8oO74EKNC1BHLNdI+Ex4c6Oy7VM0
wIbIoUwi9DJF6BowqnYUyn/KMa+obhe6/3wf74Y7aqVzgrYqvdltEqNqVx9hA9Fc
kaTuKkY/ZcT5jmtetseq6zcSUHTpXjt8mLzyKTUAmm5eQCO22HYwkD55WNNJMJP/
Qh8brJHxQAO/yR6bSEYtuyz3DbK84gYD1XcoHA388dKUxloVRfoC9/jwh3z5DHAW
zm17H7H8DOVIxtg1Kv0sik/cUx8QHIuUV7m4Dgm709aU3mItxf1EM+u35Zo8LU3e
InI++mwT76VLV06DhX1wu0qcK13c88wAUcbysrqJtJ5QJJpX0Ym93Jz8eWJdeahx
sW1Du6CQIWkD7h1Vs6EfJXYM2JT1Tk/KjNH4BYj5a4g/U0spv7bwasyRVToEEQXM
NMOXrTjLN8JIb9Q1ejKrdXCk520tv8dsGJTx71rDFCtJpmbo4hCAfweWlf5yHrWH
jW0ZZU3x93DsKdCo7lffERtsB2vmiBjJY1lAsY90clHdRkoJfkbnV/KVqQHEsyY9
Jfj72vp81BPDfqFsBwPHghZQQn/rhbPeAaZH4fBI5zbWFPdVnjz38WMYTDE/VhF7
/NNyK+XGDFJmN66eE1CZeUb6FFoK96V4OWpuVvGRXKgjIZLqyEv/Gw8M+Hmw6Yo5
sReuuRTR1GItrTx0JdUAZfR23lJkF/0XJpV6ZJvz+tTY2tRXLsUeD3Sgu1qpckc3
NtOePBE4zlldiGbJV7eYR5TASlI2Ep3VHi6/ZJIm6WVxDPD0nA1O4n00hEbZTC+N
HJT1W+CGTqUydsfgXJ0ILNmdsnL+ROkNKA5xfEjiMlCudYYJRDs3Tx09QwmkTpCp
FbMLRqwpPrjSyR4/NztkJw3DBJ1/Z8D6EA2ISrpGVeOQUE50s77H4uA4R/bn+1RN
D53i77SeKV4AL31aopSttp/LxNT85uPkyYFnw92JYqQLde52qXmTQd3WRaTbbPGC
LtJemPG1lSPCajdy1XTpAEgj/9kvs4pFgRkdSAPouMEK4YsBW3UuQedCXiuHboOy
0B9hCC7I6RzqlnHntWMgbuVLAz0gyQr5IWY3uCk3GlBkBaM2A2EomHGhUZVqTvsX
Exz8IptT4DnpX2K22i3iiUSm5qUS7w6ZoWQ8MmLMiZK7jf6+RPXOAnhSzWjjgcqn
5NxtGkS5kPqpYAvbKLHVrTZX8QEGagPErAU+83oxhffh7shAM3SfjZR2NmI9LDs/
P7kmW4QWFutDPsa2beeyOANa1/6kikTB7W9yuAyLeuxR32ZdOacE9z/UCFMGP4zn
87Je/d0hOAg6PAt/73NT29FwrBFus0ZQgIkMRQ76kXM9SUq/032IR6j2EdYD49zZ
SA+YgN3z+Lr57p8zpEoFe8sEj3QgqPGMoHzIYxPAlYeDzoP2IyJqhyQNXL9HqOSG
psJ/1yTK9U/itweIomvj3gJcT1lpRdFcrej+yn5zFaT3n2KsQX2wtN1NABcAuoSR
07Qah/0+V8H1BsUuchTRrRwkCMENg99PCR1m2+uAmQN2SKpi9Dqa8E5R+lRQVPIX
WGd7xDc9Le58Sz1gUVP+F8UJjEYGDrfE/yGhuHtcxxrc/nKUewDMPrOAkoXHpSMo
wUIKQiEbQyCIhzJMFm/8JAA3rTB3EaEzmNFu77TB2NpyqDI0lwMw636auLLM5AlJ
lYknXqaytQvESyFgGor5CV+21qaMPDpWTdAOIWkr0THOXBkiZDZiIs2Dz351kVTe
cvf9z3Xb2WAviUGhp7R5UBiRzZcIxK5w6M9uO/Q2X9hNYGZFq3HJ1Lz2dTG02/PS
3noQWI2Rb9+ePsODeLmkXoaVXgNUs555ibqP6zPCJN33JSGWn1NLNApACbSjDP8V
kfOgUI4UKHkwI/yOLNKf2sPG1vnj+nEdmORF04xgLt2V16RrccjAxgs3lZ8ZqYh/
hUdv+H7TmOA0juGrsFIlLH3e8MoVFq3KAjC2R+S29HVjXB+KenLrJiPzuLetWNun
8ib/FfVj7GnpVQdkXDLMPlSyfFVjNQkGzav5IpLii3OqWrtu2pR+o/5lHllmURNC
uSNJObuqgcvwL/g8kNX0BV4EFYNFYdMH38KvigcSMyR+zLSAK+1+WhvVXqvkkAxV
VgKYQaopLAMPRB36SIS6pJoBWN/VvwM2OaER/ppWs8GxpJj4GI44AJzDR7NTZ9PG
DbyvZfbkayMTKx5uOzBk9kvGot7lyVXD2Uo7qzyD8B9jRctJx7slmS8lY6yPkmCj
MmdR9do9u3v9dUZJKDxjFVPKyGbrFb8PJUgpswxFCZuap37pBYljkVAOeadW5bhZ
ZVFA6pxCH3kPI85pl/v1grr3H3+n15Nz5lo2Eer7D7/JfYbDa0Y6CQ1w3m+zqg+H
3bTVmbbJv4O0hA9mdN+o9HQYAyswqT5feYYIpwg919WUe5bQMolm17cDKs4MKZNV
Sp9mpGbb18+Z2Y2nxfo+/TJMsxoK3JKqjWqDOHvMVo3huvCCF0PZx8NnJ8Xy0RgO
snhRc6dzs5iQTXeUpuUFg8LI+cHE4W4zO2r3ms+OV19VAKMgGzJvWT0cRwBcEIko
ooMCkRprCpgD2ZuTEfXA8Mr4ZF+Er0htqU39s7HA/9RjnwdmeSs7EtmnPC72WeLK
PJ7DrnAtRlqS/jyTXtYMfHE74dj58YoK77NRaoVNu9uQaRVQGYQsaT3ZlNmlKQS/
hXW93WlUQZkKhfD3wjPxpDMBC1mbNwY1JSxSZrmAT9qeT1qjkesbM6QW2olz9X+D
2NkxWS5lbBZUxhtxMJKSZyw7nfow6DNMJRcGNnt6N0EE9E2mihlwQfXv+WyV33fQ
vBGDQ/i9owFkv3m8XvIvZN3LOycdjolUWuqfJx3YzNBB8xOS2AUtv+/vS7TdPPl6
rPl+BHGSoHvF53m0vO6U4WWZOolUm70dzAMdrOZKbPZZP8K/Sr7U8La8DPQ4Qvif
WuwE+fCCwq6Y+KjSZPLlIoJBoXz3+SyNgtw8aH6Cjc/QDk/+K7mJmYJXnH1LnlSK
a8s8oM4auNRt8SzzvARe+4VQwe61nUokmXpgJx3rNZBtfyIVXn66IHetvqVeG2Au
ARqigIrCQk4DvSKmieQ+7J0VdlLHaA+a6LWihU4v7PKrLx2Bq/gKHOBcTZsRIZUU
Hdw0qpe3j0xDXsCHVAOej0tpX66wjlCDBeoRWDO4RGMP0GaukBvkZejixsPzjCtR
XcI1TUzeaY67D4PlJXva+ec4IeVDoszgLo11kty9sYBFv7kfxn8190j0nNcye699
CIOI3I80MjWgH+eE5TQExM+k84L0rRKFKNrginM+VgBNOmXwsg/vbAKYtw1phWsj
TGsj+HjZ2xLh0pbaKv3zgK2vDqLgtlWcbpXCrL2Dnaya69c3EKYHFjkNHXoyc5pU
Kyc5V2NCJ0ivpL1cBBBE/kxOadR/Ec+UUIPDRKIt6Ezju5gRnFzkkMTHDOYsnTIq
Z/E3VFFkYnX2Yux7pXOv5tc6DJj7nb/fi6Bix0ORatD01hoppVuZB0r0adFRTU5l
EyK6pD3kiP1vNPbo9Cv8OfEH8tfiV1lkxX4UOLId1jiTJp7+hwt3+zwM8zds66Gq
X3WrNgnxCv//GP2d0C4SuWYauWMZ0wqwW/gKszQo21bycLOpHnoxrcGgFxpbVltA
7l044kFAKjKVDAK5oowuK/25tHuydwTAKMXjTddk2BnG+2T82bDKasLa9iwNDcya
14SpT696BaTBOrf04BQsAhJfB4pQotelr8dypOTuy4+iWASJLVtM6rCV+w3u0dCf
OchSwLTboi2EWnWmX7xtMB9ecZsRb5kE89glXLT1pzjNxhHvtLluxI8Yi+Sj1kS0
KiJe2LfKefs7hMqEMqkk7Y7c0bHGdM/S1vaB75rAHVL4n7Fz/VxEhjly6mtNlHVT
nTuRTQxGUWoGIPS7EMfPRe7AjlM/unPmYr+bLqrC+I/QidsyF01mZDec/m49O0iD
PUI754bzO7QL9yFBNnweu2Gd7bgh6AXECR2Iky5n5aOqocCwRXIMlgXqoR5almJQ
6N1/aoD4rVQf7fi8nVL4uqHg5XNSzZ2SeZE6IEHknAEQK0g0xi44c9EzurCgTh8o
/wWOeZVyCNBcpjSp1jhmU/dvU7uZIMSY1OUqViZmZSeFI8PO6SwlZHWXb/rF7bLT
DrnHzCBazInM5jD58nUsXhLqu0zyPYyZryIm/ycIFhRi69b8dNIMIO/1qvwy4Gm3
1DxwelkI2RKzw7kSAEHUmtlR2oZE3xJ3S8TZjhm0TE/Xjt08m+gJ8ODOwm9pI2EL
9XNUTZCKhadMIgU6aKLEg5ufm4PWHM/IEA7iNsNZQAJ9XRw5hnMs05IeE2lxxjm4
cJeql6P/ZU2ggzLMf3VkQpAUQW/6L/tTPMgOmiO/mbMiur4DpoBdSiKMl2ZFuUTn
B+xwZoWRh8+BSzSqTPWGIMY6CJb5AfsDRpoV+bZSheZYJLIruXv9g4t2ZQf1wRGg
yePJZKD1UFSXzEIKhOv2n3XYN5rYHbc2uPYLQbO1Xantsamp7yc0nA2CcohUyY1z
zgtTEbOpHf2xTaBo9hp8f+EjUd7lduPBVbJXciCPhlO1+J9R8nftcLoidYRYslNn
VUJZF6hdmYKkGftH4CbBfS7KhwwyQm/Su5WNHQHJtCirs538YUXoPPXhddQM2OMN
U9LPm5MNnlqLOHxbIvqw8SR311tEqWrvPp47FaG+1NJv6TSkOY4l9EvsboZHiOUx
Kao/MljgcdlzeGOv0GBKXXuzyrzg07AlT30jcLl8HFbuZX7kSZ/eUVibGYP7huqf
yqHGBISai3SIBc5TXKJMF7Nw+F+LEpjffYMj9YathdJHr4P6oI2/wf9useFpN6t+
7Xfm/68/kON9p/Ln7XqTKrMOhJ/PuNymFi4+gf3N0so2zHSx0PPble5BNvluv+AN
mImuQfWGKkS9idi87B+PlR+Lm7y5CTPWxwnuCUiGrp4AuhZMI/JmfOcxUNDZeDX0
qo+uQl1DpX/pkrct33zZWo1sCNc8ou4VONGgHkYsx2wk1lVIlKdkSFLV3qLQFBDt
GsiJDKwVfHq77rP3b5sTZP6mmyqIHiMx4jaiDIDQU3oLBVDXvhWdGS0tmBfc5tNm
EaCJWc0hHK7+8MiRvotT74z6klmJ55IscDlYG/Lr+2PTSrU7RIFOVJGNRMXN4HU3
9yzQ75D0ycgqXxCSSiEV8YNft7xKa5QSVfuvXq8h+5Qhd6bS9PFpXH3Mr5xdFqEh
Jgxo3qi5tVYeYx5A37DHanfDS314vI/UPxN2GynHdADmPw45jnXJ/30bow2HGJyy
S3TcsGOwxwJP2HNWMTNPPPFCgcr2Ef6A08uKJ6gk5hIz12nCUmMcLpFuDVd+YfP6
58B5QgoVwLboqe/JEvZqvFzYvXF1yVvPtyItAFjQDR1dP+xpOiJZQqP3zvRFNP7c
q2re6n90BKJ7mGP2W1uUfDQ2LQOoFrEY3cxyv5FP9tdkG7aqXIqrubrGLZLCd7tI
tyTrk7WdoFlI7DwE2swAgw3sCYlV6lBAkppVgNXQ4L1iAoBYAQml6lWQUqYyzadK
/GOy8YzmDZgnmOOt8TGdZ4Q7u/R74LoKc40LMPa4MX2l0bXeUJabSHDhYUc0sCm0
5oGUhswsA7FYafmzJUMZ8TnvRQXZbeXrSvEAFi5wO8e01drbFzbUojc75OiWhL0z
vcd69sx2r301fai9z5p+9l7nRuvVXCjduKN0A6l0oLWYb6JUG9AGO1Jqn721rQE6
7ME9t5jJeTQYIPpUpWsPyIHuSGXAZ4jOeZkG+xsIe31P2VUqTI391eWNYqRKCyWz
ISJbNDnWwM57XwgAYsE6LweIDj+uktYgWQijP4RwArdj62QVd3R1lvp/1Y15ns+l
I70lrlUURyq/93hNSzJ6gMz1oqeII1tZNePxtBQzD+rcLPfgqgjQBdc3xggahmaY
I0zGpuMxshvzlevYU19MR1YUalQhGxAIgUGrdZ1dH7JGcz7BjHtC0mwZneFCXQUk
Uf0VBnhqjbEroifLGfhjsb5k97PcR7WPxF0knIEGdV+RWWsbgs/y8cetLioi5tAh
270uqlXANOiOvgZDrYBoL3shcYS6VfB4Ia8By36QuPd424D5N6elGMOVshuZOkU8
lSaQ1r4o/akYlisf2ElETOzFFEHUPgVhMuWqWqkH7N+T0RLZovma9ZGHDJXaiH5Y
tuMeOFY4Z5ESERFpMYHSWpn0zLZKu3YWMuqE1Vh8fsM+/bxVkiAe8WFyId/PJOZG
PK93+EVr1mbVn5VJ2XLXarPB8MTXrWMPCPJg+geqLOYa58g51J13xtc1nvHTBsrN
MTuxNV/ZLZc3FLuKkdE1X9FAz7HrLe4c2+Hc+DO/RbcE/9O6s0ag8UpGbkXRo562
cqABGaiEwS/iRdCCp9Ezp4zAlCs6Z5b9XbNxc58QS7WsN0FHfax/otb5iydDUSDH
NTOZP6nqbZlajX/GDD7AWfbYfuwgHy92ntTTmCoZ1iNtU5C5LzhMRw2xHkFRaIE7
R8+AfviBub2eH68B71/4Y2Epbq03aFSqvLmb5ub4CEnKKqgR9QiEvthIkq+BcvwQ
VIN5K5xsVSdhkHI2zp3k2jDu5i3GiZGKn8ZRWvGkbE/UruWHxwuooHiGzWLBLClr
kMF4Hj0yoM117AKZZjvTp6fkpOJyMZ+VDZarB4ov2JsS3+EqNVQWxqtZiGPA8YU0
+82XQWAe+ZpVx2ycz6aaRKxZQqq0VPFbseHBOTOxDNHrsFyiiSsiec5ETr5WZN5N
fq0KCL8TJWW0HpMT5ULnGH7e1C1ogqSifeajdFXu+zeUtdIjEX2hPiyaK6G6MEqs
G8k/tXzNJ072eNlb8s6rTh2BtgOZERlTJPC2pnqJt6KgggxrFURcjSfh3NogHxtC
kqmepYxlSHfrY6EHbCj73gfTp+P5y4GQFroHycdfLEDtZSgnVC3HJJiV/2g4sGoM
pDMIU+aIfDJGyR5IRpPcAwjDErbp8QywnhWwOfI053KCIn0kKNA4mSnVeofpimmV
KoTenEYu+iCbsSAxMXf5BpLhUNXEOg7VRsMSXCl09t5Nzrl9vQDgTwmSTG9ZQZi8
F8c7CPxJfk4TjpceJq7IOTIzc+QTHXLy628wYMG6Ts4r7l6Buj3YxFwdB4SguTdP
/hJPYtnS/+gralH31YXF7AC+RqHgIVSGu1kEYA8CwBENlOL6BD3o71wwpS+eUlq8
NdTWbB/3XXBg5yHbQIbEBU2LxQJJAErWGG6Ln+Tn3gfOSQu99DBw8+Q8EMUHsJ3l
nwQW9VSyRJ8zo0opkgnMZHFtLbrDNZEWSewNV7SlxUzSgFS9HErLa8Yc9vt5jwbU
aoGPzbCWPDHYfWlejgJT9GgsLHXRbmYB1NkOOA3YpiTkIFGRvJhFmlleuSw+Tt7m
HjlSmD5PrvICwLdLt1CvUFIlZq1x7T7EsiCgcyhzRZit8ze+MykhElG4a3X4EvWl
GeRqOGMKBCOuy78oCyhYLncD/WXkifqVP/AbA42NheO6fhBy7FKcidJfY/krPDZR
tATpLoA4fIp1BCbBHuCgQIsZo4Td+XTmanpUQU1LQMEB+ZSs1C1+TVtIHA3nL6FR
WCoT7RUlTR5R21CeSQFtZLGMoVzgHAcVv8y4udWDBxWdhXaOxM+P0Ny5lSeK/cCM
fbaPYGSTo5xdm9n8MF0bHTwVVY/lTat40LC3IDoAnLS4mN8P3HnJRqybqSs6E3Ti
S6umBavHsoCjT7PF+jqghHJz72Fyz5Vvxaqrs300AEvnqyN00oD7T5FPjapt0TMg
qJkElS6ip51WMgSIeYToiD/OhYwIEeo2+vQeWr1BEGkB2Lj30GuFcBqowvYGGeFp
TzzerC29tmHhahxj9/d1Jjv0OQJATdKom5CLjCbBFak27MYArZ8NumO/MvyATSKS
2TqpqnzzMe4MAjZk6pTEGtzwh4OU+i2ejGT0Q9BuyPcyhlqhCyT4A9vTuj3BadDX
lHkrF0i9cweYthmW2xhI9u631MqKfyk1qMImcuC39+wWJP2QS2sp5cK5WNGSD6ML
Yd7xsokA9RlHQfLZzVWfyVDiiETMnnba96AAKQ5c/W765StdWZgXM9IUP3R1poOZ
ckx9e6h0JrvfiI3+4pGxnxQ62j6isvK86ivKjjc31SecclLk/B0KZvHKuxBZtbZQ
wzsE+zocgcwrgArJoGWO9lA6yh0ZHjhFQ1lxr2QmCs/xxGXnLdRNQlOatBvS4lxb
m2qK7BU8gJRw0eAnJKTBzObc6VGpF/JaiPjT6DqAIc3vPVCQwc60KNuGe43Xoc+G
lquaHWXzf49S4wZjFqcjYJMoR0qUPoe/boWbBdVFcOJtv4rRZ2Rdcu06RoVj/Prl
9CqL6rPJf9iBfCdOKGbfojB3R9ilzQKSnLDGgZh0x2Ai9nv/mEfqDkIbnXVgunfL
9DOllOK1C170knfi3l9uxIMuzINDULYWRn5PY+E+1KgxbKN4JZNLHzM5O+3/TIn7
xzeH9Z3J1kOVwVEK8F2zpyN7X3TuDtywaMPoPfrgpUUVsGKhiyzAIRsxCmFgM1Z2
6q03IgKZlTz2LHIbSWIBbM6qBQKzBYcsvlVHXq4ldqH5L2AfqeyCjB2BRU4yqXfo
hWU8TgcwxVzE2I/bycb+MQjoEDfden9KHJxL0RDfZTSFdgurI78dM1pSFD3vVvQL
BToyH5prN0reumjy+xOlJsYb5UnTU3lFxJ6iSqMwoERWEH/zKIWmKnc4kjWjkydp
T2o/VVixyxOsvXj9ZmtrWx+cbLGSJz3hNT92roNAPtbRBgBhVdIVTPoIlNtxIpxU
aKzaF6Rdy6vZCYOXo6ba5bd88FscI4hVX73FWBcMkUp26oK0VLJMOp+L8x+RT45t
JlDNaIlzo6qPENznSptSLZdcTsQoBYd20pTOseFFm21HAUGwURrIt1uDCKXm1uAT
9exM6xOdwrWAPJNc2+Qdg7UqzXVtBFYzxTyYhjeDGA2oHXiHxCsRJpDR6PBfG4UB
SbX2FcBMMfJcE/VH7MwgZtNRxqFh/AS4KdVUQR40XJsORGvgAXQbgCngMGp2NVOD
pF2UBSGCIyaRTYdeSaEzmuKsM97VnHYDBaPIZ8Iv6EdgNClDpizH3B9szr2rpKUf
AzSI9yHEQZv7FUcj2l7blqqAOV5RIdeG9wUJjmciR5iYDlpQBaoyn/3WQ4PYA/sW
VCqsqtlnUUZYifvDhGCbBurHiJmKhjDsRTUh1+w3abodN840t6Tkuq24JsJSp0u3
2tMtN1/ZQP+GF0ed+dcCa47WMtvo6AeusTRn2M8uFLsB1/ihN88TA+qAacs0pZcK
pQ0HeTjqLNcSoLx3tA9fCQUYJMr6vWsfLQ7ttPJNdBwB3B3RuZhssyjY4oBJ87zH
IHBMibhaJ2qY3UWxu3MHdk46t1BTQ83Nj5kiS4O1hUe2ejplZFF3nmitOJG85k56
a72qBISbo8tIhTTJu0QjyHhDWQ+EDUoazTGJ0A+dFJuupUVby/kV1vAFxfkjdPnc
2YTEXs4jYf5kXnt1WNjzGZRPvmwQBVc59PrkD7XAxTwHdnfPrcGtN3mXKSgaPc3V
eNoqOEeIiTIQEgChPWy7bGJV0T0yQvIcH3YZ7LfVIVU3yxYJ6EYVtcgEYZflaYo1
Fjrod/Cb47UF1q15VzC00FWHhz1MAkVxh37ibe2Pqgw6AVEmPo5oqT6Jh1B8MHKu
WE7nNerJFuLWun96IxRY2spolbXXrJAlDNfimP1eeK6vLFVA8DBSXWqp40ufaIE1
fsmvXcZ/u1zQqPNU2025kseK1+OLl53sEViCjqV2d2J+xsygKkITYk6+8Qqt9Keo
vl+AqI2bU3+OGb31lgF/5gT1CM9R3jgqZyuuZArGhp6Jtf+I9FNTkCaWTJ50MTjk
vgeaBLy931wLC+XZEpG0gshKAe2UrVEPH0UvNRMNUr/yoS8EhNpedzhr29s7EKrk
CTKIjWb8ysrDbatSl+F3UdLRW4J5u+jItMmB+UMIlCzkkhKZgdHEitCqN9qY0D+c
TmhjCuOL4zeLsBBlBxS8qvup3/xAloQ7kFo6c3oGLFfMl2lLeb+G+OhAkv2W63Hs
kRJ8WA8HDSF3mNxG8dSZcpoGi4TEqeaoVnz2icFA6KrBGr2FNV35KVscU+R+Bqcj
/UdaOUIPG8iL8sqEs6+tEpzeQJah21/pCzuIToE4bW3eVk0hgc38N79GAzgb+zY1
DltK5Xei2PgcFeJxCNtXsHov61S1cwo5b/g0puZ10MEGZQpuRkuJQeTTyfwDngGr
Unx4mt/lCKDmns67CuRN9/r4yYj2ipxDajmhnMbZGRduRAqLakHJ2qiXxj4vkCqD
DWHsjtZnFJjCizDVs2fSUjYNUjPGZpvhgO+4vLequcjVVMQC9RqUe0peY6eUffgE
XgazUghClx/EHw/T6LYGhcMiuilg64kEK8+7BoBIWMPCgiS8ZGHU/kteIihT311x
DybROONoO09W1/qWttm8dHQZi0saeJ2uvMKcqXF/G2aITOUt8mHyxoplkvj/+Dmu
k0W5YdF9HTR2h0SONAB7EP7rs+9v9WdetYQY7TGiRQcD09D3dAlDPcPU6Z3lXu7/
0+/GQDjBPbcGksRk+JoNTh4LDNSMguCx42tKIahX+oazdURS/hBdjK0i3o+z23Ej
AIdt4s4VsIup5UmdFrw07P9DWhZDqII+krZsX9RbpPHMRL4nz4+PJS0gAAxnlOpG
NKeMn5qrNmyKxyb2yoPSsjSSNlciyeXIs18zqX8BFnjZIG1u7aj1ToX5jyR9iJ60
R2QNXxnP/s0jkktlZ9BQpJ9mWVlF9RISiqjUGKNu4LidrV6LqWelsR0xjfGE1/74
wzZRSmWZwWuPjUbAY38XF7GxlJmwwaAncj4tlUmzk2NEWkMUR5sIx3gWR6jNaDuM
YK0qqBYPgSBJzEh15nxHIaACxdCbuac/PrSaknZuSDlbEji9Tbap1IpDbuWQeDCJ
3XzsTzn9kggfxvYqTe9Yr86hnmh00ZuV3quB2onn330ff+WTS7THcKu45Wj/cb+G
mdJV3E0FD96tn8HSZvAh61VEJOYR/mtTcYygmeUWIpzb6orgSw2m55XUOT6oh1Gq
BucXuf7njd9PF24HP/QrXI96Y+3yx1/Suc0xHny6ohHxsqIgHA5YznO3oS7x858B
HCGxbW6jPK0sR8MXxdKZVXPUsCEu+/20lOmL+yitoYVLf4whDKRmbh5sL92SLgpi
A8jPcixM0Zq14fYcBYzE3etJ3dfZ1qWDr9Uw60rNBVjLZhSINE1swRK6Bdh9rbGR
L+OPI8c5HZ00C5Vbf94r3UuPZorVFi/NBLCTPtgagU42ENTbvtB+//SddRSZMPr2
68Rw+Gl8cBrfDcTjYjYKSFQuWGSpotIQm39EIqcVsslksNKn6c3gUToWcIvQrSgk
nGxOBFeB7C4E1iSEu4RqQmrf9XPnlITaqEB74hAcTEMhTcJPXzdVeS6bYwA7GyqX
C49/BM9aAMe49SxSo5b3buW8eCh3h71U+16mQI0o6DnxcWUh1L+lkAXPC/tQCLGk
+i4/suTmnIdCxCaLq4e0lMOSZSXXz7GDoHcbeODvH0eB66QmW+9DX/0Iss8cdD4N
4hMtCJghKX1gJXXRRmSzOdgUL4ACP1Cx620aORJEDms9seL8t2Fkk4oBKbWkKoLI
gKf1cLoVRJ8LT2uYrUlfpWeZIDjEefOgDnZx805/1lYGJAMgfEr0Lqug+wNoh00q
e3K+eT67JeArAvBXyRxIFfedPjhJO0qffkJ4hZBkfP3a412TeIYDkog7gQCDVyI/
du3C89FoGWj/es/6gbo0BLHWW4QHWVUAMlM2e+3OabNnvBEOh+pFyvrCW+RqnCyc
GqsKoN22yyAC5yYHgh+MFXtWtSkhroJ71nRnNZ79mQwqeE0gvLDDUS/sACeHJnwp
GkwWClUNQI4UKUlD6BeoQDmwkh+Ugpl5stp1qVKX43qTfCGuGUS3qUvKpfc1u9zt
q1vD4PCod+xqlB1jfAuadXAzejSM/u1aaWmrjNkUsiBcPzLGQfkPDuqx0zCJmcGx
zdbWm9Wg2NxSGD23XBJGSpJqwwyNlm4ioOGa5aMskbV5XIIXXltDd2stLMNKiuyZ
XtLJ1rQyItv5rid7ZgFVgRjbzorMSXP6HsgyoYYWz5uhuEEJnlkcTgPXdwey/DwX
FKvMBlQchhbEjM1mum4/ZbeIRKckA9QT1msfM8se22675eaCxG68JfQcPuoCqHMq
BGoafnreGshXa+cHeSxoUMXI7aGLmf1IPAlKPVjHCH5uvUyva38kmRbsul55nv6a
tJSqFG2xMjwpVE/vB6VGHUfSG+oQedTZOAWoMCVGUEQT7cAZPgjC4qf8OVxuS9Hy
Tyu+wM+b1TU0Dmhponpeq//HUMn96ziOIgKyJ/sYsuQodzEwJOIaSVvqdNdtvjkj
TcClOZJH59DAAQCf7nVOUc8rOsgwOKtH8Ry8e5+W7Dr1xlT9esHeQAzExy97dAvJ
emku0r3zFADdkOFMT3IxvMyVrJ3Yf+TIUo/M6BoRWVC5Aau/C3Dhh6wOvHxgxwmj
ueqjqBNfQHHRjYVWw6mzqrZhgmUY7SYZLt1TZHqYOikpcXVTMftu5u1YLK8lYRBw
OxlXObZmjBI+Fz0GUzSJsYMM94T0n7+iOnTAf0EvXzQsbw4AO6uBxTJ8XW4qShFu
E8ZNFr6KWvrnQVgWEP6v9B88Qej3v8vD66BtQSxcDk+A2vRg4XMm6oKk9oFiP+Tx
/neQf3YTst36hoFqNg6FF+SrIeuyL8LJOicD6foJfeIX7s2TtwgHnUuJSWIoQZI5
/bgctE4eZrcEusUCLKzQwC1Bljru9tgiTKvW428FaFi+XKXpvFCzqMFzU3rBTcwp
jTvSeWfrX0awy1RN7QPAOIIo7IRxZoL0m6DOAHvFNGGG8Y4tD6oVkK6aLZoB62G5
SvflWc29dIToUPbgsrDxYVI0dv1vY/1usYJBIkuFIt2bn+PqFQXOHqKIxYrAruTm
plgC31ZlItaGxEk4G7Tt5BR3+0pAcHA15gXCjbRBtrBNxf3YmMQVDftQHwov+Q1v
+1N5KD53nocNXw73BvmRqJ0VbSkkugxoercO7EGi0gTaPdDBaeY/B+MxNOnfVOq8
uUxCx9dqXKqn61qGCOC+scbO48eVNkJE/P++21/1bUCUNTuC5OC6RdNX6P/LlipL
gECx4NUFarPfBFGf0vKgg489D2dtvRL4O4pXg5KnAxWZf2VIwxJEVVf/udIMux1A
EfwxjO66+nWgNzLmTGaLwu2NwwM7r5tNJgAzrnk+YrGDvPdezvmDCKq/jrn/0mMZ
KyMjxG2Toyf8q7GsB9oPRGJMLCQRQ/hWg0lwsWkqfFBBu8eG0cNeh7t2dpw95noB
tUPnIYdmk1Wl2r1rY8+Dr+kPRsqhhRsQ800mXMiCwgtEfxQIuDkDHuca7/i9vw3o
WiJKStL7TT+ICip/jwPpgQ+YZpH07YCfZqd4tU41tbaZ8T++1qyE/BrG7vyRFb9q
MRQ/MeXBR1px2rhq8RD8J5o8avuaRB2NHinybsJKZNCOT4ZrqhCC7emYTOJHzmju
o0bYx4lRinWiq1z+GViyrwJC9kKo62USPvuak89DEhI28Ste/q/sm1RkXrqnNiA2
3AbRJY2prI41ABlzliPLS8RoaXZTvBP0de+/9bKzn9KHo2C7sE89acRs+b6Ovoa3
m4CRXQ6bqWD1x0hRP4ofSfyISkebNk3HS8xDEn6wpjhzn+hjoDQtlXzjkZU+aHTH
ID7KCsfpplKKLJSSpbjiU9q1Ots1eGpKzGK54oY2V/Q/Kel2vGR89KJFTYGDG+hC
WZP4MEZ9emEXBIvluo6tDAOx9EYz0k3Fd2EraOL6w9KlHcT13gjQ6nXATL9kuvA1
GJ3drxIb1NL3ivJpXbteCC2gRMxtFtTkI5PYFkzt4mwm9KecvlTtvFvr10qonPx/
VwIC/jKbifohgtpzt3U0aawNBrCY5k/r7/yMBn8HBXzGc0RYQ3riJ/bbjm51lyAh
zu0V9DJQBu6K1N4hD/VYLf6rp2Yu5NMjs1qBBTme444wPwkNmMzX27Ap/AGzQ9BB
CY+lQG2wV2qGN13gGk6m6ee8o4/+WBX+oZytPgt6NGIOr5VKnuXwGf4a8ntHNh0S
4zyETJGvSDZqN7X/vuBfiXuaqFqCr5ACLGE+K8dpmPQVJAcrDM/NSHgZ2xGAGkJz
TS1jB+KWVWicDz1ywyBV/du3ExBYHhkQCDuLE1nFGdcBLmQ4bBBzd/QbyP/5Xw1M
xhIrnKK7n4dayRZy883NDTvfdUDtVFiTXV7We6DLEtAFv/xLrf0gQJwxxgSmNPIA
88G097/KlximtMBzJqjh355GLixrZJQSDhnj4x0IsW7+dwH4xTJefK+mUq8VvK9X
tXIV2UvuCfFQL2B+7+g3P44Jf7XBdZlCjfLA4atqXRJjkFFhd0AH85OB0M2mLen0
B1gPyKgJIT/ZD+1I79Llxb1JBTWRLFJY6IpXUt4Ev4g2Rwx7+hTt+4fp69m26hVC
0jGQZyZjlx3LCe+rlWm62Yh0RVOjfwYRRGCMih3HecLPUJEWQA2mrUkZcXYUA/Bh
jaRRYzGvMculYDWx+EjegEZWJEZ3jJc/3WaEgkDE49SYH1O8rKW+YzeHUrHTx8N2
OjNRroIqJJmAKD4E3S79C4ToV07sg3RcHiQpI0HnP9AXFj+FzLh8/4NB5WxFKX2Z
JfqYX2xb42Q9eF/t2DxfgNIsZJ0HZc8OoY7mZsIsNKOBWJ1anvQH/xgv9AUKsocm
vSOZgKujKroOORzz2QCWxkBGdsAOJdxCmAw8vfZGyU6vkaqIdqhBSCY1754cdIkM
rvkI5JkUZJGfIVADF6Z6w6CHpFd1GaGU6XXqW7fkwVCCERnIbX5p6T6O2tlpGAj1
e4Tl1Fu7z+6WAdWal8SL41/9beSXEjaCAUo5IcefF/qYLyjGZwWUcIqPaq2v18iZ
reEeLtLUbYTsdR+0UqOuiosNYLPxIukxjo44gzwPPUgECLNEwZpXZmm2mZHokGZp
+r4Y5K1ps1zKz+g2XSKHmhVT64fPz8ao/WsCtl3cvBo4FMFqO9E6mNFZP2+1a1GJ
lbtfYxfkEoyiI9yVKye086QgdA8VCHmdl1+N5IO/ucZSzpjzwEQWGFKfYE/ZP3vq
8z1h/7MoNSbDXKeKlL/YZ4QPgiDFFYLen2zS2Cr2/9JU95BXQ9ory2Emwh75R7DE
AIziEnQR11sBV0fNq83xPRixDPGXpNLihEVhE8qMIqcTxNtzFrCC5DedXAR2TetY
pR6RHfIvWubgBe0EnvU0KzvwVCet/LXTzjYYq1cPiWbnFSYEneihpEdJwnrKDo+j
AIHVkBigGskFqfb9YvFXU3kdWf1HkE/GFyGmhnVRZP4z8tM1em7CQ+cQHZrXJZZd
Md6fl3vll0//ZBYElBgxiB9+wOLLWUPbhD/zYv7eHGcLr8XUc1BtSlazz2pTTGbB
QVAf5jZZHO6Kx+DtAkIwM3nuL60BWOMERC5WmsG3szoVkHLIrKROBn9vuFWZfV2S
4U8vZ4IP8h2eaEfJd8IOl1ygolTI6/Hzqva7s2VX7MecsAGx6GvrJHpp/h8z0jD9
bS+NmkN6MIXbtUsBHChnsVfFH1Y0cihaZPPQanaumzLNexhcq1euGKPy6tNpfcuj
4POeiKJIu484XRl6iRPN0+S1VojwP/h5UtpdVTMYrVX7TTTV/Iyz1sIm8iRBLefI
bkIAZagv/WqeL48qZtNr/TuzmSs4qZvEiGO0l21F6AqjAhn9gBXFPEabe3LNgWcJ
MIAD2l19IFFmrfK2x0yLS2MDa3A8mkOvBfAT91RXJ8b2NYyOXnRD32HW74OAmXsM
Galn3qhi2tCbZ2KLSq5144E9fADVVgzFyAcJ4NK7f2D8GxThE0mJzH8dC2lTH+Dg
Y3DgWh76ybJK2Ig0VED52jsEMUfLHYjvIjd54+9oVVsob/IIjdqjgcm6KJpRTl/+
pvgvnK7ML9lTyxNBjAzv3aT76dvYh13lEXwQpqZ7HJf2pYtBPINZsGhsDRQ2zNNo
nf1L32nsR4m10vQf2X2vOgxAQeZwjj1rM+BpnrHxLKEhutxIikSZxK/CYz3s4jF3
OONIMq0Bgegn1UVHN6ondzfnxvksg9YTzNRC2xHTiTREd9bskj4aYWhN+BRzBsBm
KHLFaR6Ib8kzw9VMlmiVKvbJ4TE0OGtiU7CtSk4iUI2ogtW0vsI3Ni0t2jXYau1i
WLD+ecgRP+6LlYX+S+0wxddTCCUjFR5msA2nYcbHVk+s1xo0W5YjUe6egvpIv6im
V0Ka05mUm1H4Qs9Oj2C6iNNp0h8O3bWW59d/aYyoYhbpOTMsxOJbB98UAhHsYYfp
GhaCH/KNkzxGh0Aic0iJfTw5VVhNAOMvF1GkW+K4Wt7zZhpuVihg00cWjPX6A+ac
/uZx9ap6IMgnGBGw25LhvVhMVtNk2RuD2esYns9CNRGMgj2w+Rhka+MvfIvgTSdg
0oXcA88sxTsE8Kb7/PHKWdtHSX51DM9buttYek5lJPFNpzUqWei2hJhJNtjD0s7Q
SUOs6fcHgDv3aeCMsEqp+6IoPDxD5Xz3VRVAZyQeMooaegTS7N7489xcEm7gN+TL
z4AH9EiLLNWvmG1SknNNRhZ1tCZNza+qcXGmULHDPaU4NasIAvNo1Wwqy48JIVOp
whgloJscdkPQJ35/4Mpk6TRuEPjPCG9dMP5/u0F/WbNxVstMxv7R7PdE8l4ozx4g
NQpdkTKbAbwVPkb4NoHGPthl/xozPvclq1pr7Myllvhc5h/xZlI8RihMBagZ+UEe
1f/fUJVYZUyM/qfjx0k0qAV9XSJ+ASHGoWhc6ukqBe7jlRSi5Uf43X8k35MNadH4
drajdi5XXV3HwZ5Do4vtJzIrHpCFtN5o3NuCyrFdp6Gop9m5dRsDlvyL8mMjgIFP
jCuqbWFBMVMjmI8byaVpKDkf14wpr4kac92/cc6NJQSTnZ70a0GqA//mv8f7oVQ6
/RE8eUfSLfnSEbw5Hpv+RlwXT+8kQ7dFWA4cavOizD4L10w6yMcyE/wzjoKYw9C7
5YsQ9ZWZ/p2pUvdSN11akPB9uG7fT7V5uVizUGOS4kz7/KnczLtbEfSwronvF0hw
ctJ9ldm77lbcM4NHdwFgcsCipEhQC2nds1bAkGumHBgoQazrXsIkNUs+EgnkVvJQ
G1JfQPi8Qo4drLsM9g81JoOnAdYcgpSD6fZIp91T1nN2sbPYjJ2SEZDNbjDd1pYY
Pm+ziDVEr/c7JBDCwU5bWEbvmnN7oMxUjVXjQFJxxGxrh9jkuCAAJOsc3WFx2uxG
ugB9LZPGqqGHSvtOvUEDC4r5aAuiT38mVL2h/yKvo/Uymz9kaMbY3WAXPT5bvyy3
+KTxiIr8vZAshfxR/zklap0xd9wPlNxACC/L5xXvQtiFbB3zYFgOVyVdMnjaU41h
Q80qQy99pmU+vBXr1CXKHYxfPnioNuWjnExijl9k/CRTWvivQe04IHFFHjjQ+h5a
CvqrVlRvf6SJ+4SAH5IT4+NuNMVuui6i26FoqlHi+6ZCONcew9nx7GqXs4M/EQDd
rwhAvx36J4kkSDlfViFDjRXg9QhJbjPq7hXYUl9QwmzzW8BZdrTaHpaJox2S0T+K
OU3cdaq4ibcx2I6w0arzqV5ny2i/CwukxS8Cs/X8A0rvOOe7OWzMCU5aNS4l6LoM
RtBJsfAk3YNKbAt3MfmbQVM1Mb9fABkzjbVU7qubddSWDtpByn8san+DkRG07gxf
DBP/RtqD7/TMwPjD8lduMg3QOFqAJ/7YPYNnNnLqy5hNZQ6ISwpu/RyiTZQGY+OK
vsGxowuN4SGejrbnyh+3jaWJmK/m5S+tnKo//GBXGEI+XK4nWQlU4cVv7ILJVN1H
p/MxD2SkdqnIdd34N4gzwDZDU70UKZDaW0jVbybI8KWnSmYh69AF/vpMk4TeqyCP
g4OClNCZg4zsr21M0oMPe2U2EgA14Z+3dYC2+5YHOtwElW5AfN93gbFONP/m8OFU
Vm/bjLaniy2q4KcnRLAEKw3Mf8T2bacbjGK334Dmo4sdRsYxFYk2+UCsovf43fna
aLXpIqaGK81r42NIlj/FwhUlMx+NZ1Zu70FjzSAUGd5RTLyZn+46W/GdsD+w88me
+rjetxYH9wu/ZKxge1zRwOTReQ8G/XJoR5o/WYNI19Myv6Z+n9BMIo7ZRojPnwMd
Hp5OkAXMabDvR4i3qdywpMUMKc56MA9/oBT2xIxCETVTyld8FNwbSfKGrkXWAoTc
rsMmzV3Ph13pNaxFD5qjU2TWZTxz4MTtIZRK8WP5w8bpd2uk0AqFzlzNzqd++tmh
VOz5XdDQtKLZHT7XndxdG26vjJgud8aM1W8fB2KiJ22eJz3mf7Nb3RFDCUSBNn8g
W6PPrPr0RPksjrXSGWj+rIIPeV+Z4flULsnE/lrlBfjkzp3Za4mLO7tSn8LvHpJb
jKhxo1hN7BoFiLuTuCi3wuiLPVk3lg+apmA8rKllFQAw6QN5eHkNy//UG3yXnkPq
H+CyL1VJeaSyheK819n9Sn0H4i/www3lHPb7sCQZCDhpJQuRwvbu74QoAWkUNZqS
UTmOcugRtD9ZnVciRw5cgBvnk9zTGsFsD/7Dt+zbwjWcc1uHSJKpgTEgClcsHntc
zZAzjqjZUqdI+jiYNr6b1+ptq9VPTvFYT0m13xdV1vEcHYgSpMPavjBWOAqMuo9D
a3GEPlikSvWdGMBz5zwxRavyLaUWozXR3p5Ze+W72JfhL0GZNJqhIJCEEMleIwvr
NRwqBReVOYD1StF43atzMN2OH2mTa0h2YZeGj+9hTPtR63XLWeBvohDeLrD/z99f
/3TM6ygQDXLwXgYjr/y6QpPaN8iDNsvCjJ02Nm4vQRy+ZYO6RJ+W2fu9xscUQXAV
sxi+xhFuOg4D7rrTJtFDk8s1xkIVRzuRi+iaLr+9TZxm4NEHVdDiHyS4bvhNfr0d
muO5BWsnGZQc63Sg/ygioaPF9sPS2DYb+3ONlSTewbRYqu41kXZ4p3MOgGoatg4B
Qn7kqbWBS43szhjfrFlSJkeeJN03v0DXvZxGUdtQFrAUIlewQEchDTB89PZtaHI2
W0vnnLpwcGoBa02sOgk8UzzleycTFnMaNzNwwYOLMuOUHzo0MjbVOAMwcNdQ97Fz
CWx3aekiDm9y2xaG1SHZ8BbdAxe+U780Nna1DnLQ7VSzHcuYLiE0gvKXWXyBwCZP
6EPGCE4SP6cGFkyv3XriPY5UE1URilIGj5QGRNvySmKIKUoFHIUcFoAYWWAVajZI
ECkHQ+K64H2sADUfetCl9hKQ8A4+ty9zHyii6K6MkLpysaVzW4Zp+6zIH+D+5p42
HpUlf7/SBfV5+jP+lzTxlJugOh6fdEENsoSFCBZgzlLvFqSBfKuWWWge9PSoDJkC
cvnouRJvsd9IkjbXMtIJ8/+9CUzOnXCTB1/RHHTV0ZOUMw/pEaDFhzHWVVk+23bK
9I+jWxqTwURiIgO+hmmbz9iuJERJ64impkZ158xMmIunhaWNxda7C9VAq7km7xjL
P76zy2MN0t2dwQTNgJouFlPndly5sCkNIPl9dFevVKPVyFsieVYUwXjnd3kZ4DLY
ZxugY07aac4nTl9+dw+3vw19ySYldZiXGv+qxbEMGd370BsZeZBXcKM11ooilCC8
W8t4DPPoASfnyitdCqNbecEQNMiRg3TDRBbZVAjjwXbMJCHPtLaHE1bnF6/XZkfl
ZyWiuYqapweTicwsHpHw3cg22ehyk5stMoJ14YqoFA4X7xHCY3HRBmaZz6aM9SyQ
NLIQb3+Cjrkl4Mfd92tT1z9pEF/oHflv1Kfp/ItazRVq3xs4I1lllwTnQ8NN8UcH
yZTg38ZGPIFUNCR2yQTBIy8SrYdiVDQ3TVGQqW2ZKLcWnSSCuckKCLlnAs6jGntJ
1qqZsgQgUSFK1Vc9P3xSbuQvm+hTRFFayOHX9mfxv6iaa5shA1vEZW4MDDvOCiI9
wZ8yp5dLinSx1vIg+rrvfOw0D/9UyZegKRXWw6OAOP8+rlwwAruX+as6Ycf5FO6V
iIQCWygPebqfo28QRiLqDCdX/BlShkpxf9kL/PDcYcdx040rw/03pD9OUxugwrl/
W/5hX/CJjQYmTC1cQtwX1Vkl4u7ellrD89iKXl7F4X8IbwyfwVHMuX+jrIbvd80t
DGa1OrBQzakKWoOQ9PpD+dq7pKTPTjrBUvKvN239pl/4H5HjDAFwwA/dW3XUwhjA
SbhGE4TRb487QSlPyZMiJuYg5jQivi+XXTAQucdoiI+ga20qHBQQMJjmXVpjR3MW
J55l3kJGTfZRolmZ2TSFGf79JF05lLWBYJO8TVuWly0wrNk7mmbtDyqmFlpzcddD
6YDwMdYl+tGhDJ6BsKrpHid+Y3TtMGmxIiMtGa5HKj8WVeiv1VSRyYMdCTTtpJr7
WS+graAE4uS3RJb9NvtPt3+7oUGlwRldSVKohA4y6kBYCLOGHeLS9qkJR4MoskUn
0jfNzSIqzcD7d3uhyplQIcSEIKsldFsN6E0soIVd+NyAkWJSEoo3pBRNZ7JaLqNC
Ds5UwMRf7S2fiY2o39Dfkkj0JZ3m6/T7xktr8ZGqREgXU5HOPraH1cXmUKBmWdt+
MniTDL+zHWa4G1dWPbsJp/I3aqXy7cG0ChbbsDSAK7hd4+iB1Vin+CfSLoQJJ8J2
2rmuZrTZJFxwMCd6yewwJBCyRDK5Ln4QgCo+DqPfwUMY+12ZecQr5Bhwk/ARFHUW
r3EVvwGGk66aYfbfdD3i78Qr5xegMgrIp0T7/a+ORioo5ekQY9abYMKM3jXRhNl5
iel+ov17kj4SFxhajjHShtIijVmCDfc2IfcPrk8RPlgQ9MpVYcYupgekuYLbn4zV
0ONRYKQpIMkxflERmbYB+e9ujPsDmpxdI3/U9XBxqBwZU0XQpHLcvhHytKk6CTsH
sDtQN/6O7PUXjywfLoMCv+HrP5eGe3pqdeoUoAoNEIoXGwnFYVSwQL6hb5pVkfK/
m1bRkxTyKKdESRELprD6o0TzVrZrm0XZhFB1xSgbzqUZSrcjXA/B6aNEOe7z1UYb
P+WtUNg/UBqUcl9UTf4XJ/J8dXFhikk7MtxN0zPfguo6dStBWO+hwery2ZP0CH5P
KYqYcooI92MKPkqA7/ONXMmJVQjLYKQunDZOlYMDany5U2Ng+1Hti9V2rpCFMiPg
bscFXcCzoZ47HxNEu+OCkzUWmMjFiMPX/cnaYyWw5jr8Ijd20Yn9qrXFnZdzsmDI
iIcTwwC6v9Hq+43YbNCnygvwDMyg8WIFa8xFsfS0shfyaglmi1g61vv00TW/iid8
r06NqlgkpBAjfUR00DAXUdKrBMqzo9SeWkFXnCV/F7uIVMT4iKGG6puXkAwqUYgd
9YYbcGsz19Tkg+4bjCAa/jM74toQsC9nDVfiOEsxwDOLbTDPtSnhBcK1HIzcM5qb
+PXTWtbI4Kc7AH32q3Juk9cQN4tXVvK2+dZWt5u1Gz536E1BADfoxngAZ/X3r7Em
GwAnRXppu88XoZ6DLGWs3wmCC+ddTRuUeTcZ9F1NCNQc5/PomCwBVxeQFgtV4PLe
qQm8HnGXDznzqpQQvpkn4YYICWNmGfNBNEM3gBxwZlNMWFz6gA4+2BfOtWnAKkIg
xyMZuXe3Yp9FQrH1XeJ4AYgmApJI+6S17zfaahX6/RRywnBQ8H2cPmJQvwIChD1E
lr/fjM91cbrbpCfDR450dx4haXtZqx+PxmVXRioTSVf44KvMUNjLLk9HDAYr1XHP
+B9RpqALZ6n/R6voUh3D6mHTqsCz+jrI/1qLL06InQRxH7wZUh6pzAyMhGfKxmld
p+NJ52OfDU1Ik2fCOjm5sxTw7xXdJUPdTbHH2CKKmgYCMn7a/IJ11CCuwnitHWzh
yoQ3hw6hsSZOPxvP1Il6ad3gY32ghEo5CJd41Xda66He8Cx/1UWBa7wOB3jx+Jhy
U/I/im18flH0S8hIO5Y+V9C7SAwHJck6Qu03stozK5kXcmI9K7Y+ftQI6PE7IXX5
FE53kqbdOrH3aZeiaMn/mmaL2CdEOcceVQFY2VVJwm5OfXM+m11T7m+gRxpx45dI
MMdohe+n47Ck1TNm3JMk0V5qf12oPWfNSpx3lWMEj4CUk05kaFZmuR5WIjcf+nGn
+X8IhuzRpurJ2/84RXuwSaIfhuusF6yDit704whiCUu9Ffx7O6iZLRz4SXtpmcqo
v5Dw62VQWVWmwOLBFJNZeL0kVmmlH7ERkbtuPejSWAQDmSyISkZOM17ow19QrfrS
tYlDQCkynncEvKDLTVBas2p5dvQQFFpULE7mBBR7+1w0OO4tdCQQ3H8i2wxdqg1R
nsA/O0OC5HP9yVK+Ki08iSHUvtTGmoVcdcSXBCjdaW7IkydDsk1A0DCvCIVu7vLk
X3sVzW8G0XKFJ4WzWXBze9PWd5gm+KBgVNFqclfYU+oJksCKxFyiRIK90W4CmfOk
DuBFCjQzJBjAQ9aVb7Sd7qCCQ8NMtePgiFZp7jDEcDe5Pb/V8H+xXLZSVAPBFnK5
Iin3kwBjGX5YPISF0ldIqCkVTr/gDMOZDQKN4hPcfgolT5yLTfzCrCG4FTb/K0LO
u8SHHkY1AvRxpR7SoU1SU5hvhLkINDoegsDauSrRPHA28ujghUS9USvXfuN8uGZI
RtoDkiSIcvf80gYfCch9l4tC9I5E65HaakozMWckpbc9twpq9Q96KBWQs/wG45Mp
ab4HhB+MSC83qzkZJE/o27GlpgyI/WWU3BCcj9HPtTKsAh4px5cTMr2hWN6NXx+Y
QMtP85PKZQ5r6mClJaNfAcTn54NaslGtFzJuTabyRL+tIlsXOMXIjvGzE3MzUWqY
Rej1r+A/C/GjQFrIeOehzvdM5eQdwLaOxHpgSrVmIGAPAdNmw9vktWze+sOrBFTt
4NSZCjpr5qoD1yuvv8pR2mcde047or8s4enJoceD3YtbC8GUFDBXG44vuwS31FfD
olpdjnfY697+2htnQUg0amI8aKHa0M9Tq4AGoW9IB6L5Cq7FSTeQHZs3hHuoNE3d
PpeMWuAcNYWiP9EiOYfoj0W8LThPLiVBf5A57Xp+Grc0ibFfbr/LP2yHqHI6ykJw
2J7N897n5Q90FGi29S3KdKY7ucVN0afgCvN3f3hdFXIkkzpMlGPwefei9Rm+bmaI
FrUzwiYSmUKt2sSbwpQ8St191pY2tum8RWFTntaG8SVMYpU2Tzf4W06KsvN90FpD
JSRcTreqlOhSa2N6wDB9x4FZcfr0o0icHiGKv52fieddFy1G4unvq3qXNjMYQr1W
7eEUBBa1PJm7JTN2xu3JnTRbFoduJ477LpsOrfWZeOnbeqiIoD2pQUIQmKYgYthX
oqIfzAlFajlyw61b7bDtH1t2fEBvY2W4lg3TqpTokzvsjIqIuA3JTGkvXnXhKBoM
h0RmmJGpcgsLreFLm3iBcPWq1oVOkE0tcEOzokSYGkE95sfG/N0seXs3X7myKG1l
qEaPjCFubTf3vBhPbz+tWDBJWgoXDme/6Zs243981j1nV+z6mPOHUrsBZ07ghCiM
fP2wVh5nGyS6ngjImPdWTnWofsjEqg3Sa/atgj9eDphyp2eUbCzmOT5PwlInjjyw
cbkgeRDuxIKhdhZgxCRDBeoXn4oAseTPwn/F2rorKBUUDBtPDgmUCzkrD5K3lrDe
lvuUWt4Ppnu1P4vffg7vJl5FE+OvEBRCwyJWXvGuPbQUPeQxQHWDRJSc4abZP8vJ
fIFutWKk69j1fwhQCR2h+cAp1Z6LqBbhTKLlkfmBxHcxVcL1ShQ2IxoOOXLKFiAv
6bhwnVwdYid3Xwtcpf+KFMf7TMTw+RjdsR/CzAcKVGOaqZitTC37O2aJVwTY5mmT
+e6mHVXX1ODUXf2yOQ6vVJI3XYUrQwC43UxjbK14pmQdPlqw/SieKPZ4+Vrjv3X2
uxjc+9jsrMf9hh68K/9b4qZ4l/8MlJrzEDdht4xacMzlE9zeknJVOEYxwwOdRGmR
BkkW91xCKhHC4QKYr5qrl9s1qclxH/g6XfSCOLh1aQG4nE0tHLoqpOXeSt1L5ojZ
Sfv70IewOBsiz9M8siD7d2AO4SqAGdjn+q+UBUvtqJr9dyWDsr5vNqTrrT1XGr5c
m55K/Yhxmh/9uvVSFTZMiwD3vlbnDUveY8gR8Bgb/prr1jqokTl5gdtN08LaY9mt
f9iqpFh/EP1KVaUJcR5ii5Cl6z5OD/xJfT5O2QNCCXdzmJt84GBffQy77HLFC+09
YT7gCyfoMmD4WJKq8udbuH6E3mcdYTzaAowzm+dA34PfiezEJH7bueGLLqz9Zw1w
djX7yOBiVVS/ADy9T+7rHKSL00z1LKyyfOLjzwGVy15g4JxTljHMn0thuwZa3I7u
LFB7CBneBRMyZ79VQQej8p/SUO6lxPAThAajoEAMRsA7R1ip8toIg9bIIrGhqPDj
a3HrT086uQ6pmGMNDKsnXLwBqFhEFfGHLMw+qvMZnxi835k0RP+MMZ1G78UyUMqK
KozKrvSLTQE5waJ3aaPdu9N9HR6a0YhSfeyVcuT592HacH+WiUgVoZiUIJX6aRgp
ZhHmfpaWt+CzVucREu4Z5DxMlUiQ0MXvvDKLl/d69ReOzSh1ONgUbWh3jGU6S03z
XF/uWMV7ZO44/2rl+zPw4uaHkrGjtG9qpdYTqb50OtCF8HQ/sjknFT9R5FS03g0Y
C9j9RJViopJ7O89uD9ytzh1v+6spFcTGd0qCXuZvW8rM7NDYvxrZIfHbtpInBkTt
3w7lcYOzg8AeHlKBwwF0VTYdrSpawIflGMxX0Be9ixI2i1zX5XB9etSrUayO352R
RG37z/pOeRmZb2S8pHEAoD4QC7omhOLwXyN79hHBtI+H2bXnfBK5G8BDVDYq8sBc
EnputHji+5mykvbsR9w2DJhoUuvAzdQbibrk187TWKjP5XAAoMNQklUIsJ0EEzmG
zna2EllCD+NZUwzlacK6ivLpAIch41mbmvlb3GGpQXWLOWwx+Yw/L+irxOzdNU/Z
Pl1aWCu3YI+8iyyQA9cASTZJacgNiP2+btfEZLjiyKo583thEUpoXNq8y4RPTu73
MTcd3ctzpDKD0e8oXHjIuEgH/LvHXze7J7uOA5O+EGxOnEAEItrq0RU0hOdcuyht
U5s0nakaFy8xOLbnmSgwGv6nbIcqIhWzUJiS0zyL9bXZ0ri/2DChf406Wzbf/rcA
JYwiLgSjg3hYCPrduHUhCvJT0cUikVA6dWPs4/D2M/c79c+VxzAjEV2BBJ6yU8J8
/W47K4MKtbSnkHL+DsW+DyrsUxwsal1QDUXm3sQxxMd2U6wVjvI33S529Ts4/rhj
qburULO7a4FVw0/sDqa9huLtT7Ni6vmqWvSiQ70UlZMKl6IfHkOxIXFLOYzn0bwn
U4+Hk07bdhx4tUIu+rqBQacl9W/SmD7YyQ+r5XxSuhCBP+BFVkGjSarGAJkZI2k/
067HZP+JVr5f64D2/+l53bgSwGaCUIw4jOYEEGG1etMohmNry+bllPw6MJuiRhuh
WM7jQCMAMxChiO1sQZ+vLkwV2EnZIEjrdhxQ+rnxz7L6qkWUE8rlM2PlON8LKHPH
97o/chrKf+vtA2La0v8JlDUtYeN5ngmyZY2UZK0eNEPy2fa0OkyDnj4ptwxvOLKi
+tjn82XRztoLIXL7heqAc1s7dPE/UwsjjAQqcT4AdCMGaDr/F2w4BUPJj6uQgkIA
i/YO6GnnNcN3ueMaWFg/gDioD1ei/z+kmHYuDUP50lXMfheL/5I3K25YCviXVt8z
2rRildlRYJTjVWpT/0rNJhZ5NFwnVyviEqPUsxSVPXT3qcUWt/rlKiIfoa8wS0Ec
9XX8aqc5acmxanAE0aWX97syXICNAItDAXHdhNOLnPRMBTYJDL6XvygCoHpx+wlS
A+124rC6ogPKgip7SwIowGixFTf0uw9QArUHLJqj7s6mprcIF/l5XPZdhK1L/XXo
4kg6HAQ3B9Yb3LdI+gjp5jThLXJORD2QlEd6pk9BwJslvCa2lfvF9MDjTAsuEkSX
mDpmt4YI+t8tA3g9RvCa99McXBDD73eshMEkMUx6inbiBKl0cF295ymxuUaYAaLG
mEj3xnijr19x5bfIyKTH5bgt2lTYMWIHTrIzepy2qQ8J9AQSjWFyG8CfJcnsfuGI
XgLx5svVDoyb6A3VJsDuP+RcLjOosjDL7mr/oI6qbsb3VbD3HR6V/flJ6EgvnmyK
5Ul+nngY3UpcnqM6aw3t6bJbCxrWlPGA0f6aiX2fUFp8sxEcEWML1Ya9tujjIPD3
Nqw+hKYW68qKoU3O5zugpEA+fRrcGd35hmlz2y0tvSQK5qqfJxCDfE/8mWfyMRhT
gb4gk7xOAr18YnGXTbjcm9W6qEeZVRXhYlhvLUC/YwKjvS9sB2oU2q2iwfWcXE4y
Qt5FN2SDjGx19HZy5qQj+9Zx2R+EdPBnT4YELvVgl+PgkSTZDbAQS/Xyxv+EKJdp
D5IZVNTa71+hH5qyW4iQ2qzTIVQgKTSzPjGDHzeAUxmTnZBvKxqCMV9U0jra0YPj
RahDbGe7kV/FKKsxxNZuXyIL8gmEwbtkkTVPxJDbeF5HNHyrtf4UbItgA4bvL7Nb
Vd74/qhsyU9dnCAIhtL4a1HtFJWHcwfItLrornC694I/LCSO4X3ANa8zQh83bYJS
EwFIfX92Lpe9VmVbVQ1md8q9Pk4/f19VF8dZXBXGuj2Ez3xoYWbltLaf6sfozrSL
Yi2homeFI7/3+yj3P+3Iqommom6FLJrgKrgwHGqAY8Ab+7ChzUCXz3XdXVZ0gP/x
rWxGNnF/ljjADlEQGZevcyl7cZXw35glDGTv1wC02aRkc+vRY7JR7ERrqq01aitc
yHkkzedYQsPzGc/mFTKwNrX4TJO7iWTjrXbMb6BGmHcNnMCEC4YNwneg9LOCqyMS
0oHXqem9dhwWsqFMGP88KXj8Cnic/grfau4Xi0Gycyloroyf9tBmIWWjZvmq5cu4
g2aHqCudDLsbZ8Pqe/k1Aj+MyeKeKg42g4UpL60n03HmE1LB505NACfGH53o4RLN
AG/2nvyyu9acHkOFmwfEPfOu9IeM7c1sKGdbLobcLDM=
`pragma protect end_protected
