// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QZnEAM1s1dyKVh/aL0AmWo5PoJCaaMgewNfrMTyDBdRBhdseKYEWN5Ok0zUwWQoL
cBnXaND2ktQMLmyo3EQ03C44h/YTF5MPTFa4z2N8vK2zXrmjrsiGbI1A7v/At2TS
ByEF7Zv9Wd7PhsCahIxxDAw1xYX1dPcaURVOnEudXMs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17968)
x1GGGT2ck8JYTcHYlK6OMnf6pOIeaiRnz3h9G3dwDkrutR89oahtmi+TLyyuepvG
D6YB+ktSCUl0i0BYL21BLsrdjw3sP7qcAdzD9ioHUIxosJtfCwOO3bHRrqGm5AD2
8VTBaj3AkBthyxiq6ALP6RgGX7ofyUqOFt0/aO2tRdDlz2F7OCeJPgdfvSFgq7yj
9hnorgqa60dar/G0xvA2fDfARmU95MlZuVYV1JMio33jBz3AAxWIxukM80nfjK/5
z+jpWlq5nPrHYu8M7ZrKHINntobBBU7sb/RIOM84aGSoINzEWHFpDTzsmsQihcQR
9ans9mRbXaQJv3129PB/AljeeJO7J5+E05tMD13xv9/oYUN3zCG9uemgNMCYbxpz
qz536Fmf+URovX0b4f/OWByjQZwXBJFWnTQkhHOsxhrXnJjGGgyq7cuDa1BL3EcL
AMEiqTzxeTkU1QpYIBprwnRFVbJF27kwZozvCLfJOCZ8M2U3AezOcLIiSvhianjD
3zFZxni9m0yy7vTJ0BEK2o8k8XwVruWw4Uz/0X8mrN5G0UtAp+QKvOe/Znod9yC7
jpcrdHuMalRrsRjKOz6Lx40DR2ABz54Pt1urK8cLnQg5K1TQs+UWVmXLRFkDEJLG
FMHAvs12t9XNwJo7bqQiozrqfMEDWMmLmpaTmQps8xeR6pBKi0424E2N8UdXIXOf
uKVD/6rwSSQwwBkT35m1M6lTmjK7wtGkVm3hrN6jV8Adf5aU19qaa7gzgsPxzkoa
aJKo3y+YM+Jwz4sCawUrg56kaa2KrUGeT2m7eIvikEM4ujkmZ14snszimev6nItR
ZGDVMeveVyTB/lq7VA6mcdC66v/jHMp9GR26+yzKTjZXtys9dpxsXwhrlDQhNS5o
PXH/1IX/buyuAG3Sl0HuHFAzMo+Jof3AnD1reOCpAXeTi/2ZOpkbgBGZQj3NlMPu
eWLPFXxS16GFlNIhBgUDyl0sSuhXQkUaL0Vx1el1OsfjWpgVTN3DETa1sh/zeS/g
+0cpl59hiLZBer/97+LTi6hlsA6mOLocUmrRDoXpK1jZvqOiwo3z3MXbw3jxZgVz
YOeTX3yzvxaNkOG9k2IlVeRvqjaRsY7KYcPloSbWVZpvNUZf6hFsJydwyH5t29la
hgaxYEig3/ekQdOoTohrsQCO9uNbHSXDBC3EoLwpJsvgx0uuZmb6+eHF9UEsV5dJ
xrJGrOZmHpB4uA49saFBUzCglN2Nk1LFVsDJFZBgtW4rWn4xzKIKhpoRMB76RufA
RgJ7BR6kngTQOVEyErdCaKlQD+Vzr49/IvF/NJYxhNw36yEgMGqCRPl7ZDaxBo08
HmfYo7YxgwP2t/TgW8NBNkdVlNZwA8FKuChqGb3Yix4i0sZzVMXLyrnInFECpx96
U2kI9r5Dd1pBrlgjN8gqJXLAQZ/NsaNqt86MKOIyCc/5Le5RAcoLoGnDwwJQsA+Q
aJF9Z4lVhfjFdiE/nke/n/s4VoRQjSyE1VY+cJ0aUAI+SoY5WRK/4Fx+jKdmk+SX
9S7FW3A3LboEgqY3D5Cqn2QShcf5uNIHN7isXVgaB2mXUKBqkVbR1buQJ2kZyQ4d
1iaHHIPLUov5oAnNctJ0ftj5BBBdKMoHK7i/MpAJYahFOwtODE/iQN4iZ91o8VAK
FSkXW6TDp6usW0o2eTSMoP7jwPxHB4P8jhGIIosL8ZCmpUkjiGMqRP/WwrHqMolE
CgHvZnQo3NfDEiyVTq7/agunk14fskKurtt/aX/1dpyltOz0DUXL43XjkWT+NN+K
Frx5J9/eqV+2KWTHgN2rZBJp9wPHSm+Z0SMtPclBzBehu0ZdRhs9jluVmFzTyjhO
zON0I5TtAZpwx2JVv7wZNzGHqF9KqTBjp/2y933YnmEEWmSjEEs0AZBLuV6SyleA
Y9F7u5D3ORb/2O5h0FvPQavZ7PPeBH41zCHG7CU8ktTikbcGbspr+ZFinWF7XPoL
QFUzDL3neE+kuA1Kh6tDcuie5s4K94v14Ek+7UxsXV952q19iWcnhGwfMbi5yccl
2gzcayHsoXKu7qohoXrhREE91KPtmoEfVzb/JcfsnKenFEkNq/gGT9is7RjG2zcM
B7PTHJgfNETfxPn+4KdnHTHP3whB1DzHZqAbeBY3UcdP1tbPGF7Zewq/8nTt7x+Z
cMSppt2u1SEU4Dy722NxupjlXQ0p+lwE+3EnGENUyve8dovSbB67KAjDBGKSUtYa
kKFYLRKULTfUYNKTyZDWuei2hhzlFvwRiGXGOUDmxF2BetpL24BHCXuVF78dX+Zf
QVEOf+gvrys1aFhNYPrFk2yOVON42EUODTjmykRz/1C9gchg+0Eg2Ruf1sJ1HUfW
W/EOhGVFyAXFjnskW9bPCn4vBfliKJ3y1tzxxGk80TVZ1mP6HaoufNQ6fDBf8wAe
fIEn6mpD/itRWOPC+2xmWtslqsWo2HQoTTuchdj7LQCDpH+Qja5uxc+d98WPhLM+
0sZsm9/eg02ARU1uXmlJPHNJv/w+X8LPtCFfGB/LJynZdQR1W7JrLqrxj4jioq7O
co1EqEH3t/Pg2nch9e9mR5+Z+ZiNwJj6Ox2oVEi5XdArcLlR518BJpVWgU8aqmVE
pi9U9Wmk+kIL/DPzcHjfNmkfX4QaFCG69m7sVEIv9sxH5SMGRpfn3Ur3DTo5XL9K
Ydecfh/Neu9hQDWfE8hWwZ7u58yBDbeiQM3ZfIb9NybkW9mcHLSU9umnwivZiVln
W3GiuEuzIKfPN3/GRrXPZAOoN8V8v7UR3VghZnkEMjqU/+70KwGCNCfLG1z3Zk77
VCulaHCrCnDua/rqo8kAZlO38WA9NKSVUj2j5CWJXZplh1+Qte2LbWb27htla3Wc
e7DDx7R5FeR81XkTMgzPjQsRyLx762We+4qugWLO5UOTNNMkTMwK3pQZ2OTyHkcC
TXLyldLedS4kRmM2kC+DWF2qUlisGVom9oTSr0+WmcQAwxormMdKXssIORmU/0ym
3NBzVwzPk1cgvXKQORi7RJrTtACZgRu1urpSTylmtyjA8XokN9TCHkhecOhCa2Or
OT4FxNid0+KrBNTqDMaV0uHi/YAAPLGHOCTtxwulTZm9pVfVBwP/BoGWokwSwJpC
oHckzv8dbw3UvVHAwPFc8rOSJ3qkIUqjb+IKKvAt6Kj8N5Q0Ql4eCZcwMGyTAn28
IJktwYiOVkH1IhY1SU5hhQXMLOHtzkT86QU6SKtp+UwVmXduTLVxFnOfu2rnI7v6
wFE1vN/pywp1xOqGs5KUzBPElYnqaKMWLFZl79GdZCKG7t2dRBwNtZv/9Nlfi9YK
ubJvfi35PnGtsGxzamg8Kz/xqi7Htcwbu7JqxGmovNrl+4hxLTZdcnotj/mut4rm
Q4DrcJeERuv7rULS4ckF7LpwqdJf21UmXa69N8Wk7sKKhPJeVAf12SKtaheegX1/
WIq7gXPqSEXyl155HN/p++o0ZYDrLc9xoOwq/dRdLCCqMp2oKchbH/43fHBQ5zBz
IefR6ePofvHB6v19Y/WGUIzw2me0FD9aTYVk2Ej0+EocUFjPZ7P+vNmGqjEFRkxx
3wAoNe5N/khizxtxUxS08EDJcOMm+dcQrLXpAYyGiYngXRv22itSe1TYLU/VPDTT
1QgqDEprawy8n5b7O/S3Iz9JPkAkp3WYkm/rGufCnW9aXBq3+JmAobOSnzK1uX1e
cru28hsi44skdK40CsvjCekIaP9TWJS88hGErv6cHo6sGU2uT7jKs2ZNTrA+QmS0
d2dQc/lhd8RHqNzLnYGYnsGoWWhPkl32b8Y0/Qb6rkJPGjnFWY9PJ+jVKn9GAHYN
MxiCdBUx0TB7kva+ZSRWSrXuVZVFxNpekx2BDGb6A+j9Fy0dcmlXazuYnv05X2AJ
2/PBJ73yimDYPdUqnMjTVm1HINqhC9umitS+uUL0wFx9f3s/kcoFy6wuk7remKIw
mGv0YarWGzWPeE/3Q71KC6usIOcZIU5Q9pq3ssBug93o89zQGSIiJqPVvBNsILqm
m/9U2QWOQ7U2pUWnTHD9O5CsACK59G2NQUwMO+16txs7sDwOIEulFcsrpEsiKh/Q
BWBwNodTZhPMfj1VkCxcM0FgX3K0Pazmn8Fmj/bzPXUBh0ImrFrMAugOkGYbl7Th
tyGcEocThzK49pWwFm01jHmWzp4a4YkRUtiAA3gD21f8/BnoIzu/PvpXqeQJXCiC
42/UibhLmVnV5darsMAs0hcYKsqcnfHNEV4jRHuWKZ0WFcfwuFUOPKcTvr6NPjOO
/PX0AM9Yk4n5HNawLfG/aK7uL1oT2+iAp5kGKaScl+FTgxv46AmYsL/9xv0aj7oG
GewKU8Lom542E8m9BBI0Lm3gIfNVIo1KKZ9AcKOfp3N/FSblb/rjoJcQbJj/t17A
XBgZL/ybryLfXeujVY//Y6t2rHp6qNFBzHRiAiikD14Nb/5Yy9k2Oo04bS5Wdl5w
z9qaX8b0G3/0BPwd+VsUgIIfJpAZJmKaPiQd+a2ayRp3WSgz0cU4XiDiBpEYPp1D
a3mlJlv3roQ2UGHESHGRUW+tmTji9TYqERv5BL2g165BM04K5k/hM5hePqNTKLPD
6Yzkaf2I+1hWn+0cpwdiiFZns5sKi8ElPkpSg6bXef5Id2ELBr0p3U09rNzyfv/Z
086SWUBJxlVpuo4pQn11BRde49KEzD+Pevgk93dYw9Lwr5aYfI618BbIUwBky638
iquliO0t93ouJQIbuwNubJi0O0Mt7e/teE54O9nQygTU/KfnkB2TwNhELtdyRV43
pUVNqFEg6mkPvjvtfGeerzcMDQAq8EZNZGi2uDPJrCDxVf3VotYat/N1wr6783hF
CaDouP9TMptKqPDYQPTP1oIzXgQmLGUKKLuijJG9lT/133v7yjz7j+EB3q+4qVXu
1Hd8VKBydc0beJt9U0d1i6eQW/LgqWYV67WoVwpZuNmQVr3F7jk/cJPxgB9PaFRc
qFmGlW4fZ7TRJ0x66u0FIOX5k3ufyQi7aCDXQAfMG5xdTsuob188xxOSBbJ5TXT1
nZ55Wl6UDje+r26EnsM3T1rBXnqkOWlqWhCednDwYkZijIVPEWia3SVwIL5hfNK0
WoM+cw0Ku0UGt18yLjEC6cXaWLTTQg0ZsD1wDzWPjF8PeYEnu7w2k6yOVrGl7+SS
Mikod03a9K0D51ymNTFw05NT2MKwuMTNHW6zwUgEJGWyq4cwIwfc8U47y3psjMvr
g5Qz2eL2NK17u0rjZ7RtTHUwiFCZqfO7g4CbTh3DYlu0YAgIP36TGGVdI7Fi25pI
c1G43M5WEtLQ6QpS6lhSLluIchWQyfPATvwcvQSx9eZ9RfqYKWORjOTrjkiiMZD4
CuClMw/bDve44N3JUPKjcf0/KGE+GkH9cXwBFoObkfY4mXkniMPBlk1WMxQSR0Ff
QdPlb4ko65l0Tddegwlbucc7U83x4xiOXMLs1cMS4Ff7yjlqHwNTeJtQ8DjF7rKr
VQLDu+NRIExA7X2RbJtMv9qFxRWIXm+wF/0MfV++5K6ZZdDAmrmU2/oyjXsknMk3
vAqevfiDDDiUB7iSfhDtELzybx3rGbmBlpyqD0I2ny540flPGVfQibO1OIF2FWK4
Cx+nx9nfm27s0rBlQBG5NaKMlIsuEoWT3ugtqBeFAVxE3E1fgen+xdpiOIFgEMm2
FSKB+2x/aWGNHqSFS6gAyLEQj/eBiNNuWRZJ0//J0/00uE48TJb1bntnbSfoMW0p
af1e74IgpGzhvp27pc3WXiTS18ImeVlVWbo6+riJAcarlYd7cwd608l9ghU4b22s
8BV+a3/jQz6MnnXeotirBY8l2iVihKSxnEAysG5vSdWOcOUJUj0hrjs5jKpbvwtP
zRQOsOPSZ09h2yqparMLKMnVW8GMWKyQ899BDG/MkRc3QyxkofU+o+3DvX2s6PqK
LNc6gPBKBOVQGGcSbg+fhY8TiQF8b6dLNOF+nENPfbDG+FVyzZ1yncRmt1bIV3Ok
KCcSCWOvBSAr+F+1HEmxIP+I5Z0wpd71srrg5nylNOuknroBWvef875YyDtueynt
qh9yiKbXqbMkH4HorM8M6BoHcdZNd/9fXh61x9oK17Zc9y6IeprQ8tBtgQkcRnP9
/a552Gauz3tkbRU1NxXsmgOGtxVCavlMtgupcehTvvJPNhh6ttw7FcaYauh1AXj6
qvoD1ImkUch8FsVSI7HkkQoIYSffsVsOs6WhJD2CxjAZtOmhtU53so91K4RI+SPu
VpwMFW01bg9z4DpbKM5xPNiZcgHI/2HawnMALX+Ik3HQy859jI5XJxQAZvxOxAPO
ia2B3b7DjpBboOFHgDy8VTuDziEwTZhCG5Hcc90nsdIEMz7wHfgeIHwXmBh0ZJhk
aCgTUSAUyEJ79JMQdpVlr0Fg5kRBn+aXJxDcTkn0k67azr0aW3TnreQUnH7BCi88
QiDYj7ioy79mezCaok2JHlPv4oVHO2h27MX0wiXJlxhc5sUv6S3SRNFYxk/x0KW1
wt0MPbebBZR6n2oVtUSHNkoBhfHZdRauqXnPG4qc8vyaC/MDjStUkD39SSZiEiOn
qVeDJuCVRM1Uz8t4zVz/bwBXcHK4zUvJivRmerfCdWP61TlQS89N4dwwgJ09FZwL
0R2k7zdb1UIIsZCiP+jPSYiNF/SFmycrMR5S531Y8KcN0O7sJT/aTFfDNBPFOnPL
47fKs4JZmXtS7XI3gp7WhNVdj4+jWYtaP5+A+DqYgxKopFa/+RNl2qcoh8VxLPPz
Yl5YoA4PC9VNvVBO2EQo5utfkFuoEI+7Nw9GC//xo3QhDKDadiy8RHjRsVTFDaAH
TWuwreXJh0galRclL+r1LIS9gKBbZAR1xqRy0VMRH34ZedR45JMxDW7YYrmniYIx
GViy8RtDahUYSHwGjm/LVRc/AbLosUzXxRZhFzeUButrz3W3Ezq1NqNzuSMhjxkr
9mZR0F52vltKPcjsI6feAXfhUUFvCM7L27OVDL/01DGbi/HBQSTl5n2NAexVHmRD
0vSkYsMNzeEJ4aDpG5EtUK2HIiytSkqMZ7cJx9xknZEW5THedsdaR4sPRFITFMOj
4tVXEkKqtrwdOMVrXfh9bTYOtzfJph+PXu5fNEtA69P1y0/QTDrM1JXA/3VoGdAO
Qz3FujV1fPiux2S7VOIt9J1YonBM6vbmXtvJX7EBSFczHizYrm1Tbg8TrWO9Vm7E
e94KA8CzsUCznwNcFTgecyUKpIOW7uiWC0G+IxkSV9LKVs5zKS026O6wo+UWkbOE
LT4xICt79+WqMiGfBu+CorX91L+dSRyVLfiUj/mLtUnlZks4QsPHSuECIJpeIH+p
ut7euKX/4Noh4R90Gz7Tou4EB5PwigKFOqt2+NavtoazBkUcfsiHwq4rr3PzFOeD
I5RKqqFNIs2OF8ddvoNKvd1OXAgrOrW2oC50yE5Cg77he9RKgazoZAgx/xbMbBOz
Xpt3VarJofZwq0fno2jzfItlRaZcUzAFi8XOoF2McWvHqMH2OavcKQ4qFiZmOyOz
TEzJQCmW+VWzR6cRbYH/2a0LPnIaX6VagXfFKes6I7Lpxv7o+mVr7kmRkdecHzaI
cd8MKbbk2Z/C0Qy96wCWVH/gsjG9Bd6/RpcjCUhlJPSNA56RdN1OgOHEuoetDIDt
Tlr4VoaFVdv2+q2gjNGi2WBpwsXvVpm4Vq5xJsldARmbBBr3/ln49RLVEmg8HGuQ
JFYF6JBOVaIkmcc8fJ2+KixcD5adt3fqJSxOMmVCX71QlvnzUnUYAAG8sYSpBk/3
gaw1OFAlgDrQOq49ddctrc5tVnWY6I04s1EjfdUGpI/5F7Sy6zzsHWLQKvMSsl/q
Z4cCAECbxpKrisxAfX68E7zkyEgd7uijhsIuzIcjTEanGwMgbum1b4SFFn4lvATl
81iewogmp00BYgjRKS+l06FXyGIFAU/je6KQiM1CSSBw+F9FBiukddTS81dLqPpJ
sTOqzvVsVmHGhQ4wQ24e4qPQw+bpXXkymMAeyowbWz+zWCIQsFlL3V62MEoTGyIX
GCU3c/1LzMib9waxe7jXUIJdJB0KF6g2sRvBft4i0LJ2TdJvbFeKdBJjNAL5Hysr
W06vd7xPLeuQdiyjXxtSJ1VghQkhc2RAITV+iBQVJVODdD1wqj48hgGK6JkCii1L
cxZti4HhCtxDjJP7I880ILd+dZRaeJNCKqt2mFFuaYiWYspRiTmG3ZnIuUE7xbXp
j3ktJMj875nRKGCiclRQpEW/RyXK+3KLG5+dYqM0Ug4AP2nH1S0kHyEM/xAlmYc5
6uKOwooYtBbh1fZLcBxvzBg5Bzg6tiBXliIik3b2ASONtAULAWk+Db2DR/Vs7CxI
Gq9z0FhtCZWKDf4txW2m484iQb4nWC+iMHX+QSx68I04D6cAHAzVXOX3yTjwcbW3
kuNis4QBTeHT5ZXmKKrYZT5dgGf4m5th6tG/t+pBFMyu0mEC97TDBCmdiJjKrfQg
L/AcvG+5lxi0OXK13XOR29m5nz+zllefgiMYZXmYvyCxchx6/MblhVQK1alAbrf6
E/ZKTExdz3PtN59cUWzhDUI9AvGoSUB52mBmbCcWAGCcJevnwaOdG9vhs0KcFZ6b
UEvt0jtr+H+/tUrXM02kbRZRK2bzqOtGovDdgFOkw8dyd/undXN+/NS9V9Ob7t51
J+JXWK8v9e3GouTJh8NwCDHSVY5+aplTe+PHymdH88pkVqlHtKhXH6ouaapB+8dX
YkAP227M8e5SZ2FgDYhgnPFa0q2e4eIAmu59I3W6wm+N/mQeusTGtxSClWmUZUJp
DnqRAQ37FJHCbqDaKIdem4EZapN0lFgOtoAhl1PfpxCrnCUcRjgLZlxtnvwXisi1
0cD9fYqOKNTpgWR0yZ4qOmnwB6OzdY/3/80jU2LkDqCns/PazXTjbI1fDalm7KVx
XKvvAPVeIIYr2OFPjQbimuucqUbe3p3UTdQJScKC+5kQBpDV4+oevjZ/pmu6Ytqr
kZvOEkss5W1f8WxYLdsHLIg0JK2FMUJoShuSGKx1TUmRYuLJ55AufM/iKWqvXLep
hZwF3YUrpZWuutoezpuMZWbYVeKzV2TveLxDqoib5/fMEK/YIy3Wb6//gva74dii
Pd7F5phfumAh8BWQYFVUcw1k7WOLIlwTxd1LdmnfvaJHBxDJyf4u0I+OkGAGWq1O
BYLGnMb0/uSY0E++oCAQvxjmfVAgYZqyG2J0nFQo6jihGNik2emewQRI4DTvH14r
udlaMcAuNob04YYM9SSXmlFmPOQJE28Lf4c4AE1mws+x6gI58dkXDe7v0R4laR/T
2hFWJfPOAnIZja5qcntUuY+XuPPG1GqYwgOr8rJVADiQDMtHtEiRPr5C0tvvNomi
Py0opPEAKfwn+fCzRYV6C3WZ9EZqg4XVyqjZy9/mEhwJhdQMO8tFM1y416pbYMo0
iVRRLLtAypwjmEmOryLfIqxmiQAKFWTcZD3N2deabjUoXgi3aiwvZuWcD7/7mpqP
fx8B7q1d1i9Ur6Zm1jPIZDFO9jK9lY/G3Ssw+zyyHaqansIJH88Sm/zKTNzLWQli
EVMmK+OD4pwhcDrf+p8DN2MPaLnSjzukyJuGtvDq2mmmnaIswztVIkZ14NhnaadM
1O8PAm0wYRlanqf6gaewabCzy5fqiXTgETo9OH9NQTa3OIu4GpgSaE+5z7HlmbYq
w4Liw+UT8CDnl2ePCCMZkI0GDrx0tbjifmYtdz9cip9cGaMzoz4/J9/dPL8T4B8c
O+vsuINaaMG23ZLNqilvCwDc0pC/DwcepLYGKRm/qTBwODf2SUpD5CcjyW6h5HJd
i2ZFIzFn2z1P41cLVND7Qv/EGZArZr3al16xkY0cOtFN8OWo7s6POmRYt6HeCnu1
sB6vWBZa0yBwoyB5Zs0BzqXn/VZD4Y8vRj+kqRWU4RtkV+khZDJmcly5YR5GOFkK
q1U8HH1Zk8peutFZZ6CL4MXzdRdQOMpV4r0CIqxta2OhY/gqhbtR2qP2q2ezX2AA
MrB0zKHpCO/BauoTtp/nrXWrH1Hn74zqXihr6plBBK3CXyZQjjATNyKZMimq8WBi
V49GH7Vllti1x0wOq5fPLUS50H7ezv70EvjGrv+0k95rH0y6Ey6p6+vIrtXO62DH
8r8nbES/aS/9rkpgGrDe6KvabJ/3+oVCmfvQhUNBSpOWulpWy4ZE4cY+qJNdzKGL
qY3fZ/Z0zcbkCUzQEEPg4rjO2tDYspkS7om1NAZIcvQ/ITAXi7mw8NFVv0QzD3iX
r6l1kcr1g+glkpcY9SwaedttLvMlroVdHbNbbR5Owucimkcs1OKFCCBn5S39EeMi
yAEAgHIwkVu0XecXYmzS0Lm9wpLPfwTCXb0l8kC8bQsd36ayDcLpuAgegW9EKmtR
HkY/eixnXdUFJiYzVooP4dp8xSgKvInnDp+sJOGrNVbXcmhEb8LzL8O4+/Qwx5yF
Fp0tsw1r/j8unq2HeJw5VxlXyhpOiHm2herLLwNTxt3ZiznhiRyAeBHOxoPEbIHN
AibGuLTCD6fXuEFzr8drq55V3tFHuzEZmPQqLravuKbUoItBxqswwTQG0vGSkg83
MHz9u6zuTvLqEanOM0A/dZgndWi189HvmNXrN9HiBQpynvUwfhipFd7AH6VFv4DJ
vIbIndlr2l2BYJypARIL6g2R5T0GGgJJF5cryOpo1tr6tXQ6fQggv3QRsbxvJOFD
LRG6fCMurwz1pl/whULC4F97xg8tZ/5qn6O2qX+3xlCzGJYw0USHWuiMnj5rc+PZ
6kQBd3ZjI+oAUIMdCH6YzOWgmttktQNLqLGUqPk6CUUiRMYcmuevCQgBekbI/DgK
va/BiIIgwNTWLFfPVMHHg8Q2rvDM8qIxH7LQnqtY+AAWQ8jlgY6Jgcdt8+exOKIE
cNoPRSH9Mzjtp13QyQaRmsQLVcAQS0wyfTXBKHkJXgezxrwLVZiCDGasHEDJzjcq
J9zuhce6jUoa9aL4raaZ/hib0oKoM3ST+JN3dS8IrgAhstSB9KU6e4FEoIWT6G+M
YO0sR7Hq7xiecqAFkW2m59rtsddu+BBlwLb0dyokutVBiSzGVwCBDu3ol7qTP4hc
XCD7BX2mH0xB4tlswLWQcSRLnb9TCjI47C5kurMaRvDtV/VVTtD906sgCEmWIOD+
P0IjVl3I9EVGclg95wTe0qWTGRVGD1YJZ443EE2R8rvL0JQMz12YoUx8Aw2Qb6PN
CGIzcScuilOK8YytK4qsFQxmCLSQBiFanlIRj6JPM88mVMArdetQL4eHcEz4P4EC
ygiPX+lX374hAYVyO9Dh4ueqQAEYgbu3R8IF6bjsi9ndK9a/MWhuyKvHyjTgYMgf
l451RDLJqalNywr2cHvfzeX0MhpgKc1VNJEmAVt6O2ogYMF1CQN0uMBca/0b1guf
fe7bvF1NisMuKwim3YSpT9KOCBYMK/He6ykSIDYNWoblo7neGrKJMyPv7pNanlL5
QvJb20YwUK9/tjkJYIwHHC6d1PEi3DQb4OgPQbb5o018raHwxVEdBTGvuq12yozP
dt5YEAZbigXS0X1lV2TgDizDnNePX4ta4oE4ehA3agh5+MFLH9vvZX/hzDttMiTZ
5teIxvefPP/5D/rqpAgiK9BFDX06BVTtgODenrp7jvrELwJS332peHq7+3YnZOiE
mR3nTYYr/x5WKCAO/tq18D9YBzcSUHnw/+ZCRvi27IGLvAoWDAcWyoH7UuyOq7GZ
mEG4mWMf13Va5ey2x12Oio+LYM9dPqRGPPX3EWCyw8FDrZlIlAPyRWq/Br4M8Pri
UEzc9zG1rnprMFB3nxkI6y+r1n0+QPmG4VEq8igSEvILv34LBQ1nEG7HwG8qNAwn
M+IDkvfvG/p1LwLTGG4Yva57VzQBHxqDuOjdo8wiacDYp4VI0p56zFUPRqWV7Fuy
xVhKthl5r2dZj0ynSvurX45Nge/o5oL8lZ4g2kw0iVbumFknq2mIYPhdAuk6CU+F
5iIfwTmYNiYKbIKc/el9CtIDIrVAzNB+Tj+I0eBCu7fx2UB1/dEsGsvYVFFrTlWO
QxUDZdH0lccm+FawTBfCesIWTWtyJr5hvNNcESPN7RFFXJc4MrLct+C77tATOYsY
AQGAW1PjK4Jw+PsbetqWLv+lVpDPapcbXqAUsTE6GKCDorFag8VLjrAtmNZoX/DY
Gco/nKNWMJ+DF1dBRKQ2ZTSc9u8DYCBE4B891VyzoDZNwKB9dhNziYN29FSBZyed
/2m/gbMmWQUG+cOXftwBtlMtmwqJylkwLAe1vDA5AEaDpu8s4pXYbFDNP4c4Ubf4
05oh4NfQfloy9KKBgXWSkjmiev8L46yMY6moIEocAkc1qKvQwRbRHZk5bEaJv+5b
t4hdVfMrrmRFEJAwlfi6u3jZ9GDgxjmxiFimEEkC46r8fMeEpPnuqPYs6FF7Frr1
4KOv+Md8dKXN3WW4TFK7mTYWibR/ereMWwrWhvWwTSHL+vJCUxvbm2E+cbmNQdKS
2lPEwSx7QNcSWLAPzxTjuaxfn/oi2L47GWc5OlZi3DJ78+SIJ1lgBzSkeIgvIqtM
/d9jMCa6tAqDf3NpKZxBKDDoBtPWLT4WrJfmHPpeq54lGJtRHzVwSezsxNe847ik
MR4eJ5p5wXpqOHNq6kjYNkrbeWkg1oG4Bz99p4WBW/Viqh08ZXDqjS0yCVYHa+Qg
SUW8jtKtyK7AUjKhjdR8xXnYChqw8Bqo6qd5Uvw8zD83zwMRSus/4hLwDmYblyO4
o1/0yB8gcgMnyDZxsGS69/WOVGdiO76YUzYlcMtWmid/3PgmhWS0QsUdCsIpAKOy
slNK1paqzCTGE9xNs0IiF3InWCxM22XmojKcpn2o4zp3k0AZOcDiZDNuD8w5LP8C
25D3lRLddyl+r8XO/uXrYunZ82+qphkY1xmqcGdl4BBsuSoGRaMMUgoeYnL8t+sL
6QJrW+SdRrBYV2GU45yAj6NnPqpFxpNxgg1nYoZGMgibunaXL/Jye+ymAXiGY3Y7
udzlCnvjILyvUuIF24s4XhoDRw1xWsVbh4yG56ymCiQwTsItqHYuO7lIyt/IJwRA
twpi3mWVviHypl3dl1oQegoRg83EsgwoH5W9z3wH22JnJpjHo3sctoP+3Vwkab9g
tjORyODSeyX6cEZQoKeNEgrJt8YmlY5DpEOHtK4bxVOqjGH18RO2pyQ0uP978W6s
TR1V4ljSNs4jyfOJFouEOZjYz71NBnrJpO8bb3webMvZzJhaPqC1TeOMVzpcbJc2
z1NshF63vWI4GHDpfejsSr4gPSeUST4UeyS9GyXNiGjkyUypFfmulqLh2axudE4k
SBieFjh2S+/8a9igoYyAaDpnWyX2ty2yvFMSFwyUsmsPeaRh1ZPNuSjnx3mRgbTF
1QbacwD2MO4GZzLDea1XDq9Yi6HqXmS4WyMmy0oVOEb8uTErC7IltKIwZkCRAjF+
66gkulN5/MOwaPJh0ud1AXfU99DlMpTr8Wj0+iIRCbDx4f3AaPwXitPUSp69M08N
JGygj2uS+n3VgSO17/XdnBv7+hOReJR0UgOH5pmqqVyEYyZGqSlC1C2MS69dAbCK
v4Q479w92fxEfyE8YS1d4SRGCPFpQhZIHelg8tD78dQNSUKO+aq1yhxGDeqgM21O
7WtAuabYb7ENntqm/IKDSS+oA1Dj3/rN1hIhcLx2TcG75WDjugR2luHn+T+JqU01
RDITgEbYXWRvgvThfr8zx9tVqdaj5XMJljEfUHJOivI50Gs8ku7A8LA/kpYYiiYZ
0DOoUN3vfn+gYl9ciiCyYNyTyVLN99mwmZL91StBM3PevD9zHhcwNi5o2N0Fz9Hi
8RfSw/mlN3LAPxWBHMPHc8FVNSXoA6sVIQk7Aalfw5w5iydbpFpxggCBmaqQbx5b
ZRXHCZtdMHaiuocvYS891ESZETPyspLk7WBu+CXpb/ZIwLRLq3QQDGAnu/lo0pSP
kdBUURgAsWMSUDydbRD5hL7ANYz5zQDDaz++rIU2lE+SAHc8ujNnYxtNBRpZky47
PYnoWsU3PWMlv+ufilPjASSeNa1efTk0TAanp+KEJJRCjxvk+SfFbE2AALjFjPOm
Ce53mqj6bUcqKq7gnAW1QL8pL9TGiENZ/iBVHA0FQ34fROSsqE8d0MCfnG4PDwat
TKYk560mtUqxOc6zxbTQEFB4xMKzAC4lLY+4En4jM21piZMGW3J9iSURMammUgr9
vpVdHoQhSNW+PpGMQjpBwLcOZE6QTwIhSt5EmfpwytjUcvOrHJfBbxc7ks8OTwcF
mQefS1aoEHLVGSBJMdxUOGXevL3D+V1QHOLXcJQdgzvX4Si1vfiOVLAFDUF2k9XR
ixmjYeNlvPLebmfAl/Z1/u4GpH9E+expjFnzRJAbzRMm79vEgol6M1f6CL3WNNL7
6f3De/SXhzxrF0gkDO3hNcs3RD7hk0rAR2DNTumnAJ5R7hgCvb0j68wRpX+HO0q2
jgqvddmVmsXOtE2wjk+QxI1dqpsA3XRCOjYZ2wduUuzJaDfueMoBLSh1MefF4tLm
GfXEsDAb9qfEu5kPits2/IkC16jYUebMFiMXnnB9oiuxV8X3ImOEFK2gpg6l6uvc
x/vxs5cBPzs/X2ElBp7Ej8D1bOHSuF8SSAguCwtF2oAqwxOVKekPOU/I59paAydT
Tww/3XgpuZm/Sqf0mD0XmiE9xFz8tzyb8lk05v3Luv64tMeDe2HAFh2Hh0F5z5Vz
jwcLoOOtDo/38WzQrg9fLpk7yZczJ7/M1b3BIUXIBiN8dntsvgDvBZ+WUpKIC04Q
rGZXG3GxyErObgZqLn56gsw7O1g/txouZH42L5lTBD2ugqrP2zQiivWpz+X90sj5
yvEhNQU3DSBdEKzydmkJzC6dHDj8QOXjAaMobYV+3oJnF9NzEERbpVnCDRa8Z8Tz
lygbgeKaA+Bi3g2dj3+/hm5oiJgi//87I6wm219TaviPoF/vKg9U4eQTYRIcZDZt
+3ZSk+aMVYQUdOQn3t3hz2G1LnqAZrRBAx12PvAu20sC0T2DdC1k1gtcyu1sNK7S
YfkF5tScEqEs4czU7j0ALGME9k7zjKw1A/6pMLH63wbgPZBrv3Kzh7T0dVmPpcPQ
YjSvbJBgKEVZPobX8JGiFTsBUBKm9jwLTwkk0ClQ6QEVfJrRURhBQJGouFAP4Ji5
NDsiuEKGDHodRhXhe5oMQ+eU9cYjeXK3lSbMvj+GjjaicACi+xABvRAmOh3N4+N8
gXm9F+Z+k59YMmsI2DNiYY99wLc5VRpqILJejfTZpVjP3VHxZb1ooRa/OLxUciAp
3Uc7DZmOb/AEHvvigmvmYgJG7VEeFyJiQ2ZNVuDbokNk5PXV1d7+JH3Npirq3KZW
VwTkRZ7pW/Ysyy3zJmucY8qUJyndcdbNhMKmbbMDUEB4rxJZL2jnPWIXDvYBn5Di
q9Z8/Qo8y4eVSH9X9PfpXgRpMP98oW7V9li2kuz2Wf8CFq3BfikJJc9QioACzZZt
q37oEuFGyruTad3mq/Q4W3N2FzyeeVE31kB8pKfwDqjq5Dzo3jHmaqVVZTjxqigx
8KK6kQcbiFsJKvqCcRK6ULYDvJN9SipGosM4vLa61CkwhCEZ7/JGfqaz/oCjz0rA
ZQW7n1yDZE90GoyOYd7By+nnVGRMU27LdY+lCYcIv3REuNILzJZN+hvlReOrXZCa
MWJpI5YskT+Pp6M8iXJLWlTwkos27uzmOa2JMigP9DQJuS/d6DslHOGO5vCRQNeN
9toQWbVlPPbRnySN6fAuiL8LPE17mPWIX+rS9vL5JuA62ggKnvL+3umGxnaoI2T2
9y0s4CzaKM1FsKq4XOKyy01+xRb3yn+3XJR1VtoB3NeYfFeAWGOcBeBLewNPYn+h
6QLGoR6I5yTl7wD44xuC9nmta/HJwnUs/kRrpd/i+9UlcUMooHF3qyLVNrCBKsg4
irVXCgC7CuiNIUxd0RzucihdIWdUf4qY1o5iImolUeQ1chkEmejpwQR8ZIiIBKLU
0xBErrNtQSmF21OMHrgVov5Uz5Bb/o+yw6LO8dkeLyF0KdyXyjmy3Rwmy5DyglFh
OvJpk4sUxdzA+4VU5BrttRvr3zT3eUHTuTMr1szjnDQjlY4msakmcfzFRFww9p4Y
fwdV1W/k4QZs1E2f20cRlD911t5bwRRZARwoX7nC+Q1pSz/xC96RS5+nDPer9v9I
etIr060ZHszaijQuRgnzqudQ5+awX9G1+aRAY+fSeMXdqOEvEYj5uAyZ/XJJDCNp
PntlOkkc0HvciN42yfppaTG1WAoGHOCb49nR6ytScF0UnON8tIO+ub6DVljjxsj8
GEu6ko28D3lYfFzWWgXiJNKbbrDSq1EOoclsCxUD32C/dVoPHC6xuVK2t5/TmOK8
c4opI+gKjWZHuUtKDt6Pj0dm0LL8pp0vmkQjmiadht4H5/jVeJMqOADVMGB7E6ou
XSCaCBzYAYP9ruct2WiMlYbpCttFhr6ZuYe2q9iISKNASRgxoUYVpGPF/VrDXVQn
6G4+rq2+n1PYyy2xSuVa3MvApOVFmS9GeHnv3F9jtXNXyjDkjfIMbqnm5hOFqyWM
ZlA9/xjKQ8r7LpN0Cw0XJOSl0RCPTEKMOSDw9Z3Zin0l40stW/G52V26WD6Wgjdq
o8s1pud8DmCHFLnMoU59rZ/abZ17tqkNuqSvLnCFP7j7NTEv4N6B07ahG4OnaDDb
yUB1ZUVaAR6jOtmooAZuObvbV5e8DoV34833cCSj2PgD+ZWWVyum2E3IB0QkY9p6
N8hKxD0GBfz2pXNx+mOSV3ZRNCZelfKbJ2k/ee5z1I8dPt9UfjDNNSySvFpQs7MQ
Oce/fn+E+Vlu35pr43k5m9t6mY60vG2kv39Q9QrqOsXbHqpifhL8XadiAcHZisch
GekGLSMK2sPp7iM/fn3MlurNcjIZ1nOaF8lOgpg7JKu05LoJ2F45jf9utLKwHmgq
adsMDHMyw9AKchSzFzVzhWrlMgDaMEarfhQQviAPCiXJmdTVXasTwwymc3pQDpwI
MU40nT2s6MptriiBoXcR/FzIKoLYb9dpqh1I01LT0T4m6rdX61Midv4iV8/OUb8T
YXbKvyBaMqglblLZ1UMcf7nuPIEDz7Af2geXPWGevnh4/HE+BOGug+hA4wZ82Wy4
/7XZORUYm4tU6IJRO5MiIF++r7l/zVMtPwnJx5lR0jVvVOsKW16fe4UXtzdM2ULD
hx0p2jpXxdLXjbvBTv7myqtZ5R4ZxFLIDjMXOpsCw68Z5aiRCvh9sBgTIQuHTaLP
tw6AW2GkRBhXw52r8UI7wz4BVSY7ciqr1v34TMCUVR9//iaDHe4QENBLWeC6cBMB
taTW8teE3+2ABDjjBmODkvt1tlG7KlnatK0UU17qdTl3PfdTHEBZDJS9FXAtbvPa
MGH/R+B7F9EyLpsYIBl83BsIlS+OH/UmRkgL7m03UvA+6hnD4u1QRNe6wlrAYgFh
KYX7HnzlQrMaas0JN1r9oB+erNpxVb1cJw7GdWGqoJoMDksoGTfRE0E9qDPb6uqC
eeWC+BjujU7dVQEb2oI2vysOHKqctAjZOuDRx7c0P/SFz0MPwVZkyDFCBQdIAUjB
OcH5WGvfa/x9zjNTQuP1gvoRQwjTnjZb/85VcOAx6RRMp1mSirwBs0ovy2eBpXJ8
VYfmOgmae4/y262hfVGVcsgCUlUdTYN0eYK3L83l6gzEu154R6VfXXThG4FvHnEb
B4yoUIBkQJTttWnzziHMDeVV2kaAHgpvrBbTU2W+1uwwUPRtpVQa+zLdih9HJZ2B
m+fAhkgdGL4U7/3ReSjh4Q6Hwob/KmtT1uiL7OtDKVVnkI6Z3VZ1QZ1AedJhwin5
n1b0GJAofSpF8f3acImP0qs37pIycm3bm7RasG1OOOQadluJyW6Q2pqeSOdfUzbr
xcnKhfvMFY5A/eguXxM5ed/FxjhpGiEkROKPBfpCtVE2Xi5sXj8zI1K9ukDK0p40
1iD0uvKIA+btogGyRpDVcfOQLoWp8p05ALOMydLuk6mIekfHRcAZtog5XWPXK2+H
7oJGzNKVCtoSe1ztpyubn3zuh+pYVZfVZshzELbA2itB7obzwu37GycLHxVDsihL
q3B73F0DGpIdEO4kM4oQxIFSS4Z0vojsqE6nwxj+lG+qZy0Qde/pqw66HSyQh6EN
1j+urslDMwLMBCy2Vn28CX8nOmZEnBSnLb3OyPvXTfdiaQA0qeIYifLDbzYFEqHf
MIGBwDyM5lHhH6ZkQ2MtwRUEIwCYn3ymS8QLS1YdYj5/Tyqz8SNCpfpZZSYPcp1o
r/mCq8QF1L9F8gH3OrCz2azHp2MN7d7Vmn4YaQF1IIuaKVd74YN1InXTj8zR6Fy/
WlUl1bLJFa8bJ+CkJb2JkU1Hc9zmCCOxydwiP2ErHG1rN9g2G2NXEtVsR+1/CKwo
xgXEyjTQOvwVVYcVz8tcz4CJH+BmUMf3N/4pzPAhLFfVuZ95Ka0H3blvFAwN8ai+
afZVlmc+gx9K9qjhI0R72ERBeLJ97rHr2zaNT/1NHGX5Mb/wu1ALfRrzHgSw1y5A
lMrSNcHNzk5DQ40Kb2AXGZ3QP6j/vrmER/P65OjFpWLfG1MJeoDjLuFLq5+PLSEx
t+kRaGTxMFM3JuKK399gGCLR+e5h3doGGgeeWaFvIM1/OldeMuvmSAw5S4rSJi42
t6zA+pz4iqlU8qBWf2K3lfWSZ83WXIErbop9fY+bfrlF+RP2gpRfiqDsQNXqrqKb
t/EzjmE3X8l9pl2OeONkhulaE5uf9mk2RcnhQxoGbnvcSKQRTUh04PgwDKP9SN1F
TmRHBn3p22XxT7LXol47gN0SZUnyMY4ApGht4ZaiBHeMisjRlHitqrH2+SbXQAFp
IlPxuPTYfOAgbbG58JSU2lWy+9UWKvjhUcXIy9zh2k6+lJOVghbogs96bEengmk5
B/WoYxO6dOXf9K3gmspRcPw3VksHJ7RTU0PISC8M1YeEKoG/mcH/yfn/r8oIGsyS
s53nJo4yFadOcgGcHrf2u/1ITVJWMlzVKazBuaDeTelO5jhGS2Wj7NA46eGzo9Eu
iBtEcL1/uVUepEeM/t3GgFMrJDgZzjJXXE5GBEr2mLVn5TPAf38XHr1rNqr5QaFC
AFOj88hceQUHlqycUCfwyQ1Fa+nluQDCv/AjX/kHWlORKJAbOVYSMPy7dXLoboMD
8NFWth6i53IYvdTq2wOTR/KmfMvyCSmDYwu9WlUeFDDhpirnTV49JtYmLb2oWaKh
F4Fx59uoa0hidxnt/2As06/mRA4JskLlzWyc+8KZCNgfzqa/Lwb1yyAG+Ol/vID6
tN6VCuzE55lw8453hsHrdUPEANu6Xcy0SXt93gq+30C1TYa5RpyEZao9HKB9IRjT
74/vkALwI2jp7wp0Jy66NcW/mlctwM2qQ+JV3CQZWSIGkjBcHuhBeb8Kqac7Kdal
Et4yWSsd4feO88RzUxU/eOZBQCqA0SxhO9IInm+YJM4CqqQffOHKvDeXh533w6pr
zs2+X428d/pJpw/AMpS0gnOsS89vDgT/v5cAVmyrAHEib8JrwSHZZ0ose8iom48v
l13D4ZgugmyqABiTszQYDHHNlX5texh7J7yk9NusCDI5sASzUr8DC3IZ/P0MLULC
vjDl6qtCliRnSl197MmjF2VFGs6s/5brCiZbkRl93dy2ELNF862KPctn+EU70+Ye
uAVJZFEZ4m6HFIfZnpAsdoRci4ArAtz/XZQNHx0382YWlLtQaz4/5O0W4056c6ga
cth/r9TppV8jRDJCnqoli3j8daCJe6/lVRR1oIB10K+77nLimch1AB7qCQ9n/XeJ
uxjOfh9iWV/Rlu19N/2jpj2Tdwj7iR7Lp+dcCgjlNoAzdtGHrTxhqhBd7WeB6z2j
sgryXlXKEa7Mbfut/9cRprDcwwvClZzzIhM9xLAkl1kJkjoYj7uoyfFdTaHmys4v
jY4O9RTaJkuyfTAZCjzU62/LLuePBPvJq5s9BcS+YLiAfg4LrlkH1pctpgQZ2Mvy
HOowQLPDGDihppAeLKSXwUY5U+3FOYPY2/G5NNCaqnFatj0wLPNN9LLNWcQ0NxJH
xauDlPKtZ2Lo1pQ+rTDmf9q2rBQzNXjKqop9/cJJQVkdmhEPqyOsSMZp0xdnE27G
lrGEDRpJA4fRbfIEc3w/ZBlGgCSNgZKwFlenC9aLQZ3NmVVNtUwTmlczpRCcM+rd
2DzVkYOOTozM8uYRdsUkdXLQUYu4YiJOG7aVdeIrDb9TSFZ+EEjPp5pqQUkXiYwq
Wk33fNguHjaVIbch5V586l5Ck9v19jXRFjDl7oZkLeyJokJuPY+Vs5ZrmpRUnmzp
ptPSXpSWSr5p7/hD048fsHuyPa+oYOZ9SC1lRHeoH1cdi5c4Z8oHU5IC4a1OvQOP
TT7KcyltmYLhnZoUimug5sSNs5iZMuXzUJrqswJ+p58PYwgiReXArovRrRLOsVFg
NDZQcqpwfI4ClZzS7L3xuKb1Yf2cgzqYi6aXpCM+Xvz8cp+pKhOYzHTH9SuAkhxq
jzSGFdRbWnyRMmQN+UDXLZHsFmPNhh3pf8+9y1uXkJ/9w1LjWVbbn5fXcrEBfNO9
wysQDk2Lml85nSAcYQZixIH6LCv0iP0XKz4kAFwTR/mWf1M8WtvCylW0xgM+WXKr
f4QX9e8NhWB0y8oIlAQ+w4R03NSDpPyEE1YEstgahhFcGhGI1kAxOlRWdqmyoXok
zjBHyLeBsZfun/BfC7G9wLsM0NXL1tDVe3q4aeCAbzODFB2mbGNnnQqHx+DnmUWv
LlR53DGVFYIinFevJrrA8bl7Fhx43R+3+BJAPEQDjEiOaL7+h6hCuAv4K5NrSweu
oZ9ziUr052s3G6UhIHczkfq4nXN6gWFDWsCgwJhx4eZTcAfZaTgQNVlnwVaK8AE/
2w57I3oTOn/OGeRIDUkczFbtwD3VanhOjzJMo5Iuus4E9aRtjlk5juyLA9bcyDrh
rAo4UqxGXUwW/zNk1iOc0lxm3jmCV0NjPqtSGzpxF6jGIZBICISDQd7Q3d/mdVuQ
XRhKNkmhSm030o2qPa1RX/4q1oJ6hm+jDFvG0Xvb/M98OvzHpOWPhctVjqjFCe9h
bNSL37nZ5XTyz+F+UZkjpByPKQWjLswXbChQOFOvqb3MK3L4zmojDjq7M76X8Xn8
0Ilu8EkA9rNIYOQcHekz5GNIMjPrUf4XSy/cqLHbZkV3bWZAkoX3rI/cy3zLaidI
pYe3YQaTl0c2htjJSfuc6rtugL52NV8OeAn+QyLbVhtGzekCtOyO5iMwil9t1mXP
llw8OBWXb+7gVsepDwdb+OecCl/k+m+DL1mIiiRyREJ6BkTJ1P7MhF9tlaQE74WK
2XlGFBXegum5B2iM0uO7ySGhZBBpi8StqJrbnnm790YtIxZGLCuSGySp/57Gjp8d
97sxoXw8NlxZmxfhqCMxEhz78/IOCAhUTzjvN983KSZdy1wkugeEOdmg7sws32FY
fze/Ne1iJgF1/MqjLvOt2MmRQB670Znx+Do80RXFowUiZFe74pVMYuKet2vDMxTS
HIIXY6pLXf0YvQyfMArDS4hPORdwNR0ojGZaRhV7epVOaKhRmgVLr0DKUWfJI+7q
w9Dj0z3G8XHg5JNM6mfIIwWih9wTjxHQ03aKOKoXi3zRmJRF/SgceHxVEdwQBqFb
AjmZd3Noa/QXLJb65n3vqSx/cTlruZN5vYKaXObqWDQd96oejBd46gOv2kYQYTQ1
nmAoJ+lAQgmeQ2w3pW+vgY1L90yf/oH7HjjQWVhbK6jsT9FF480z1m5HW6m7T2E4
5C1TfFOoY3u6pVsMxUOIoPyFlgWTuwKxaMtuoQVAJjDJuHMRZ/tbeYID68iu7HqZ
eNbp2wwa+MWzplRNs/Du/yjgnSwuyZ9UlPO6v0hc21BAeCK05/TAAlxL5LAp/p34
/skTbACzM+L/1GPf6eFtjaJf4CjdxfYwVkyCqAioJWCDNX1DVZEuLBchh/4rxSag
8cjjERUQtza+C7k8PZyqyrtQOsWi/EbvL55s3N1+2gAah2yhBJ7a67f21zneS/3g
ByZ8qWFqvrFdCK5qs3xrJOpcUlJR/MjCgYin6G3a0Gg3ep3ZczVym8EADBXE8yhx
chtNLDAD/wShWjE2cMwE4QYL9j2yH9/XbzLLH+MrLx5/3/et+wIXhjJ6QxPpDxdq
i/MOzpHZgYnIVCFq6JGQfyAm0eb2lVIRb6gja/sSH29VdjKzFAKhD/HXWRuw1kwd
MOwlUNziLbdF6RchO9RVCrig1xlGB0n1w/uaTzZbj/p8oRszgAbBYoITLHyaekls
27urqsxtEgzWlmlsE8laJHp5eQDalM1x+NOy/r8MqOUCnDZu5EgAnGvrtU+fSCgd
PGSoUvE1rzLqkIa6iEiJYTywJhuK9p2OptIc97b8T4k02VzHocMe7s7N5P9S1Zwp
4dY4bjR4KYIPKHjoGbrVwH3XukWUeQ/3ghv4HHLl2IvvrvOBn9kpV/j6fzcm5t0q
gF2YstCiLkvZP6806zR6GqIlfmQFEXuWaxq8ncnM/+IkbuZOAcamCcAcWZlIHaNY
RQXeek/+8/Rv90Sp0GfwEAOtYVhAQLc3eudeaPkOS7cDiLEiH1OWGS6JPq+Eq6aL
VW5/deVgKhqKUQjEBeoVXlU2bWEP1Yv1L1PeOrloLib0QfAq5NuUT+dodtfWEkQn
Y49jdsyVXVhMs823FZj/hGVJX6NbZbZovAkWlFGrZpuXjoPwNUZxNPi6EQ+H82Sw
64ZKHwXmBt/y3qtoOkuIWeWK6pnu8oGiY3cQGoA716OpFFj1FvUE7vFCs9GWYoNf
li1ip1NJJK4rNC5jTDZQ9BGdfVEZcbd+fcnOizbLaX1Dyv9JES8CXH84xk4Etx35
3srN0Lkg1OAPu6eYb9NNcPB1PIIqlHmOVKZ7LZv0SfNvCkzIw0stPQ1yxTKhbjmP
z8MWinMRR00oyK/zjZkasVuGe7J9OfU3v+rXqTx5QWac1OQy0jrozGky7/HVj1EJ
mdKaHrbQA+96e09H+XjtjKFnK2wW9d7f0fR61GBXoDiSoP8ybipoZVQSrdTefBGI
zN2ARlnZvnKtB+59455cpFJXbXUH15Pt1BTA94Bp/WUdMD0vqQzbKbyoF0YujKcG
TBUd9BcotE/qSf6byBE9N2aJq9KHzq5ilhd810qnnEptnP88g4fTgfcFleKrr2Ij
py5OsFJ/93CFEIYkyQOuO5KOnT9TSP0wgSrXqKSeUoJw//ZLXKidpk3F5RzjIVfc
ac3fGK9IBj6MrvaT2Z1u+WDaPrhXnIJIm71A6ka9Ifq0EgvEFFohGM5VMCpKA95H
N5THHq9OtYrU2EodUK51dC5mIUETgtPADt9GhiwwzNCLvrDt0vWQg2ibUpAEhZRb
sZOJHqXc2TE4/tXS5qZpqst6fHAaC50bvZ8L6Xb5MzaiGAmVOLaYhQI3u4CUHbg+
loP/OfTg6DubXlQ6jRNS9h4t/RffAGgEC3cvZUPON9dmgGVqhA3amZy0cSz3j0Pd
e1mZstZpvK5G8DfrET2VdbEq0AXcvHK/+V17rfhr/VVD+RaYzVIZgxuWwqGZO7am
Fvs9r9/+eFIg6UJG916pb4HiFLycaVYm9nJ0CSr6eHb+KZC2QIkRFvO/Hn/K/KCI
lFREr2PjrEp1315/xz6KWe2mY72JS1j0tRQIUjh3GK3NxzIvid2U7Zb2RBe5r567
DNsqBwsInHbnVir0TARKTjH8QsrPxYrEqVDfvTslPGFLNbKvpJRe/9JCbwcKTGS5
E4CR96o/2M7BXVedyEjz9SzdQ51iDcDEcumYcWzVzXbfthmmX/7ecQYZaNVVhsmW
HgRZ+eRkzCGXiuxWgc7UPg==
`pragma protect end_protected
