// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jBcwkswTcTHV5FcC9q9OU4gH+9FqufbFTJmC4+xs9FcHFwokmdkGSq5FhX8NBlRV
aNun7IGOz4TEdclCSabc+q7dZAeKHIjKV/bZkH+8HqwFteAogWF0LFAQCgAdNeDl
7ceKL2cb5C5exoB+2y1kJ6/KTV0CBRsorQaio5y0+2o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32976)
f08Z9Qt1Qua/X0lqeJF6pdjui6yrl2DGhLH9z0LZcu0ataHuh3u5x2VSzVOToCAd
elpVtOoXyjZjIU+wzcAPoXWoziJay8rDi+FWt01uF10Dc2WBHR1VX12R2xJoIYGD
kqfUD00HwOrqfI/ER6dKRMs8ydh7eVQCG08qylx38PnDA8YOOllMJ3ULH6NzoOaQ
wd3YfZisgftL5sftAiMctusOtN/qvL3EarVK22L/4L+q0hc9ybwjbQ8ukeIWuYSi
tDP5au1pSy6sXvUvESCv+X7uOi6MyS96LAgGTiE6pxXZpQwH5JsbnC/geEwqWpV5
YJp6NrKGtE0MxREHk5RDlGLzUcRAxCwbzuUF5S1oENBIElKKfALhJmngRed8tdTF
vxibjaJrjzDAe0x23HXcReQNFvLuqFBHSSywAnyZihVTuQn+mlKFrGTOJBNSAiWU
/xPY7yNcLqQ2srpLkSuNGvcXQvCEJG9avrTXyhremOBsf6I2J3wHCvSsjLlvdxAs
wrmKYYohnEoGN/EfFMy2LqSZynN9c3zEryxhZapUOIiyK3Oqrt9N1MwjA+NLWfSd
4HrutIglLUFer5X2FWQn+yhyyG+G3IAVcXBammWy8SqszRnyuXBAQKeE/BPIBmyN
c7Xq3IccXHQZ/yGHEILvLiHffhkdfT2p2SqwVV0ayvUZUYhupcwu59ScjNeJxTib
cRX2CxMz5Jq0jW3qrF9rBgoM2dtqMdy2Gz+AUpWXG8BNz71X3Nico3lH2tMYAJkj
PReOuyZwd/FiWpaSwK2e4XMJXKfyosMpZGrpxQd4EpPWHLULxVPmNu4hDKn+nk70
/Ng8FaQsp0a5Lk/4NJ0Wf6+bYpZAO/a7ZPNU0dGIdEHqPm0yyfvzq5k3QRFDcAFE
Zt/28q+fYe7FrrOUmUgGgBikbCiHV9OwGvbXNnz5HvfLO3Y6f0ywJkjaEmogZfzo
uGoG3whQHzOwgm6Ws0wBkJ4JpYyNXzxFPd9JCT/CL8jM5It8+OSsQie8LJUtDSIK
Qxut5RxF7MBv9+fp8VPMJ2Wrltq2D/QDjSPuRn4jx6HP/4LvJmkNUM8Z8wFk1qgL
fzEQHKj38tGlqerdodlxj/AQXweB71E0xv+4c97jwyiPBLSV6R2DRoATbuMVsuWU
3DwDjYd1cKRZ9N4amj8u68e8P/M500xZSVrwwm6rmuMf8+4Zzv6hvNur8Q8Y9ar7
IKTk+YjyQ78lkRw6ec5uYs1CB/6/5u2KtL7taU06sfq4f1iXUTZl860jfl9ylWmr
VnWeeIQd/NYG+iQ18CcSmu0h5TnNC4XIgAS3Z3Q2e+NV/BDAsXTk4ZC+tUS51EDW
ncqsTrUUiaRZb08WrTSxG8saoeoZdlUKl5byOe/OgzVMSGvtVyUChto+H6o/nmRk
D19GXDeizZyNSLDY/XBJ3lsCVfb1uNTwc5U/dkOo8btHHkQhYM0TRJER9R1O+J9V
PVd0ybuS83d1jlJtOm9SwQPUkgsSHZWFRV4qsP7G8OnETs2fHD5FEeafS2af6oDt
zvnSTO06dazql9EM90oLsC/QFvZ7FAbcBvV8iH9xDb6ydYuHCqlGI4zCaIO8NRr2
y694oxJmsMj02XIlkzUXSzSxnqgMCYCa85MvVoz/lMAAh5EOCoQhBZ3pPghahPKY
nTm0tHTsHEalDudlveBfKQBGTZMpcIBFQl4VFRQ6LiIlwIOtxzISEt1Wbwb2IS10
dXNLygiPJY1Od2RJrRjIcmSUtF1wbetp/0f/cMOxgSa+kw63VODBNhi9vhOEamRY
wSjYkfLcKxGa2SuLroX/FaKSY+j5e9pFoQv8qBAVs73NK9Q9Mlp0dXmbdibp4Z/o
FQbAOghmMc39EY4cbhWPBsiym5bXewvkmyzBnEgMndXIRfZdi3CHoau4yT3p5Rna
U58qie01T1wdx2ECaWbb8r5aUi476rmc9AFDrrnuvMXunH63Pcfz4RojIIF/q1Tj
0n8p6Xj7If15gxIUH9goKOZ8iaGg+a2n7SoIRj16PH8+gWK1XTBmePo3H1J9wNi+
028U+SZX7aJh675ggvvNL7NjuQkXGZk2OqeoDI0vpBKMFBzaX+fgqVnCLg1/JMkD
0Fiv6Be58MBQpW7rpQXH7GC+H6vFHFCZEA4f0T80Hv48H5RwffIAJrvtfz4/WnV3
a5H1ZeS6oORWTzlzhwVYPfZQacONKte7dBn+SJstV2Mc83kE2bhe4WU+lClSi1R5
53xAfuRN72yP3S97uJGL7VeaJgj6VY2g0cU/MRzK4iRb+YHiLAMUdp7CKTy9wsvn
aktBx3jv6E9HV0OV7R0SBOr1cOQyflfShY/BorUJvAWS1lJT3wrxrNZZLHbw9kE0
LVdP1/ZdUJjSxrYc0VaWswc3YhSLkfxJeSTmX8EYDe3xsSyvJH99qgwAnRMVeywI
SkEBWjWozKFwckZjsF7MML3IUQx5BneyGNvz0+GUwMXCWXPA0xT5uUeTqddb+4Z0
lOhnEycvfq6fuRfE4+jcxo0cmQt7Y+vZJhiGrlXFDT9+KdkxjqVOAMRp2q3JncVa
lvwD5U2TpzFtUJ/U0j6UYr4m4Gy4HrtKZnSF5gn3fCrm8rWj8KGj9HE84o0nXiz5
vcNS1eZVb/Qc8OR9RlWR/EuOxCN/VAa5YTkFH4HOUumKubW0lv8Q04JCTX9Bv7ip
fku1Z4WA3YLQzsgRLZNYXb+WcfMwqKTbpDSyvUnS0OCRtgE2ulYmoMtAsf4Cjixo
Lor/iFoEC0h1gnnFl9SE++rp3Hg4fqX2Zg26NNhV5PszgVVNXDZRKV2mVvDEGXrv
AconKr6KSjf3lkXycd3DUf714FfWczsblNr4KTRF2vUgqPebC+WmpEqbvQVZfmDv
nxJ5I7tIP3GNKzC8Ovq34VtD3th/1EedEI1SFgrHNeXHFVHwOnlABtvLszKZBkQ2
sock1Qs5w0cAHIE8zIN52LxKi8V2jkT6HQbpXLC7noR5CMLbEWdFvpKjNSJfcHo+
BdIJFs67Ie9ouj4Nb7vwNdttMFJ6WrHiFw+binzVyMj1O+EfZ1tNy9A8J6EFQgHC
oQDKYINnaAdxYmbvX9/4yLB/+wvqQQrQ5I4XBBxhGTAqK2W7s/9qgelj5k00hnrC
TRAAvXmOrQu1UBtxKFObHpf+Cs+kawJH96bgflJsKUVq5RB1VAWTEllSfOzpdn+Z
rGdcoyyOksLhFzdrjY6HC80nI/J1qbmAJy6Xar2/pSpQyIyElSje6bEsl1tSN3mm
6tLBdpuQF/dV+1i/S31wZsBwix+h86fNCjeHeA8skFsD8QkQshOGcMm96g8ARC2/
D+284trBImb622Are3NISWLn5fUbVWNDSfHf4u65ZEzM3bvEZgTspMKS/4FTV2N/
gdSmz1W+jekVa2c8mX9tF+/myESVaMnLHjLmD+4OPrjWMgrrQj2qto08X8TV1mR2
YigedjiV9D3uxs59K3GzMz4uDnisqSYhfdiGJezuLx0L6NpoZARfckFeC2p+WXHn
My4eAvBdYoWUU2cYfymYFcfMwi/XjmlySDKhbnJNQ43KMM/iNPaVSkwtuHq+cUxi
fWF3EoLXMMZlR9r2l9KKHTvNAUlXBAo4XiEWZqc0ootbLBOcqAN6iZNdh0f7Gb6S
cCUhNK7sjYRIaclc9bJMCtn3mBVMye9OVrpBchzqdq/2F96TKZecHwbnwCG0nsHM
8lRj+vpvfbEQzYkD63zpIa1nBk0ZUOxIew5lCw+qGndDXQc+R4pF3zxxNd/N952I
VvmDpDoXz4eQw1bP62/Q3O39Ui4VbXY5t+y0kqW/lorLZ7GD/7GaMN9GD6Wvl51J
Yb5oY6lZ4aRJonDN55qCLh3I/d81omtdzB3fAeVGQYhKYC0BGIo3U2uCpDhtlgAg
YjQDIfdPZL8nAyN9/lrCm6wGhmUR2lDfdi46rH8QI2uguuqAXRQ8EuWY01PsfZr3
n0kTdc4QABZauWJDsOsp3vUeuDzLEMEqVLIU68ACAHOOfZp96SLjecEK9rECCoQE
ISpiov/g0P4nVSvVCT/jPN79XqEQytmXsBAj2/CpQuk4NDiC+gsnWmPpTwTuDuej
2y6ROVSfLS34IG/wqmc1ct0DVvUoEKMgc6B47s8UUv6ikQ5bXJfmBkxiczY8AWlz
3uJPDpFjzFnBSlKVaJV87VmAPeBytMR0o+jUpBLv7KPTlN7V2+HvYujAgnEvIFMk
ZRub7OKlO3ySJp0DN/g+SZBsdarNPWRYVVaLmwb9nqaxOCthBOat63yA5LZyRy7D
MFxk2D58hwp4U34t2ZrqlgIRiAi0EswFDjN6699BY9DWmQsKLJulfotNQAik/aVM
GFou8hthKlwjt6HuTgQK1FgctRLy68As5zKhtmwLgYCtKhJQX4FYldpgaDosadpN
AH8l9tNk3tanKp92oxhWc8G0/QvZ0mv6tnasdR3ioEOqxfczaTcYSDL8lQ2n7mBu
Nogp0ktwj3YNmYXYKy5wq708ugu8JRhxGTKzfxtn3m5RrcOCaXnPjP4LuYPaG73z
TlMPrdjKC2d37NhqmCA/+Rxf7wNjHwf8l7pjMK1DEpFT2Jd3NBqFDK1cHHyQqW4y
MSiA55MHdpOsqrCImIx+5zlMiMKvqvQUOzas6frhalmQLQl4OJbcPI+ixAB+BF0j
FIOr6ZeOpb1zfUf46V204EQlwJTMs667AKi82Q6fneqPOrNrTN94F0TcO5vWfxel
T0enQk+gHMfRQEH4wGAAIIcOeL5G8B7cvBoT2jPa3I+a3PeLm193XKb5ceSZeICT
HESQj5/xO5ufn0NGgDliZQ1qe9c6r9sSJpJBMuawtIcpRrFBwjlTbrH3UivCQQon
woE4IpdmwbLVjVJrXsrtVPflutJqlxYAVLHGDLqyw6n2lZlY6CVr2Uv3MulFKGN2
FMjHggCePRRyGXgzWVxsNzXGfusFV88RuBc1J2eY/J7DDwbC2BCcQjBDODa4kWuS
x4koVb121fhYiB6DAdbjCOQ69p4PTpYWL7gBnCUmb28zZX07R6xcKqMZFX06CRPF
PBehEfrRpuZ21iVz7FyeNygh4DE5svwvF3B45cTJA6vksMY//ZbEzLejZ1k2GCv7
2iUMGnpEm6vsvdTNWgLcA8yp6Bz2DtdSJqanykPmaBI1uc8FZLvY41tZFWu5yPwz
0tEDBzyeL+NVMXslVULMfJKWVASJCx6WAK2qNWQ/Hgj7r5fHJ4PEwxGid94GPK45
d0ryC3RkC9zGO60Waxuwb9J75f5z4laX2W+w7jdVomMCVJV78WJVJ/7O8Z4FqUGC
/ceDtc32Y/IntwOB3/o18YlahhBbCFC5G3hvC8LCYD+kmuAHdAarUF88b/DXfz8r
svBbNYjNJHvmIuHvTeaI3h3MdGgKmulpAOAYvRvjY1bPSZb5DDcgHqmMrxTZlih6
n2vwmDKso1KG1J9NTSZBE7BGhcx7h06wNkQFsdELAuTdYlVzA3SBJbRUYmiCGZdO
xBfxKbCs5W0a1AhLN10ClPPj6gVBwVOkn4R0q5McQhDWSmxV0ZW7mEKuQB7BBROR
UKobMZGeRc7hc8IkkJMQ3ytigLADos20YaEIq+0AXOjrycna7+FffQMPPGjkdqVT
3DVTMYMRJJIdb/YnS6xHYrGjpmni7qwS/7lG3Mg22p6RHNmByigGnOtkvaOj5AUw
cpuZYAp08v/Cegqj578/1hqbMsrWzXZELuVpOTauylj4mZ1qAofuTkfsFv/PYBy3
z2kI7QGwnMFsTFjiAG2pYyhR6SH6uB9tq2LHq6VV01LkI3wPGz34mChEfJ+0OmsI
/OMWzOJHOXZSeQVED0b+3Ef4+dZHsVeb/KhnyAQ3LEdchoL5HMtmTKHqjNLuS6A7
aK+4iNBbTPf7u6v+sBe+TzjNgLthhrfGVOd4Qs/QxABGaACHAfZrtxbnwz+qXeO6
kUx8Ur63xThuPHjQXjtlBn6W9YafvX3yfTXxP/UQvyiIWjprqJ11b5kLcL2DNg0S
cKmsmnHPBfmyd1Lhca7+ydoR7edXcM7PocENkjBVNO19Bbua6mrKbH6A4s3FpMxB
JYt3dkjOC4+9owSxC/GzkFCoyHSkW99AtqJeOX3Q6giQWld8DE0K/y7/ylaVU3q9
Gg8BEQDGso921tRekt8cu1P+9szukF8VENqwivCWl1cmpc0DBfe5ORU+Hpfbx6oS
Srr/5NH+Mk4J5OpYEVozHWYV1Iebo62myJRr6n4cH2+tDx2kNjiLYZj4xhx8bfpF
F/mE8QO3NkghG9BCYEpA7QACITvxWiOhzgG/KhuA9RVv83+0ABHELzAIfpcfnxv3
uk9K/O+kdVH4MMrdko8Kay90ahUF6MFcRwWF3HTBM4wv/ppArxF23MgeGq1X5tDB
e0UdhJi7pdDh/tuMfHezy7vs4STEW0dCVUs1Gwlg6LvzltIjnmWRSqqYHU/yJ/u1
07f2AphkGhwZgSBCVCFPc4OTAEEUO1Jwe6Ua/P25OtrkTl9QXHWXaEqJ6P9nR6+x
FlYqLyG9T1JtcW6m2ac0SdmLrfIkEZcky//J0wr/7b4Y6fNH4+8i19FSFfF7nSoE
9XgDiRrNpKukYKCSIzXI+h+ic05bVHBedLNxSnrFWuTdcQJkg7M/5FwF6fE5xUTF
nifGZfxy9XdFKsZcgWmAyGkai/ANS8CljDxUMYohfTanScSUhjE3VCeARJpM4EOS
tGTP4CGMTZ7jxHI0e5IA7MPgjg3vAe/AjPsw6OPSYdbH/PJH2w4hi4ibta/IUH1G
LPPOpM/WEDeuQzc+Uwv1uyRQOeosKEcaVBvNKMfHAGHFSyQHL9zPf84no6M0DtDr
bpLtdDfm7A+LYOJapRATcqtMSZx97g8h/NdoACQFrMtkLek0D0ZoAhBiL4c3r7+3
2r3IerOFz16CLf9Q7HG9SKimGjv7/zY8xSMgwp2V8pK87pQEooJk347PWd91Q3CJ
0Mtfopxj54HLutdEpsA1Hndoses58dOceBb89uu8BLlaLlHfds15JYrwtdvE6e+d
dpP7gRmJhJmFouCVJr3PbAQoxszbfQOtlaqR6gJVAZ8p3hh9NwkD19a4dOJUHHLQ
KHyLwTLiOQMdzuiJIPNORswjyPBvxloRmWqd9EBd5Wm4ntSDxOOxMjKG6LBD+O/X
W21jW6TNbbzTwGxf0OZdhBCK4P/sqyipD7XrQie2UZdN7+ru+3FkBkitWh95U6fm
NNNX/q1Se+eroU2YldzOb7B3+35tFkI7H6cueIFft/5HYziq++kBoqI7TmZtEPSz
oeYMW9WmgqSMDpX5Wojq14Xgomctm107evbaJ3EdM1SqSaeWAgAd6xvV9NBssYso
cDOpmuem60YmJIIwbwiz0s4/GEc6vDPfUg5VZNtChAsadlyYEZh738uqHodiqWJ1
0t8qZx7l5cnsfASen2IAdtq/ENCy7dv5V43jIwqVZmA6b7oxDF0ZlgE4tMDPzDUR
QUvV2eurppslGvwo4NpKIOwg4gXmGyOYZoUtmPExWo20nxWjdcxoeVAUPECrhdN6
xF0h5JVOTK6e9WlVnLE7ru1Y6Kg2RRnyL4tiUurFs26r3DpA3CfMdEvZE4539Zb2
xDfzNPiCW/SezFuNfsoQMYeD3KuGKSAS9UrGxEFav9CuH7D/X7lOs2D+ZjRueT73
X7IZsyqHIsGCgXcRMb/RP2JRl3Rohf7T3VFo4bXI4zHitWzizqWhwqpgevGqQU8m
74wu/ivOLaQzueX1GkNJYAHAHArxVLmGqZN+IWPWPkU4urCtpwu+YXLDk2RXEccz
2eW4fH9id+Xc/u1ZzJlXAuVTdVEeGwuBZHwl89aU4I1+W6626az/nGZVzNXG2qXR
MnRnlMj4L4ZxaFnRN+IEZYDZTyEGQawaHnI5hgqMpLaSFY6GT0zZbkbGMl36xulE
u8JtCAo9YJxFnqC1GrKIS3ktP6vgJrmhJst8N28mTTrWGVk9dS7eMYpx+QvKjnqi
yCLesBHLE3EIAAqk9SoDEO/CjOviWn3/3WaAVIRb4/Ll+jS1iA5IauZ8C4CtN+8H
e54XhMQaLSIbZpPFpmheUOvzril0yWrHG1h9WZWREPSbvxuygMjECiEL2hrHnY6B
hSflW7La26lpFnMRsUV7XOg6ccbRYv3YzTm25vl7TMSRdVIuov2zaqsP/gq+dagp
QWElUNikVaum4vQQFwp6DDTowE2Of7ruBhAJcGrX6h7OAv6RJB3d9dCexJ7iPSw7
nr1hxhDIqeBFN1BAypgNHeZBg47bSgXQD/KA+0t9eKsM+w+US/p+v+rtMPqsA7sl
85ETDXHniI8i3kMtKEZxlDEN9hBFrHkUPft73cJ9YIrdhLxyjXz4ct0hgxhcnPwO
DI/vimC5w4zY6PaQLgast3jd7Ou+m2vkTz7aaJx8ocQUA2p2ZRLs23miy4VB0RyS
NlQ1+UsMRbsbXXp+IvZS0Nq9bSf3oySz+p+H8fmc0fHRgVD3PCDKTUFq9wYoD2yw
Y5t09Pjp52yf3WVwfUPhNsMxvys90PXpR0Zqv5HkyOkE0T+I3G012LuLw2Zx//XY
4ODwW6N+cbAZEBIv7NCU5wbXRd18NMSohHA0sxfdEFQfKkAGhkjmJxO0TQ94qZ+8
IzDwT8Z5MdArYQSnNzrMBlljn8OBslrMJoZO6ahPV4/tmXM5M+9IQ328aQgQzCe6
koXrBDyFStizh0W3Xe/a3kB+ryPq0vT1924a6g3IdeKK/DET0xbyJ+dgDaGNOUZi
v0hz0o6BNn2vWpKpN+9qGVPvN3YAmiYyxjomynU+Hcf+gEEQSSXj/j3HhYSodbKa
hzrnBSdnJT1jL0bO4QdU0QNhbOdY5LPuPT+1RAt7P0IAHA4+ffxhoh1FYeCrQc8M
cAZ26clKSS8p+ty8h4/5NaU6CHfVklTp69XdVZGShnRb64X33vT91Q6/WFX6WCX7
Qgnvk0KFSROxOf1Q6gxQ9l41MA93kNCPhSwf5MH1BNhK3lcC6xariTd+DQOsj0Os
vSdzaXovw/qmRO0rphWoFyU+oYZZiG+FI0/8SX8AR6+qa1r8exRNua1n47kik5NM
Ig0W3S1cxcwbpy6lpST18R83Afop9D/VLVH1JdJ9E6VClysYFVCLRGrwxKCXfyqH
o2KLQppAK4Btlv70EAB+IL35eL9vRdfPQHIa+ZAwFDsSyYgOnbALRs9kMxqpgAEi
1BrJ47Q93OQ5Y0VmGDhkrdKSqVSMGxuznGzM3pTlBNOXvJmbT37CPRh/Kx2jUffu
TyesG6S4b4lrYq0TlSN7CJTG8wUBdkf1QMDjZEccXh21/fe6LPJuVbW2sGTwX004
O6/9LF3xRZOoYQ2/cyDS3pA34nuayD4WtOw8IkAf3co8T9AUsuNpQkKT42HCutCS
Qwx4l8O4lhi/b+JfJrwfhkZsRn45Omxt6oYTELSbFWbOWzOgdxpNRQusazh3tNd1
V+rLgFeyC717fRvTmOarv4nhbPtAS0fETHD1lAb65rcsivqgLLZGl476gprGyrZN
9imxM/qfN7iR3nSa29G6cq/ZWwfLqmAV85npU/MKWxcRcFAdM4LJxlKOe02kw8hJ
D0jpxgCqWu6MjGTwmGvL9jvKZv4G6pF6ndEghQ92S7cjnWoWjyqfadNIGbl+gQHr
hz3Q1Y4RS2ZrFliBW0cCCxFMPpVLrZKnAarFSYt/5IGX6j0OLWkgp7HJgTq9EDeb
J76x0+6Ot3KmlVHe2vnfPT9FQrVNEMLVLzSwTYSWte9mTtBJyqb9pm8kjiuBER5L
Xz+TPzsTsoAuWs021GA6/U2LAgZbfsSYrYPa8PiJ9w3BOfhpigtOx+VR249LqRXv
JWIEfhIqhU37PE2J5jZA/Uim2yVVbzaBQGpxF9+4aVptM2AUzTSq0ISfASkQX7F4
5OeyiRoeHAnfrHmvX0GPrVNgqKFqR9vg7v6mmBZAO81WCxG9yz+5tg7ATazz2IaG
3QjXlerXG11jd+6GA28PFerYx9fD+pX13+6gdNb2UkU6OS4rGVOmQjB44LF4rj3E
i/U9E9+WqNgrQ8dywPTpOIMrw0XCzAfDiHuZJUFdPrLMvNap9ONuf3FXyzWdDcba
0Tuz6RKF0g3UOHbYl7cy8VkG6eeht7M97aukbNcRA84VL5x+qQREQsi2LWzCXsXc
jt0ifITVjJAgDQr6fN+PRR8xTM5N8lOBZT3gUsSNK2j02bQOfghwc/q5+iPyqRiF
F3Qtt3Xck5TntbGBv/RrFKHLUQHK5El/7ofhK1rByiz/elVqW4Ua2f57s9BI0WBp
slZ2A7XxwqUKB/71Ti0eG9Q8bfiORcdAohXxbfN8azVRIyZCSQD+g03qAmN+jdZX
qarZv6RNsWVWkryn1vrABuFk/ai3jW1daZpt+Z+Y9HLc1qIFoMzmOZL9MdBHgh6s
4tySInKG7FCVgcAHwPYDOT6FHfDdreQef5ceD899wvfhJQDRTr0g1LZ6PMoOkMG5
koqNnLVrzRxIFMCyDAQt77WZ/nh7cx3DKotqsWQq1OPD+c2x0EjM27i2ZoGBHEoB
a6WeOiO2kHCm3O8fcKm5i5KnAlGFvz5fw5OJ2YHD7umC2BMgwod7+7sYJbjYZLfl
gaFwSjxF8ZXds6MYDhozGR6neEsnfxgHhboRqM3O3oyKWb1cdvHfv0LTtIs2Y/bd
RrnrlC1+WmjncdWfik3b+cxpa0vA866+xhzfafWV5M1b3Gw1wiRYYsDOTcAGgXhq
KcJWaQG6CqDmwapa0rMAEP+k/SOa03lD0ZC4xTbONuKAt6GxG0xl+eqgHjPz/CPY
MKQ7IKCgLMqlGYzt7ZZDBCOv8qn0JdSz3m1ZBABheDac5lKVLpIhYFW98k597GZ3
EQ2M5wB5oZQGcDY8fSgvVuWa3O4pAkN4i+4j9ia1N7Le+GcE5izNPu3QLMAGGL/g
9VgqV8jyA3Rj3L4E0dgBbz6EAipr0v/mffmOD5kToIq4G/t9ZLXxQ7LG6J8Y4q/O
vGjQvlNI8sRjubcvnYbTE4d82aARBR4a41g0C00Ry71XSAYlRNQlvIxw60FVMUHs
t8nX7QCs2leNXP2z6nbXGO7Oe9a+CtE/HnPJxvmHhKAmM2kCpr+TxsMOYLivWwOU
IR+XxqP7588LoIeRDz1XFHpeZDLYFgpCg4d04be8h4WeRsZ6hKnIU8IQ8oqPgZ3q
kuaZmGUtCYuZh//OHyJl05/X7Amy7sF7VH//W/KRZo6nzR63jlSYN45EzG4P+DXi
qXAJJYeX4R3iv/9QqqGnV2bK+rdqS7yJ9uo2sMchDSIxxQnDTRtpG72hK/JBd7sw
/8Pz6mgS3nVgqBaxkFChcYyDQcMmz1/NTtfLSBEZfPGBYGGI8BRX+dX95YzcPxlO
VSOpkps9QEwGSktm4h2GvWKj6FMaCY1rglOp1/y1f0D1BW4muy8k/fS0YfUWKv0/
c9i3y5YL2WV7qEHTIBwCk1NyNhcvarOA5utvfkPQ2D4+ngnX5KaY1CRRWjokJo+0
3o7ZaNeOJYTzuUjdFPTdIt0QtNGUmYXkTsfsVZAhnJwDGXVkpufLGCrS2/Jrn3Jh
AqDI1tTgMQjL2uDvL/IKf5mFWeMxXVQVEswGB6Lgq3EdX2/psZZj/+uv1pXL/UST
Z/vJesaht6rxL58SXwysrRtOr4uV9wyKvjIOMQGk2LcE9cHmUKlao1pWV/hguaXZ
oNB0LHXn8BDZ4zqem81EfIo648Qlj6+Fep9keFClieBP0a4Gs6FdjzYHs4bVhaJ1
M0yIcmiaDhcXqt18GFyq6KT1+NICWhNIh3v0gZiUSiL0P7evgIx7YrARkiJ6JMv2
X7kXhhsv0XH0S0PlQFJc7PfxL6erOLM+ib6RV/OLoYV3TFWzhs8ejq1ugQsyTDcy
md1bo6BOzCqeo5s5q1puup6YwbM5d2VnbUwVfCb3Lf5uf3LRwP6gtiarlMbaPBMq
i8fcmNtR8XeStYuQJAC3osmj9+BR2y5BN4M2i1F4rdltrA1fKwaLn8htnTn4mm8K
cGmrDKWaMQz6fkK5+EerzxDtjOlog7x57nmOnJULiFfWtJ38V+Q9T0ar0njQa4A7
xysea0ruIlFZmf3GTgMf2Iq/JcaLBxBUorfIHKR5W4d+OiNMhUiRiTvMsSTFIJrz
9pb4Op1ir3Bzahto2TFgzSr7gI9KHalbmeCmyrs5DFGJI6G3zfAwTLpQ8fMRzD7I
l/G0ja7tZq76EaDyPHW6oUWwUxXms+aoeFS0ZuP7VCECq3ukpaesogYXRuAtqaVA
B7doi5pjGQLmWNYYB6VRbGezWxkhhxOGB6Vc146rPjefJF/Tel8ySwdatwVtniqu
PwapyGnDnAIKua5urs/WqIiosAnOLeexLJCyRRbevP7eI6NB3ARjbBpKKZKEHoKc
e5vN+UW7OieCyi50ThMkDq/GxD02tbUWhLBIwf+DlzHoONDva0U6sKbY18nBeFtB
MJSLDcEdO8IXCh/C37n6VT8KU/DdRERYa5OuIPPjGR8UY8RhKrarT1MZDFVvMq+b
YMSouNLErM0hya08ZyElBuHqPJPhtZ2m3We6Fn5gGvdluNeGGt5x/ZpwxMTxopnQ
th/ryuPgVZXoxfoAuk5pfAzyRADc4vQPS7/3WKRf4Z5OA2JxZfCEFzbsnv8zfhSi
pCRCY+vCwUv1+sqxzxcjWg5EkcAALrdAdYDXB13fBZ+2dHMrkgeyYL+6R48y2TTa
LWFJmiABCwmmViXol3jAXABRWLNj25Cx/bBJmdSCEiRg6yNTYFX7Eaif/RlmBrCB
VvENUVwoXKdSzZolgb/yJYpFMRqlQaCdqoAUTDSDHmMweNxEh4wBwd1d9T7fI2Rc
P68mk3gCIxs5YI9yf0IRg2hbEVuM7mcVP4eCwcjtN+YQRzgBG0c/vPDenP/VPnFs
wkstjnv1/ySqxP5lpVQ7n3jaDvhCVky5N51y4tLQ0O3TGfc4iv5SdRt+91P2kQwN
ZBRmTBg0HQF77q43FH5elzHg4JfUES5JGnw6/czugWxqz5H+a3hnLeLMd8upHsTt
3Ng32TmSBZLpaFH/GZCXvmmEMtgsUM8t2ORXo/P0DAsnCh+reSKI6feOUwnyPu2z
uoQhPzmG9glvvYlpO9jI3d5sOSlXbZ6PoNGfRtSVquHYXa03xi4YAcgmIODgytqo
rXoaJW4ZhCmtaNA7uNdF0KShbyibVAPpzHWshLPOF/fEVhYjKVZDnpY6KQS1o2S9
bYDOvvKnmZ5Nyu5s5GFW5yaZbZgk1S3rN5hmL2BYGF6fKjA5i9GWDOWPgHqoHXVz
m32oVBFCBpYY7U2OXtL+dT4V2ztdjg33hk5NeOLXNZQ323KwHdOGwt9/Jvkp2M8k
VJsOWsuyN3pnfiL40x0Qt9/+IwjWE+XHBI3yissXHuxdsFjbJyLHZo5AyxDMn+Nb
5e+0k2bFm4hIQz8QzaGTxnqDq9a23OgvBapCup/+DvTR30roK0LFAv2ZiWUptggY
Gv9gLaLdZMoDE26XnVXh2Qb54i53EvgEkXEaBMFM/awvm4keAKwYL6CyR6jLsC/Q
1XW5LRkRTV3uI9zJzTlXkRq0Te2dGA5H5eTbszMWG2rTyf/4ZIa5ua46Lq6udfMQ
q9CsOzO58KMryKoAoQyLIXRFBUXsi0TzM6J4nJ0Lz/xtcBCWMUOTt8yfO+hqSvpP
thvzLwPP3v5rUzBRJOJ07W/1wFj06sg/zacZ7csLUbuBlEAYKU52kWZOsFGlWbWc
5fSuOoLLBjCY53T7BN1g1MgcIe3HeeOwWCFLSv8Ghlx/KUeRWrI0WpvIZnRrJg4W
VUCWMteaLd5+PVR2ecTqdqJTrrJHjn5kriDcp/2YynQJJpaoqTQdf3LV/MxbKA3S
44c+A7Is9bJEsbCIKg4R3zYgclsclMSFOnCGB1dC918LiDnEA7xa9m1L30ptOQKC
rGA61Q2Q2BzqZGePtItcpVNR3XRr09k+SlJeqlGYpUkPMRFCeEfyR2gtmZug/gjv
BQaaNuarUYTZNkfQp89HYIw4dR1+JnMiU682Aa1JWiRWyDYerBnrNSoRZvDLYeft
z8CijZNh0ZCdW8TiSxpBj4nfbG75juZ62709M+Pwh+V3CMpWE9B0O/ZvKltkVWUz
RuCQXYKa5H5ZUOJ7ykTeGn54HJDk+PJpZwqAOxq2EP5qgQHtIYUD1PyQMbuJo0a2
Cf0euakEs5SuwQEPU3ZiBdg/Hcg5NskeG6SqfU1uj2Ah+m1lePEYV8DPn0GMHIyN
rSuRvwxrqP9JPX2LYwK4wNDXOfF0KuQ0Tx1kclteraxZwFUhb635Yy5YuwHH1ITF
Kz+sy+tyyy6JvALUZT8M3QgBVGe4HaWPQ4iPnam/MR7O3cMxwtuFgw+hdEeq4i8U
C5doATeJzaG7dmt4/bm/iAL4Um83+kW4Lhyw4uJtQwL2YIfX6Ao1h6SyuJIDhG5C
VnB7OwIPrhVJckrSChmPEkT7D1BBky7uFPpW1ScDM928gZimJKI4DOqka/7xsUAY
YTMrGlHHU4znzhYv+kP/cOrn45qqX2m85vLvkigadiBXxkL8DhEcBatDTy3xL8hw
Ne+LfzxOLjkpK+GXGiuazGKHJEwTyHjTYOaKG9fwsC9nEfNjov0X2MyxRj41ggex
U9RrkrA60X0/eWlNL6tVgh9Uheqp+J74i3brnPlr9VC4+EzoUyE2ixqSCjsT5eqC
Ec0x4dXhkz9IvDGhp/5HXjkFuZTdx3CX3vxiHfTJ2tspLc5rCH/W6EcpAPmrAbSm
kf2SVCO8Ex92ZxJJ4wHwkQS0v5bPynXcI1EHE9Y0XJ98Eg2/Rjs0Pk4cTQG8aPsy
KNC+yz9SwFUlWjm2dDTgCZiE1EOMhheClpB4ueW4Nk+9+C7yLoOejchpSe7nQ5+j
JDOqzLFgQz4A+rVvFB9kfxgtoRv+cLKhQC154UdRipBUj8E4ug4MPRGZCZZJGQpP
E7OrNqQnXInuCsq6qdSSM9dup6iOwenN1aHXaT9bLUwzRrVf8N/lU23r7W1WppSK
Me6M+77ZXtj2HnLdgaEq1t78TP71IvsYXTZaQs7nqu0VaPoZN8M804/A8CecjGFm
+0HlGYLuxrce7231b3xdfSQ6FeSddM3Vj1SxqF9GUftSdnJ4iMNGAxGeeqpgLoHF
3Sl6dMM2d6QpaN+RdXh0J2UWeOYjF7QsOlOsTb+cyi12vB3EcTkV51q/vFEu1Sgh
sBTV6sz2V1EFoywWaty7UX8WoA1oEzTszN7ojhDRxSKW7QE7Z9/YCS8aW6VJPX0Q
w5WzddGHy+THyAMGnL2L1SpTu1FXUPTiDA61O9SSie9mBnwxWUK9jkgGn3jF9qp/
AULtlAdQghcy8r+BGAO5fYd/aUulhgXF/Oe7fh9jTz2dx+qc3SY41zsqJqGsFFbh
TfPk52qM7c3f8HH+To9NmrnC8qlwGN2RqUyWXN+9Nb/R4hIjZDVGQnflbxXoRhLv
dgitpU2JlfxBL3Po3YTPveligjEn70chVAI7PSSepSZE5dFgKhdTejTTsL1e34YL
JYY/u8NlUkeRB1yHF/fOUhU40G8VZbfdRoAzcLCWWvTm4HxUN/3yQGY4Uozn14Bh
zjS1MVIPgVi33qgT+V7OhjuZywZfdEh4PnAAfK2QERCYAnki6YHVZZh7RFQ8O9mX
yvds36og6/TmKIUfweP7oJMJrW3zro9U50xKLgcHn85hria6FQx5VwUZqFg9/jbB
LgB8ihHjW8MzjE7ecoTaXFB9WV/liz0BbvCp7NXpOLOW2U6UBrZf/ed3rAs5o1v2
gGgsMyjpu+ESd/VPHSHEobiDHmJWVrnpI/Px6wb5jB9OtBH96OBHJ45gjM131DOv
ECy2zWP8dA0V+QjROgBZ6CC9vhGbeY5R0jvgb50Vc7o114Eoaiq9WrT3qb2iTgoH
0rdu0Px4OyChMRtbX2lcoMXT7u1V8D1EyipUt2pyfwd7xYd+TYT4VXNMQvFRtE6l
dbtLFB3l6IZ0Mv80cBYyTOhlY/RucAPYZsmBKg90BABBEeojastbruli42hPLf4l
NKJL+M5joeuUjnrpcv9Y3nBf+V+QffyxFewH7tziugOmiBMb9KYcf8oVy3TvuJ24
A6Kbf1/uHIwCMdxuw0SvFlyjo1dlEbCM2UJNAr3MqnyZDTNb5nuP8YpjsWTVTe6F
bhWzDalO6BH2cZuJCDvmvKl3dXnj8a2uUmocJjABcubCWvkyt/3fCCTpn+FgeOny
4Koys+FP1gH0Hyavy27G5Q1eqtcGfI5X3n30/4XNj/DVVJz725yt8s7HlLOM1/bD
M3N30RqBmjUZS2nriFzmPzhoaoW7E7uhGWy+WG4mhnxv5iOFO8onf69a3Pd3Pug+
V+XDFYhC7RjHqReb2RI6tsqOySPH1tvvgvHHARt7r/b49raknzVu1cHTv4Qj162D
l2GmcTQdIj/8arZjpWl+0mtmpCVegKHGlfsh4cjQwJl/0WC21tydwlwp2gViVIKz
+xAdkyWNA4TM/nwV6Nc4HAygk6xwnKjIQqmQEMBGI4LSGjUw3Y4Ov9fuaiVojZy5
TpV64QqFCyIp9qTnKvveeR2Wx8v2mEb9FQu2TFmzs1X1VjkHuYnxCp4eiPc3bSsv
7CBeR2yE3sfLk263qnOqG+H9cvmvBo0raZLN1UR3e4K9sei9jzEZ77NANNoYts3g
rocFZWqJ/3xjKuHgObYu1/+ISTAZY1mzqTr6Axc2O2xNKWTDpIphtf4C+nnAyzbn
T3BxaCMYm/ba/4FWOd/IvdAkMJJhU2p28CTCNlmb5TQ7YpkO0j2IUQe8bF9UCKxz
wEXKFbHla4gRbzIxQkTcoeDdMuDGyhUmpNzR047kKNLVyT/yhI5xB/Smni7y0+uJ
PATL0/aiOCfHdBYvvkzHxn4WqSvYaPg3LBHaEMPIcsjmuAIbiAsOq0hMPkWWYDwD
o0oifzCy71e6jSpz0ksZEW707w7FCO3U1j0ZYPCaR6g0x0OUsNV3em9rJjznJwXy
8m8s/5awtmUfvXgWqlrzdqfYLgBLQtQrcng4wAl9Zu66pEVwe3RXkd/bkrJDCxdy
79SPvy7kG/T8SlGAmFJyo7mr0XhlPrGXFbD6AfNatJvHQx5lb5qpAMAHrqk//cnX
MdnXuzXpOzRF7PJdzUhw/J9AzoZszxNUUSyYC1bJOtHPHjgSXheAl+qX1TxjjQVq
wVGKu5+uVzRIOZ29Tt+vGoyBIJdcyoKp1fTzDPo8xqFpfW9VybKnSHzXu17BPulO
Bhm/1ZwLb94DpATWcZHRkpOk4cDGS8+LvVyOst4FaHNPbkWKss301waAbTvPr+U2
wTsRXpKwyhWub/sTGc+sYoQbxPJQcE3G5kUO1lJiXsWKe73i+URXbvgVxrfKpOji
trEcLL74zGrQu7z+fiCAtlfJpAGvcN1MDQQZwrbsHabt+NPw/hAhFPD0UWd+IqMB
bWLH7kfpTUyJqFKvBOpOVeEXEaZDAfWrO/ZppXuePOv0LU8vcKTqIggid9PCJibS
xI5nI+JGczQ9o55nc6SRYou0BaZeq0CE4lpgXihO5gTqcBVbhKOsHyYgiqSyZfNb
6ZnQxZ2GFLwh7NDZNSX+SJoZRrfFqOmxTpgxMH9kkrVhXFZo8rqvQAMQuqXqRiEA
qq9IUs3jW9JDvdsAa4Bilmex4Hnq0hX5M4gybtsm/kLyB2KakH0d11KKCK5PAdG2
eDijGdxvsQAGF1heksqo4L2QELw4Aavhm0RLyrC3eEX59UuGlzsIXM7TzX+Kp49S
cY8gAt3ijfucd/5Vt4BbzNjwFRj5RWjbMbAJYhzDC+0o+Wpkz86pn6sDOU17fdmP
F7B5Gpb1xkbM/MZFSPmEKCHJ/BAhzFFe5EH/Pee8OkVk7b6nZqOW+LooevRZligI
M8OsJBrOoIPyVvgzB1uHwpApQ6Bq/Ok5zux/F8vkTNH3u7jEcDLCm5qpYnu5CQsl
idTGkO1Vp4lHc2ATSXm0Qin5lA6nF7o8wqpym7y1sr9YM/lwUH/09OVzN97I4cSN
+SF58/iaXEYpxxiPijyebfDC1k3c63cXDPZ6CmIyIKYtzNpQw0hl1VL5FNWHOi3E
Wp5pIfZrVvsIm6aKPFRTta43GzSYy8glVJC2qv75KsD0BvKV2CTHn4nqY7VG7RSk
Ll+bgeDF6LmgfgGpQxgMkNi4OvIVxIJsUPG6Kzg4UQ5h3r4nRtxVhV0yDf4QVxJP
65OygPotPiEGp94AxTbZKTgnDpO+1IS9VqQCFZ6/bUdUdXCecyRbFcNe95arnmFA
jYPeJJ9kLRXfkd7kbWSuolZC8iTfMD8uUzGaUeKOfN73FCmtjZ0nWjrDURtjVMIv
2fz1e9vl+cOi/YuDIKi07ZIjv/DFffsqKpjYQTgUQ2FOu4m76/Ffh6EhVHr7LI1S
/D4WdwtyMOtWtE4uXhPMrED/AVCAF8ZbDtoR+GNaPaQ6gCCxbNGaNuLM/s5YTPoQ
PEq4LYV8Co2PRy5gZsj5EzonbpUKyIFYGFglvYeaOTvWdwBQCCC5mgOVDjlu9UGw
f/f3XO4FD1ioW1xKX4g4N5GQ2LCzlZdRbPFvf6uCssHeIHeL3LKRRXd4rjf5/cp0
q3bP/pCbH2cJ/Mb9ssBb1wKCBMicpNLMoYCvB5DuYDqLHDNOz3aTpEsR70+fyg9P
3SPNV6fkyClXWkTBGqHQLMyr98/FgVelGTFyZSZBGtfZKlKMb4VO1Ti4wYslHH0g
8nQku+ksGEwWJPQy74uk2E0bUbq76J7eXRVwbtCqW+/vEv2RMEn2KJsceTkCz91b
0BGIr7QNcPbvxg8y1n9YD7SRe5jYBxbA7LgMXvzoNuwyJ2XsmOT6ph1Kxqkfi6b+
nMrAyYtYtgSC6UimdR+T1GpD29kPfFgHSaWGttVmbmFyucXXaE9gKGs3e17uHMM7
i8ZqgJ6zPQVVD1fGosZ3660a9ZjGiCp7RzJD5Os6pXIKxoBOhjEpkH/nlknpvNKh
VcGCfGWI5DUbAsjiY3VUKXKY2pjBSJ6lIu9MbWn4w8CTisEIv9WMOzla7Ql8IMZb
rUPM7GwmTH13H0U2agT5LbiDlcLoSn0cGTff+hgTxrXCzN3zNtihyPnAJwMd7aHg
f8gy/aN1oJNw4ksBHHKDwsnwMkj85g8bGt3W3q9m9xA7AKR5x2ofvcsJuug0rbAF
zufEHu3P5S9M8w+i92mcIlKrqLbp0N3b37ttXDpBogDtqIok1mtAa35QpM+xWfVu
K8eBLYxRthltyjD+0iF+91IP4maUR7ZvPKJLCsJHQKjIenTw83QZZTQCnjRKQcMr
VT8XtKaVHqAzq039xXDBOJYiZ7ShmmlumOU+BxWvXenBiHqMHe4rtVg6SDtt5Meh
VRzV+Oe5S4HfKaL0VAYpb802McVc6EFNRHS3exB+jg3LfWYffVg4/M4rTGmvlWMz
y3RiR7NPqP6aL7PQLis2AaVxBek00QcIDtfh4nXPVowC+fEYL+/01YwhRKaoOcD3
sHtfhg/VqJRiNQK4OHdrdlf5tLc9+DdW/u90Rz2jRpBmUGZyM9BfRocySO7xdshp
EXCBIevCcHQ+9i6joZQcfj0mpiUyEIrDh4W59kfIMhJdC1KVywsCJUWNI2CuU8dM
mJFnOim4H2Qu4UPZ+b6wSlOmNdxUkyeNNxTGmn016ywnWXIoNYK0aNiO47pKCZ5a
MB3GsJDlA2cxNtSNCHsMd6EVSOpeKbP5HV91jnw4H4P5xLlGzF/DexRzG9v8KDM/
DvImt7u4mSVH9KZBCKYgSDnkroLaoz1tPqsG5KuBQ1FoJ9P5YgjKe8pNWx+Xa/vH
yxoSS78K6MDAgBcW6sEyvY611hB4Axr49xXTZSaJ+QQyt7UmKd795YgEuDrpMTbK
18olZC6kiw4L8Lua8QG0QaYOQl9N4hCculedGIBajuwMUpLdu9amioeYMoBrFhWQ
FvqGYGfZWYChjVBZbHt7eFKAjsAEhRXT+8Tj9/smXD4ujAnFcsNn0m98XeLClDqV
T0RC9pul1Ci8uhNrn4G/lnZ6xYd1Jy/45sCuCgZNIzzCJi4geOSEgMzA5LIefsPv
Z8E5T7ngQNDcsFWfvlp1d2Xl4ZKntsvvyHqXzpNxrdHQ4k7IuNpK5BgoNgC0HoZm
0IdO4lJXGPuOLTkim96XMIp8B+LOWTLDdHJCaqlIwKKhC2QZlIMGTYKrv66HpdbB
cZcTzHBwvMgciZqmtGsAQL4BlMJ42wFRzctncZ4Q2wM828WBopmZRdYZhLWwRmb9
+14sTDFnJuP0WA/w6NuxES9Qi9qxEddHWZdCBJkyGgrQ6Y+PnGwdfH+cxAvT7svR
iafqxOQqtul1LlQ/3asZSF/3Y94v93BlMr6jYSqn1zRKR+QzJGL+4/7fBoZUFNIs
73VI8pr+PgWkGTZWd2yJ9W8v+JGvS7hrEOK45uXw0kqh/g/YaXIRTDITt5EhdhsS
qQvlkhMAPxO4169AfXtYQkpoYWdmKXud8O6L199x0ewGwzGhoFMsiyWWSHBr1M8z
gJjJXcKn/iW5UwJ9XnzYDI+AK6pLSAiGkcOKgEY9KGUK4uZZ/vIrTTDJyZOHwfT3
TywHvEAKoSI4BhQ1hN2zgX1unpc5BbSMLQzhFtV7rj1GTEPHIZIzExz63XnwuiPK
oMQEUFI8BfAlT9oCk3lz8DyFDlXdRGFd0UpFY3iZgO5drLfEwphztPuDpcIKJxpf
1UxL0V0CTapQ9iO70P2Ev2NnlcB+VPoMDH9Cb9z44p5i819P1l3yczq2XxFLz8eU
AXM6xyMeXHvysbpEI3hXlXSMgxs9MdSf/2Kpjoc8I7/ynRxgyNzVge/OZr3kyrxn
xHi1a9UuysJcFAzkOGj0bY3QY5NMXwhBLb2MTkIKH3WYbz7A1TmBDE/BS72csI4H
3R6qCxhiJP1YsIMuvoDbBewaI18Mbuw/uXbXivR8GONRA4YYg7eLT/sdKhYcrSvX
NAucfMMc9OvBkxdnq0q3i8clH078DuPzGkAdK4dx9xR2WNEQZX9oJqKvhv9Y8tLs
KJOoIMuYXM86BeV/ZyS+Rfko9Nv0n4x7T2RO0TjbjeaUoTub5qCkfHK+/URG3PCK
iKyzjUDkeiYLxhw0uWMu5bNOeR4WiSG/1reIrg3MJ6VdALczMcyISmijGa2eEqaK
7xMi6AvWC4d349GG+U9ynW4vCLuqFfIgudTCZIQ+tnbhsAZd8wyaSs+lfW1tbsAo
q4DjeNZiJPhSz4+7bnU01a+XeGNdSl6bjVqPLvY9K/A6thsBhULctpKNRNHw4F5p
5gPU8sKTjXZRCQa0bLWdXGizig148UGw8wTaRRNZbT85Gwrjnkr9cAfzLnOp8yE1
F1grC8FCjNEwqN6iaDF6DsOVaH7ms1Rb5oyl+ZhzVeuT19qrj6AzX4Ktf55uA/Vy
6jeO09qNCiTU4LR/d0OdBH8ez9XHZutYfZjSl4CYSgpZhDyaHr7E8asL4sxWeWpn
pqJOU/9dgmNI8SNJgsCXNn9oOUFJy1Cr1uCGvw3OWzDL+fOOD/m2EjeYqLcholyf
R+VIWm5oO+jcYlIs74rj03bJG5Qi5XL/xjc+5jS0SC9LgLZ1AXGNNFCOUTD+DyUw
MC91DPiAl3n/n8wXha2XqIlgy6cRLOx2Nuh2hJYA3Kb03jKFez6xBnLPZJvkxkm8
vWoH/YMWsTVQXkGiwVu2ejqY22LYe/q2/+P9IqiDSmgSomm3a7VQjGvpbw2UxH0+
t/lUn7t0tdA88+gni1Yoa/dHadwLSAsA7BR6mbJeI9aPSicgWVPktatnlkR7M0sg
xRAjq8YhJ4xtRdYdF2nhc/o0bZcUNxEfuF35ZSXnbdDYIie38TR1hNkJS6dzvZ1X
uv/k/YGB0LYZF3Pm5n9dEBKxjKOydLk8WMyvfkLldtR9eoBT0JMOF6ZpUTkyHUdN
vpWj6KusmY9KtSRdUsso7SvNKu601Q8sHn5bgzNpO0pYyp3c7ga8sZ5YXWrk1otQ
IsmBeyAVXzaTLpYD2M0iSQGXu/sLnhsi2aqVRS34rFXNxF/9zl8qGT++LwGd5Q5Z
bPYFX33KDl3FhiiioGxUaZECVwfsin0XElQh1qLr+6VvwuGtK0Um18us3AcPXcrb
bmjkA1M+8QU53175YCDzve7xzLBNd9uQqYI3Kjmq7PFj8jpCDRD24MyHIgIHJcY+
wjdrB5Xc+g4n/GCQFLpihMhTZMuhqzuzy7rJaBpmrAz9qCrYqldekZOnStMwMj3/
LsTPZtA/EL8R6RtQqr4XzI+yF5wUc0Aah8/SJSME1/3nA+RroYD+5gL4QzY2X09a
OwO90IRf3Jd1J1oQs4FJTjjZPEIL/maCteeibHOSwqltEBM/8h9nEuaEFN28HIUu
DxZI/6uRv4rHjGjAsc5+IWM6kEdF15DA0PJ0PJVUxGC00f2tfK/1D47lkA3n++Vk
BZ47no6scE6CPvyrXfKAnDC9L5EAY2RLky9xmkHSMJO73Ztj/Fi6yeMeXynmMTo8
mQP6XjUjTPlq8IPbqM28N1dLprteoOLKxUy/k32DKubzTWt8P3MmLAx90JqUzPnZ
0rgT8yMU7ujUqVUb5O0QPwIx4hCS+CgNZPOindIF23cX3CCxxPOTIphpuwoo0ZvQ
CEPltTnY4yTiCZzfMucNjCpror5l26tu9NwtDlxuI8TnqDfEMHKIQgXDx2diRNT9
sqoQ4Og+umWnWR9a3S2wefIEpCE9OrN5aEyFOuHxr8coc7itfo3cExnKXd/7lfzS
4HCC3ldex+isfY/fWQIIFeYikH9iHFLEQrCNCK5wA+0IrPB14z8b1I7GTB6TBxgW
iz206FwFme+t/8ebcMw8nXgFB8xzc7UlSbW5vaS8yc9EdEI67AtQELSzjD+QNMEo
nkC7/Hh1Hi7ldP9gnDRC01fiZt58OulYxWEP6X3DPVCRXv1GWrLLmL9YL7ufihvV
+gPK/xQNNTgjwU/m2s+yl0y1lXUdcx/B/CnITQewsq1X/rgVymLlE0hn2b8B5x3I
YzYM5NJEXO81wJHdRT8g95nkAoom8325zkt9oNItaK/WwPKConETdgM+PO/YpG7A
G3bm8liQraEYixDqu/jvvij4pnlZgDG5mV5Cw2wLM4tqKSo06p3+zH5G2YvNY5UP
4Fge0Q4LeNYBSY525W1G0wiv7uT2fCj8G+hk6rNSrQCsGX9g1MHckETQ7Z/6RLy5
wJh6Ghn/MlMAfGBaEylI9ikFbp349NAScsM/jgtdGj+b5Ffou69wMP5AB2T5AKD5
dqWDMxHoZkYfnR9qeos28GfEXIkHn93d0n6OvLzjafqxjjhzw3jqnCbL4YZm1alB
TNKooTJfZ6VQlKidqTW7x+5uJsUJq/29sQQL/6fp6WFXvqemECTQSQGPRtXoW2Rv
Me3ba3YkAAerMUI5Hw4MGDSQ65lb13vDJrIuUFi2yAAXLGtiQaqYXr6Wk8tloHiX
+WivT1Eqx48tL0pt+5vORM5kOnl3zy1PjVbHtNzURFyqpmTzD0AbhJbqbJBrx3ch
sCTRqFzyoMb6Bj9ypg9LXZFT63M6kQepTtl+MLjkybuy8nvV87VFRUJvmgQSdSEI
0M7zQ3QVUTLlRou+ABiT7Tn5pcS0bLxNNIflPuStqLIcjxR5mcYGxpqyUN+fkDKJ
MDErWwpK/MlVr1KnUmc76BXw787Bcat1EqOfmysx5m+mpcJ/PiwtAD2HWr8CI1ez
1BL7/VDaHqguhg9eMridYWgfZ5ir6x2TPTLTMxci6NTOvjjpJIxJMMPPahR91yUw
uXEqP8FIqiAUAhvPkGJ8BGS9gZDU+qJ25Gp/q2X6tap3pPJcaZ3oUYllYhl6Cr3g
KTFSIJzt4yzyZHBt/cv1fq+xxa6DWgyIjX4m6UNmXytR8K1+gYTXXCraPg0HpxPi
miPjm2kco+yz81P/b9G4aPWGHutSMbDI5lzHoSoSZRxLmtHYWPytNCEqbmAygF5g
kUKSK7H5N+iVvZUuxOmt9+A8oHbz9dz0abgTdSJfjvAGbBtx2H+V9Ee008ct/6qA
nxSrCgjofWHve1+T0LZyZE7uiWCEVZqfX2fJPhbikUHuCl7Q3SYkxcO1spek7/+T
JvtbIEWmTsjsa9Zd2RCm6bkxbLjdiBGenJSQcPAfpjrE77qtICvDsVegG4eo0aSZ
MlJW+IfrmS4sXe5ByLT6dALdXhMqyRolEKo+3aiOfCmvWRV0I6qtlc0Nl1sYTBIN
lRuZeNUs4MlbAv037aIPE5QmDsVeR6usL82n/mqrzsPq8FecMmt9Lz7R3/5LOfC+
2Ta2HOvqF7yCa/VODMX4rMAsriz54ZqGUgVWc+xF+PAI6IACS87m1xHTF/0PbL5v
9n5nS226bUoTkAvNSadXGqWdovJ6kLRE5T9FdI2uyf0eqGJA3pbngYYuNYo3jTR/
x9bpEPPFMYn1HPfGL1t/ZXv75dHDlMq6xDflJJ0o1py+0FpKaauPoLZk7djv0dCu
mjYbTIr123yjf9YTZMNooVX8hUfZV2Vj7J4kNsXgq2Xlyqq3PfChJY5VCbpFAPDp
AN7Q3xXocOgck5OpnDWR7nVAy4ZNmsyEOe6O6IJmf1nmhzyjf/RQD34qVFTqNNYm
LqUFy6i3wfxebOeA8/AH/xykFtUIG9KIbXRLtKcdTZkFvoKlmh/QKy2mwhVJ6meO
NMP//cq9fW4aW5BysdW6cnnYe0KqBp4VPX0C1QtbNSGYgVv0KNeKMs6LUFNJAMGA
D14NvJb5tesFaFxegy6mxYy57ZX50WaFcJ+oLVqUXilJPYPDplCo1mtqCy9o69kR
yyXfpMrwu9ZucCVNf+pulC5NaPhH0YdmoEVnqvwkXBp6jPQr0Zq0pW5PPUSSih1F
3ik/HCW9s7yHD5jvOVYK7ig98bHyEGcAg5/z2rH2L7QPAOilaNEFDUgUYLxbM38A
3lwP8gsVxltdA/vnqmcMSPxtsqHE/5HwGXXB1oCHeHStmf4ULyw2tpySMMJO4N0p
yfLYvJeJd59f6TLM3tMIPjuJ9f7seCpXnlLL+8Yyzptbk9gA0n/w/c8H8CxEiAaU
YLzoUtQxNDFDi58I8lORkPwhyJEdoBiDvfCfYY01YTK5Sr6/uiWi08g//VZoo4Mq
CwDKZM+BYrhDNRPrNT2JF8KateO4L+8FDFwpaX+jtdRmSpv3rbv+KF8ge6hoIX8Y
56r211hhgYGSadtuJfpjNwirLZeapAhk6exhB4OeKphuCd2KaGZzyIW9uIgxGfo6
cR89P5Q7/ZgUKR3nDlrVVtQf661xx0C/yn0ZUsUZUu4U12hWXqmYclIp3JSAzVpN
Tkgg2yzUKhyw/mhMvhO9tpwlqj2K8RZ9r5F3b4+vZE9Uo/FiNxQc8HhDuks+r9Kz
KcqQuf5k7sfRa0GycO9kSnb4vaABSySn006qvFZUQa46JRTJaj574Jyqr8YGChJQ
BSlq+IXBls8upQfuDyIJHvRjBqK7e/DHGbz5+VRidWU1D3UVmCWYOR0bJyZ36BnD
an/8FTSiXzsAI8dPWa/hROsOaKVnPI7f3VDdcPa4Bjbp6qTVup1jQHnaVqoId/Ka
Sl54WBjjP2mdNIbFKoUZrYWdM/639kHVdt4EUl7uLxgPjfKEdTSYE9UeNdeDpxKO
uPgIXuvmz3fmd+K8CAR2yZGjlWgGCSg4UYJXndvylktVuXB0TyxqlGNOl3Z6ER7X
HXUn9s28dL2Jrn9HnKH/l2iLwi/UvCEAOiR64Xxp3nVwhnOnpiTVeIdVN7oTOq2o
I2MuqtklureBSrT69NPcrv41BvDrwE1aAiqiOnjeGoGGtBVhB2ZAMq3NUcsZClXQ
fVQQ9SAzwVsxnC0mAn/ffmVexw7JBk6lfsCpHmUkM/xE5QHSj7AatvhC4UBLo6lk
8kLVHCYlfuhjNwu5GLe+aQS7GDMLdmjtXczqrz8nLDxRKQGEOgPZJfUylx7nqyiB
OXR3564fUKpqmtEBdaaB2HcZMPOvMdcqX0F1BDCbwd7pppvFrpOtZz6ZEm0A5I/m
WDLhTQR0k9+Sd1mzjRZAwvFlwB34XYT20X1fYBCzaH09JoNhEZ54MnvoHB7UTIXX
ocpNvIdpccNvfgNO9DF4Hx1lN81V5a8cFg+DEOqzMcWT8amtfzvNEY2Y44VgGAdS
tT4mJ/vUdnK/olq51AktUrb33RjLOnwoDNw0br+x20E3ojzvEXEpkqPFJoQsB1E7
99MH61zhYGkq4gj3a0GPiSE3RgGlOp83JncG8WqwSstEj9qjouWhT20e+T8t1vI4
axuai8K4rWVYtZHJuhG2bN/nWiLqVAnrGsu5iJhgvyX5queWEm6sR6GBwTbcEBsz
DK26XfhlQTUIb71ucwi/hi0IhPCiUAOlgB0uTVPUy1aPIXmPbxbDc/wgvw+p7bPL
5l8Akhef71j+4AWteD+vfRRs08DLRfg9JKWqCl+VYgO6L1H1pdB5SoWV2COBJDcr
hd2y6y7/ebMbAN+PK1bqVhSqraMu+okGdBM8QpMbqCwcwkfKqpB8NfoP7pd5WQPw
KoMpgWy/8RvZQmCbrKSsjTDrc9+QE8NCydx8NzPLAtlA9Tq/u39LFm6kIs1ep52T
HV5iI5g+7N8nRYjNLmJKo75iMR4tiMM/RNb5CMcuZt6RZic3oH7Azs6Pu3Bsb0Yd
hswYSnxo7g1jRR6aD4/pT30dLxXkICTnsCAVX4kX7R21IxoEs6a5FUJvdhpkwDQN
nPSGPvPP5zrSrgli5A2zYspVDM/W9TqlfBRZAg7ngoBt+4Z3isC42jMemsnBb+2t
5SqYxx34ieECYmpyZZuSd65EXylCBBdrbvu0neATD+OzbJyVJnVzswLHrCDS7Aaj
LVFUN+caz7s0MTpFm5/px6TeUtbrO30l1rJbNraHgkbO7Xgw3y3F47EJTZcpHc5f
f4MB4c7iuKZwvd55S8gT7JW9Ljfs9v3imViYEdOzqDXd1oJ9lMqhBRdM/eg+jDNY
Z5C8jNRjQ7JFCreLfZ4oS8vbW5KLHyhwPgeoGSzrFYh71mPWs9abRhKaLXRjoKKp
lncd1B2+ED4NsRDV34c/KD4eZRt/U5uyLTL+FMAETtZTZulMu0EZHFp3tScnQGNb
6GnsIS8v9psAovry8KXeytIEjK/Fo+p2KqNk0rmxLfnZbGhe6LXpoVhEZYU22l32
Ix6m3tn5X0VfPM7MnGKFEwPQTpb87OkDkgCcq13S31ATy0GcoME1tmxsoJ9Upt2K
BDvAboeF6e48OK++0fOQ+02hWcuz5Q3IuD3ryfv5IoqIH7wYgpv8UroD9HD/DCzB
xYGeK1VObijl3J4eg5excpFZ3n4BKFXexxIcwdM2WQB013UB+V3R7wyzIN1ETxsj
127r6qSVx6u3etoAWvkZYV7eE6Xckiu6TzgzGpTWGU2zbQ06uHvQwt53nJZZeR2w
veNUxFWrUQRD86+Cp8oJMvLBcz9dqyFoGopeOvEsy62g6H9zzAoeQZR139t4IuSm
OdVcI/5oE4vx7BM0Mg0gHQMMH8TIomIcsjF/SPkAofcZ+s/nl3iZGqHIEUYMsNfh
zWpCliddzIJJissVYOsSsgyW3yFEfoDFmoRxsBRrLe0JeQKs0+EognNTUsYPZOkV
oy4j6kYUKpO3Dem2zwS80+GqOy1pmtPQMOTKx43Hcvdga7T1L0aDn1ioFk1aKMWw
0ij6nvJsNX8fN3ktTZn6g1jR1jyvc08rxtC95KbXhbqbNsseBGiCTcmezaKivp/5
rPQFXXmhT1VdTcHZq3B8M/25Zp/yo1oZdWNo953eBbQfdie2mEvmgOSSeb8UUOVh
6eIhYmDouCcfoLahRDV0aT31Vid4Fu1UB9hv7U3eLhruri+dGmIVrS+s19jcPMRe
KfwMDEXzXcHCmozMcROC0ZECA+UwAkCris3v3XDecNH4wu1ITL56U8aoOm99XfMe
6BvUDGj3e1IjA4I7bB5dPSP5mf/VVUuKfrVnDsEhpeIXd23QD3V10r35Ow2dDfEH
J+dTlpNeG6wiL92eUPSy1pa24QaFRnH3pfJd/7w3HF7lt9oYWVFmYIsnFdHrMStP
l6NKOJMdgX5X964r2syn7yIeg/d9edje5Qz7zJeMULSlBt/TD2wNpAy32zYIxodk
ZzNRHjBLA+suMUtUYZZmnKxM2mhD7VmA8T87ngEJIB6M/8GtU+yfyuhznV1DTiRO
GY4FIK+OiAMqvVcY74Wifxf6uKbRg9n1waf01Z41p9r1RqreNCmFQd1NiZb0cghI
qA3wDhAbJPEuv3jY0ijDLxtg54zUW628jibRd0jUFi+/nRQobK02o7t5fEvQYlmR
n9/oi6IPS5DFBDrWAx6HwFVrJa3OjFsV9cBGBt2zmHMPnMACb7c+QxXyzssqEdrd
sBLc+jUGKNpqpdo7qyFYWF7+4iNhwYoQ0n1Or5FPzVf1za1GrnwOKcMasu4Jp9ht
pfdLjKxJAzpTNYuZR+U8FoqqNpyoL6/mxqExNCSPsc0x/PJPuWniMR+gAh5o6h7X
OJOegKRlXgOXggXG2MuyaTpuOrCDvCAm+U0KlP8N1K9+tiY+DydHKEw0PXPutxMR
vE5TXC7dsk6Le198IaW7AaNMxPUH6Ub8qFB0Iz+Hk32BDTUZcRN/S9iFhSKhj8ZL
ytgR+nWDPDwuhdppMAlYmDwiag1rEtxobhuOBwth27XJ3Apw0o0TsaldKoWjT1Ts
B6xVd7CgSGBFRKfHlAGSRrIipMIG+cZ+nnmQCxtd0UfttjwQi/44ZNUaEPaVW6Bf
ndQcPYDMSCOoQNDbS7fbksWnPJ9zmlgo5p1bZoMj7QDeuoR9M20EgtoHudrGIvnt
8sXqi5LQgIUDWlHiWLiqOkfKsrySemfl1bGaR/5dV1UmIzeoG3agtSwbJx7pP57G
Q4ewgydwruT5U1XgQjVoVIqnkMb+WUJPS95O9NAN4mMfEciiam4DAWjUS5jykIdV
/pXqmqFutxNc8zXpxkCUfq1oL7yCCsxcZ02hVYEpkJaz+99kNbn4X358lTu7Qp1p
vv6DbYB2r/PE/cd4KWVEepBlKO0JlP4vYd/7fLlohsIxVPRORAacHYDB0WulbWfY
3zEctjC3e98CZbuW/5VulZ1h/V6ewRh3Df+uBzyusbT90ggYo3nspWMrb8oKntEH
y6jIg2+x/wrpTIhiqBFlGBmWTO+LTWPgqdZ013cw33F+AHb4UsgmT2X+JN++X4N3
6lNsm/1xFGFrx6VrXCODWjjoQa/eEni3Bt3SQXBs8CM+WssWcSZoMKk3stzcXUIS
kV50bKdGHU6pldPLTVfJmmU2qYRLowDaTfsCS8xSH9OTPqk+oiXAXuvpJ2G3nk1g
tcPTfcb7rqZF9mQwwLKqcpF42DViekmdbkJ/H8ZOugkwI3afbbWSo4eTjgxhXRqL
zAho07Zy1CshLW9/n0qu4T/uJ5+8YwkfYOEkTWKOlfsiw8szRna9dcAdYhOzviwi
+hQC5bA0WLK2nahmKK/S9np9lwv5UhpZuFEtckjSPClcJIhE9gSoUJeTvXIbv588
uux2AShZEW6MF54CnE+1ko3MNxhB/+7Sbjb+8qSELNJkYBHGaMsoLZG9qfDYNFoK
iQNOtxcnOpV5x0+O/0+LTFXM3Rc++IHKyYtclr8EjDu0dnF+SfIg3+8dQUzn3NlY
MqBnAY1lolPUTyT1MefdEMIcOImhPwtTAhJ3EkRMZgN5yc/W6lambqQVzSmmrBuL
efZU9ZuKur4lskKpNnijmLI8/9CGcdDGVRxKnSihHl/PlsV8hs1kJ//JzplnRC8x
MweYBuxD2X0rpc9hzqDfLo08+1jg2qHiFwszC+Lt5BOdSt7yGEIpmNQSD8a6fvnI
G488myw9hxqULa8yuG6Fq4RdOLJhkGBwr+rYZeoGj02NpdBx38rJgZXpEwgvNXU1
bUdqwd0zu8FOZjXB02ZEV8qbGX3slsb5hmU6ofwQrdWOMMnBXLavD9AAyEdZX+yb
hYHuBmaZDI6kr4l2luOcLPLDkwpnMEDDqy6xYMS0FkymhuTLSbZE27W2XEcoSDhP
MXE3DKzYCwN5ytCGqlGPSamtjmjJjcTZO+BrWR1tm4naPL5FK2YxXsIV8G9xwOOg
oxYJbsEPVIi4MqXZ1INkfJxsxDLOoc7bkp1rzB8p3mmFkqEaoisyZevqX1djOJon
TH1kz5GELpPjLQ6/oe60QdPehgIVIewaVxP/07UXJyIuKBqKwCqRxSjWjAHiamam
gKNc68/3+gs7yBDMtqjmXBEd4S7UJPmZ1MJcK6+Yoj/Bd0lFJ6DPWTlxIXszptQm
TJwyE5meCtax3CJPm8MYm7Q50rO5JxtMt8v/2swbR8SoTBMNV1xvuEb1Cyv/oCxg
Y0ubnvpLmHPvZVssNziS9xJ/jSBq0FcBzG33uiIYNF4EG2BoGdrLCmOJDV0LKnvg
zqJFeZk2C9tTpKFhTB8QTYr/lpoNZ8e69hFkEyGcMoVUbEvMPtEirhJULD5LGe5z
oJjRqwesOgBaPjvpfqwZkk/sszTCpheyGoZR/pAjm7wZxedzka99ZFgP64zx+AC0
BxS54Ku/o21jWmtSZhs2WARjTQDYj/6MOVyxsQAPJwH/1ZbmBWL7hr0wn+bGfsDE
2GWNuJJCFhgBtGG5vVOEBwFU9BKQ5tUYN0H9BEOv2/2OH1zI2XWtlJcJRPH9Fs9M
JVj1w1x8JsIW3ZaKdBo2kqAzcJ7I48HYvI4grTMC8Pzmh/LByeoiMoSa1q5+N1E6
g+LeXpv+MPzkiot3E/pR/RaZWCIYKD4C7mmF7wXOr9KmUxv+WoK4GFkbwBd+65SC
BDVGYFMDqumYa/48BxD+DxTpsIzhYaW0IUBIgBMGwl5zgjbEmVMTUjDSYRzTiCG8
y/uqm86w5dFovT3fDqDMjdmtieLzBSn3TwfmqVzoM6SaDli/QqSPgeYMkDANYeO/
JQ59jx03SyXp9BGqMg9vp/i1KIyklukkc2YCNH4ISTAmJGVjkGCCJD1G4WOSI29t
CYjdVoUN58FzLldw2KemQblO3ZzX+OWfHVd9RMgHAgSMV7r0u1rZcXpK12t1xdPg
cHeZQPIOJTHIQbaeDBwvJCi9UJbXDIXen75AETTzd3Fo/3u8jEBHbiFW8DlTtPw3
z3TO2pSFcyG4D5hcSSxt/bDRUW3onTpf5L9OUVMgIMHTGWIoj3Hc8cusBePaa/2M
197AJVbB9vVyG1B7COJFC8DqapJP/S4xHjownuam/mkzutiPJm/Dp4ZnNuYou/MK
cndkQ6oROwVXhkVv8YFmh2Zj+PQhx6bQRhayz7stXkKi89jStgpjcSiGIgnaBbEf
09XZ4xZ00ors03aLpOz+tCZ9UJyDPHCtPGH2WbsXhwLd9qKT+rMh3vSwebhcta10
Pt/DxgB7+W9HwxCIAspaa7sJHCTZE0Iaw++yVB0lGaaXUUIKhswlQYkuzEHAFc1W
fWXfG0og1QwFtY1vxJ09D9r6R5Hs34qUbmf5PcAdMyJEZu1uh8LEvfhFKh9PIxiS
/Zs5mp5INioefoH7kpgAoZ6tLTEBMCYDW+xairA24ClaVnCuLALDuUk5sssKW5c1
ernTUqXJ0dez/PJDIG4Dpum01LfBL6FR7X/CCubvrywGPuqBd5FXDESQOpwgH46+
3hTY27psWf/smH+BM+P/ZV0z6w9rRHiFgQGBUmT4c202d2bE9aUjwF0FcmCaas+V
g8a2vejR5D13oLLOH3IFak+cNrab2efHyLwRsGULFGWibuF6DH6qx/2U3gITL2IX
hlpM6lcO0GFcv2qwv/FAxSLMIy21QSuRmZjPTWepVVS9MmjbKxjnJ5879sGQhcg+
0WPvErLIuoyj9aAR7eJSJnQjNvbstuYYjtvbpl1gHffnS/RqI5n5CHKxgy4cs3mP
m5NtK7wiWR6KgfzbhzdD8oAzuT4297AFbDA3VpLXK1KABG+BRGmufEmhM5LEVCJC
FDq7ILU9vMTq2oRLfHBLk3RxuCltLWSZvVgz8sxM5d7GnKtufGgAhieQK3xOZsge
+qVM2Arj/77WJnpbwlkSZo9xQN1pwaaPiqZh2BWvG6qjMpG14xaSq6A9B3bhqe9+
J3UCzHjx6n92/mSvvuHU6koeo5bbvp11ti36vCycm5pC977VekJroTWNfRHqT0Cj
8+GcZvI+8QhoSGXyzGiUkI79oZWKYANqf0FujCEQIGWCTbt6ZY6wzol4hXpSTd6+
fSZeXqQ1AH169QBgjQKnWmwtjEsMbQQMjts9n5StpVeWPHO1TB67uzXXw12Tpwx0
e1HePitn+DVLb99B0b/jzJjWKK+eRrg47ZAjBz6Ny4krPgHIqgfkgwADLhaMRBFj
FpnnbrbnqiQItZB9qLkC5yNSYMUH7KghjU+Q3gNRiNvo3papJv1lhNfN8zqRelx0
sPbyrkVkmay6tSvucgNUZrhL3S0GcNCUKLZlrrgtuG7mVA0/qT/t+/lyldK7H2sq
U22U71SXK2bj5DmJzLEjGPwwBEZow8i9RXoRIOfCPIO0RFPt46zJgfdfpfHoVNBu
bDWTRht8VVZXTYpPC61WLIdocCTniA7wLGKAKJ/SYhP/NGQSGAFHlIAzmPF4y32d
8IhQVWmNTc195wFcAjx7+rycdUCpxn9XaSqJjaRYuZE40mOSVYxIjH14MP+RhycN
bpEaIYgcXkFcgXxajijDXpFflusEP/iSFjV4wFhY78wNkmhJ9XVMO2aBqbeGi8Rl
aBjvNtK1hi2oBWDSfBAu3TjrvyZ8ezwIP2P5vxDYa1Y8jko6SwKCBn2qm+uhJ/66
mFzEf20/c5T2SH37bTSt+NMel45UTOp84O6t6yPsLwA7JqE4odSji9Bs90V0vP+S
oAlvJ6ipf5IZbwbT1hmEhZJatxOSNKSq9jj09QKw5eIDHqCHxzNsMrSMseIYUZWX
dfDONgp0WpxYcfSA9mGAEZ/F0V5dxrnWFeMxla/zbc8/ekLlzSmsyxSunWB3Y7NH
rm8xd/3vluqkP0m+A05or+hGm75PlwS3c/H08KJhiSBy/LySxnSksdd1UYbZxJgn
aWh2CTLyRJahVJmxbF/VXAfX2iAqvy+wVtrVlLa4PT58YEaArt09PaKujEGf/EYP
33nei5M4bbv3q5K9aUfa5XyteD1G8zvoaJF8/9+GzNRqghRbTAi5rB8Imfaml4Xs
7Sz9WOQVVRhOwmHZ+PGXe2AJa2BmcBaXGHeNQPJCRsF/iEoRyBDXYdJA7/hpQNz2
MFaPo6v0MvFLo/D2YHNT9PC17Z9rfiTNqF5ilPnrRaiqZIc230GzvbVOT0ToLnI6
iLcRIjJyzSvwdYrxwuHKzmjCsMueLNI7hZ618+NzQFY/7ld7UaPIXLaZK41ok2Qd
0TS1IvIO75V4Ly7/XOmQqFTEU1ggRL1X1XSgERITqgzQ2eRe9Vet+kOHzHXnU4Ye
FH9vXnNhSQ3JQldU0RIL6uvLy2+rc2lK3tjvfmabIKu5EqJiXhB8Cq+2srfboOiU
HOOY8E9SKYUVGYr+JC/DQvo20xk5UT/8qFz/7ScKV5wBInUgwRA9Uvs6wxdKryi2
Ufg3uByHB3wTURvIXz2GcdrCVHakUooZ+v8wAVS6cx77IMiri7XJ3Tc4awRKYI99
lX//nIp0jq9Yw0jMFnfIlw4uDW4ixfn7/KKqH6ZjSR9h/oXAVeyx3oUDLreLrjsT
zWNjxFKKx+QbhH7/FD3BeIrBPzSEFP0ZA3H0OG+2UB2+GWP2AfY30PsEm+DLAHUq
pr1l6t7L2RhRTIZ2ELBcivYR6MhDx38yhKU2aBA4aiIH+11rsD9I5dCy9Kqtu3XW
z7UEeDXw1oj9sq0MibIlbIEroMR20onExbpqsoCAbQvetn+J+SFmI7ojNeizF4mJ
jBEmUwLH4fuI7exStPW4sRrJfTD9BehjmN23/UBzitm72cQTnIvzpcV4Q6gjfDDw
rlfSV4LEXSrS6fnuomRnAXkMQ+MpprMvMhtqmZeOlgxc02ygwX8j4d7auG/DqFXj
zzdMBYvqFtKz/b0uPX0Aq9j68tZw0CB8hTqz9ZcfSKgg0NpXWcK3UshWwvu+fvmB
5wO+ZXAvEWsMLETPSxwBNrGgDrPZRTJklOntbIxkkPtQMugxQLWzuVO6tJvWkjDz
smwUpDt/E5xiwzEKjqo7vgpSVIDNAXuI6WUHRM9sS+jcfLgs8G9cUeaWSZnoi3c6
9BwGwgV9R878DRunE70kwbLgnuGlmmNRVJDHKwq4lu9pqguvbRFkp+jLnexPBih3
unyHbDRhwSACrlrEH3X/XvJ/s/Jpw26RElxtT6coVaghcVD44KPlIA5zGqPk4jt8
/Y6+jWm3zvGPZca8FUrQ6P3eyoTEqx1MVn33VVf9G9Hs1GcPj0+4FviNcqeg8hq5
MJhTjTp8xgcLgJ3PsXrx0vRq9+u4SrlSXOqwf6LOYz37KptCTx+MSvLObusZY8vO
If3V5UBWlEi5ZSoZ5pluc0eQBRIZUL8cWaXON71Q9GTf85hcmBkQwqmTArWfhPJK
Fo3kmiO3le7JEiWNsUEgm22HxrJWXohYjAlJCug5BeSuEWh1aWa6vu93HRc4BYNx
SIc9BOpvSB28a/bZoNMRpKTbB6t7bXwKG+QaEij+psrzIhFKm+llX0AMi2+RHZ8S
6qCo1urnwBRDFg75ew0QUo0lcyc0o51G/n1ImyZQFbbJRhmlj8g1Eq76+h8zV8tu
A/15ROJ6z8UWo3xvAkHaPZWoa92/tl8QiE3EijP76bebBb22y5CX8pImR7vzPKNu
rRbo5vQnvzNLdfy4TleOxEOqk6v3PESZH7eL/6tsSnsv/oOboCJN5giXv1DoMSoM
QCczOWCPhKsLNRLL33Pgm3S7cjwfyiN7VCqTY98XApFQ0g5j8M2QJwXEOVR0BQUv
CUpI0DhGG9LsrPV77PcTr0Y3UvC6zUtQwOss2t7rdajLqCEolc+CPQWxeuDHhYHg
/rjtVPUDdm/crDGOZgjm4aU8SqQwLjamCrV5DqL98M/H2QCN0XmvGN8fwMdFpZsI
7cnKesYP94G8CVXU0RwGg0NOLUw+bB6L5TOvliDKO/t2Vf/M5RJx2T8vyvqf8WdI
JNjS1p3cH7Ji5NK7JFecVeJMbMqEXf8cFZ2KFXsNVHh3518TWI0FTdZES7vJJWKv
iyy04HtTZmh3AJj0+lah3eHotOGtux4PGei3OGYHC/ISTVXqQPM219BtE+ixzlA3
eMQ4QOFIJpMp6OEk7rCB7NupVH7dO0GvIMzqlR/LOiHt5qFnApwkzWCq2GNnVFL5
l+etqPfeXbv0/YrZG0zvEKn59SrJJbmxrhDU6q9NMX17NAkZs0RqmvrU/iwxDqly
0JDGJfiN8sIOSPSEAAqY86B40pmk0FB9jruqaxhXl398E/0DfhcU/bGPH2npT5CL
W/b526QKuAhNFiB0FSjPo3pQwpMFZyW0ehKwJr/w2NrjmPj3l8tnXs3qom+wLm59
ZtWNtBmtqYSHfQFCSwtRVp0fzrY1XeuUN9+sHt7lK7wVt/HAHgMWLncWU2ew0R+r
ClhhV7Tk4DpdmHWpzbnOfCGvUdjeDDO/Q6NhPWv+JZk5KKurvPCnK7gNVZztmfpx
4cqgtJkw/TllVKIVBYQhj0O6+Mb001bvBLmSO94YPCQ6jS/ZKYOtd0ngEDqzOUeA
ZikrfOwvXcaSPB3si30whDnK236pJIsRJ5gs7RF3Bnk0A1NVy3NQ7gTMy2n8ISKj
hZ5x6hSJ3RR7d2koFt1jQagDcEOZuPY5fw4KAK5MrujqMrUWdem8Qiks3QQKCimP
MiMdqnLxzGFjbo47PuHTeWakmRpmTyeA491gz6/Jx0AQshW7qjqsvR3GFh7Q9dLk
EyJDL/NDZYwIGAWdpwPYCCOeVMOJRONSe/HjSji2viXqYMwNb3tW0wLsumBQIns8
0xNWAK3hyxU8n1Hv7JF0+UrYf6HCtOOFRNUfIYu/oaraf+FV5FusGSycVC3TyHEU
hYjBN2zlCP5FN61jcI01p17C5+Qqi8Z8v4C0fy1KwERXX0JiZRWUuMy37hVIuqeL
bBgv8gdnolD99m8Vws9Vo9RR/Lmra+rOQ+aFcf5WJ8IcUWk5T8JxKyGmL3CrGVDU
CoFHencpMQRWez+n+Z39Cn6GpUtiB4A4Bi0QbfqD6vfJRjfKtXGtp5NAOOJqPnzo
qSv2GuVjtMj0WtlyOi2KkXH926Gcn/K4W4apdeDm8kg+ZLQLQoPRiRRAOQc8GsMd
lQa/93hcfZTHsa2srSsFa0WgYy+w18x+HKfq2wJ1oiD+mpou8QN7QHNz6/j14T9a
XK9n5n/swOUs+oljuEyqO9eyiHviweXfkmAwHtWp+39cjlZBUxIEyKaJXAF7WfI2
3YouSDymfeGR4ZeIC3tWnD6z1phKMJ+xqW0KKy6MsZoW3NtSzPNNqtJaM42jSvIz
0K8gjooqyIQM4D3+i2yndMGtBp5QSDgkRkGEQtvvwW7I1zr1nJAoATQXQsnfxn2X
m5gr0FG+5nhfQorBVHhyT/elA6HhXAMzomAQrinJrqmV4pyEgp1o6JbqOvC9x+g3
67V7WN3vca8IDWzcl+snxqb6w/rUVNFekMqdPEHfZ/gXnCjzMnrdYWgcZXzx4518
1CELurNOvFh37aOMnJ/U+18/W/+GBxIHuRyAZqUcAfsoK14JkXtEbkau/59CcPSW
j77f+mnbkJqCbwOWe0uYQ4ok9Z7DI8tpZhIXewOJ+xZnZen5NLu/oJ6ewr5emPbl
jtT7iFu3j4gYKaygWOrv7Kww7sAVsJWWa5ZZscYwfu7tdVXh9xDsD7qVourw7Bdc
76qq2MBDERxhhZ/1hoELpKyQJWpcVjvY9TaeBcfLMkzQzP7G/azyVqj50jknFBnX
Iks/sFXYKhgYrdDp70W057XDaeBQDvhhVx513N0jTr1v7XCSbL+pPHTwcOjBbjM+
NgHkxLzxcNg6vQnrvO25q96KNplwdUQ4lympx/GulA+WicKvRP8dH3cVIzJj4XAL
2gK9riJC0v30J6aUSimSBk7omuaMj1WtN57LhwT7DmYK8ro7Pr1K/Y8wjQzeoEFg
kZzNSottpIFep1HfamJVZRQ15xM9A3TwRAbEAVmYZwoSpD+sFTZcfvQ0EtYs+LoC
K5UmQvw2VUEEKBfFz1RqnL5gX2PHKvoaRxgZjPfliNO9RRA8szxXO9q8zRBaUHPx
oNk8KLBcHpMAMYZd9OQKZysULfUMR2ml084BfV97JBLmu0kN56Fl2CGxsF0rVMPq
ixrMg15Jd2VraVcZf5ACF1LaWchYqeuIu0l9QVx12M91dL27EWcx5ibf9FpwHEaN
NHRWUKBrSpoZ6Fegc/5WrBpRG/fDFLjCpRIc9x8mFDhIVCRsS26aww4cHmLL0pRw
WHNLvHMNqWAg7Dfhc2bHoWLDuFSdl5zLkvhkcKjcf/4ywOy/UMW8xjV20fdOoDxj
SJwyhaJDk5KAUfoZyhylW0ajEiTHHbzuHZfmjI6lWANQivrSMQ6tQnCntkzcRnGb
15x1pIpfawaWnVsSd+fDajrEIBwaOsLTavkmdbpkdDjSgtEWRx8RGgcD1LVhlz2B
3T2rjazIEX/F8paqphWN+b5caY4sChjP17iuo7X3AaFCzBjgG7xxERBZG2l6ylP+
awrqgfXgpfZ0MVLTtmzmLVDTk4AEnnGoo5doF0S5zQjGSZl8WsNXZbnTvE0OyhUn
J/beTfQTR8HhpxuC0HSU23kVGsmOC6Ejyffoo6nqK9J5FjokM0FFC1psAMnTaBsH
TbM4+1/yTDLujp9vd5di6y01Y4p6v6Jc7RM8Qcwa/VBu93WQr6NRn9j11oh9HI5z
Fb9BNOm5cP/dzO/KJ/gzrACHrp8yyVc/qjzaN6W+TZkgGzYS6on9/LSGOGGbH2r6
Bbpzy5rBFrga0iYdO2XR4SuSCj/VA9T/hVGmYupTvoUg1M4n9/PvUGkEJbxpnIYF
+yF6ZLp1NLO/IRz9osG06S2d81+nhDbJo3yXZS0qHxeG94BGsbjRlIq1K9eJTIZD
B5dIdsz1T+FqR22dRi+/Yr1tnIf3z1Y22emtAhomVBCY5aEADh8U8dU8XgeKwPE7
3zQTUmlw7G/01bbQ/E9ACr13nvMNF7dSC4LOE8jNiG+UekWJS0xEz5rpGArZDDiN
tJsb1BAoFB8YKJBssT/fbPEk797BntSLY5F0effRsTOqk/SSrYlHdiHKK4bvRnYy
AKjV4J7mbJeDYjPqqm5X5W0o2W+OjWMrhx/UzTwQzORyI/vBsPYibViax5j/v3Kr
tBKgQTvB6gcKe/bPpOwoRF4tWiFiZ8uvgaIluEV21v8QbmnSpvZce+H2h1RrlyDG
qeNC+btStT+HWcFko8x5Td0z6NK7HpR0/G+Uhkx0VQ2H466a3xxDBx2ZIZfm3lHt
3wQtLVIxFREPPFDToO3mtP8aT1mt2Jn6jmyjee3AK9XacpOSs309q7xWGnt8ZhJt
w5czvNib51KrAU9ddk2T09VqPhDwISHNFYUEi3wZb4M7oBQqNxGSWhZcqTkKN89b
jb27n9hHc/yEDBjsKaGwUSUFuQRJ5xK4r++o9WvBKF7U0Xqzs5SoiauFWd21OaGS
JM8atazKiK30HgIVH2g6BTYrq1/HFcrn3zIHYQSuIa3VKKdQuVsFP4YC567QIopl
+rcAkw5b8xZbfw3byzWSWbMb9RH3+P6QpqmkQ9s0hoTZpRPJGbSwZLAfZXAyA1q8
3B23y/k+S24amFhhRO3ScPELLqwK0Thx9ZCBGmEnfmsQXnwfhkBQwWVCEf/ZlRK9
L8qIqPH0knmzq4lnnJcjqi8S+mlL6xMluKVrce0sqLDFiFz/2D0eemH2qE/tPW/D
LqU6nYLHKjGDrPa2NShjiJ8iCNZ5oG0MRNAoaQkAD6PzN8Bz9bl7kUicr8zI7DBi
JHrAMzuUf9d/5Na/cf2osQgCJoiRBsQ5XKYPEKVFRJ3rDTjy+pihZEdUTEyMXft9
4CyXzFRs/i8rmoHzwawAuP6J9g6tVMTxZaAg+4kAfidBm6xVWJzta2kXGQoWbe9n
FSvdUSX+8seY7/+L7R86bvubs9Fqqt9mxUN7tBHBc9Deo7OJVwNzaHJwWvHzenD8
r/pZJL62idc2gBIKNeaPO5sQX5Egx1HdL/Dw+AKkXv7UuLA/2SRp+lAHrMGnkRC1
4G+pMPttHAjk7ZzclwLubyaXxoLNvaq6AC03C+rDLkiiCWHB8JtU8vkmXaQHUjnG
8tf71xem/OnXWiQqPvnkNmOARSOn80Uij9n99oSUHoCGrTWuO9BstUuD/Fvd+4ja
ZFalzvoe11vbnog+7PmEcqc7Tqtvq84zM2V/Un90zV9I1tj52JkqYA3aHqyj+QOr
jWNsRj0/1RbYF0hmUnraYEDYRj7ukOf21nmpM4JZ/RWS8kIcG/x9ccU+K0VLEz8b
UJlBt5IhQJtWMtk39xDSCA01eNotvxh+lsOO3xl/bfdJVCFnBDMfkqqRUjtHJTiO
YP6vtaM7VV/vJ+f+4nYmbk0LZuu/mYjbh2rx8H6dIoY3GQOPhupg4HIC+x7aTt7g
Fv/+JdRUvC+4wKKpZ64eNwiIN8jd47KAFzr1exE8cW/Kpndhw54NJOZtgdaOyqlw
PSanuHd3P6dyogNSFMddZWYsfhzQe9HEvzftxMkoaUTsTsteU17QTYGsz0aMlsmt
hhnJu88E/DacfKkzGtifUd6bj8vWzzCjYIAS3jJTnEZ2W2TgTGH72oQCnHgAoxnx
gIxdtAPwfSbKy+9bmU6OhRvxuSnht9A8bHMpyxF6BgFUJ5gqcMKF+Hpi3Rrod18t
g7sWtXfPyYUTpeBQ8tYFcO90o22+MVgqUWPmRDCQALV8uZ14xXvJamwIwgt24niG
2VsDtKIT5uKgE385O+lzoKdIeDuHoyEDjkOiWCsJS1lZ+1r2XYnSt74fHdb7sjdp
fUcne5fcDfbTyMZyWlLyeYMkZv4cr8MevGizyqQOZYBBvwBLBpGKr3xxqFfV91Bk
TM77UoFAwPXnFE0Buaq5kH34UO7ST5KvvQCFsccQQi4PoueUJpPSexYMKeVV/u+n
RxU4SfjPzzexqnX6+MmbsNBuDm5p61km3po5F/Me6p1bavpTN9eU1XMZHBLBMs+u
PTC0EdRr22MN6e9Mcq6TcgwB3jBIuPgATCpHQ0KXa4jHqSIvxXOIV6cbXPo1CfGA
U6IbLs9lg296fef6YPEr9gV1E2ZxKA51xM7IfTFSKz1mgJ8CPzeaD2P9XMlYxC66
jai2eKADm/JKKKGPhpXni/qo4gjjSK3YEtVQ/qRJk46xKDnpCRA6/nlcwfheme8D
B6qCijf5xZX2ZJVrXWn1Ep+PhFFbFZ7CCInDu7LXlW8AC6CRewQubKmNLTfUbU3/
Gq1rQcv+yH+YsdV4Mqt2ExbsjBE/mWmmIDqjlT/dH2Klz0ad3URI1dx1rDl5kcME
hTnt3+sjN3YwimiTEpXzfuOsW+RhdU74TUwdcoFVr/5ozj4L2CJaj9FlN4Ytlfgs
pwE+iRAtK5V2ZEEo3FgaulxPjyzHm6oyN7MevmgOERL2AYn9q3+asfaWctqELfRp
xM5wp24QHhPFp89lT7F33OeNcL/pT4mPnj5mGFyR8bcS6wd60CbefZvwFWLCJeqt
JoarJ1RAm3654ch5gyFTZPepJKQY8RaL88HwO5fpsMCQDtJmM9RqVXvHdF3N0vHr
ewLerbroN9/nuLC3U7pte6+9bI3h19MkHrIWGcq/Rj4iz9yTVPEkobSmRXF+3Qc/
Sv9/+4RARC/6z2brMn+40cMt/OQjCbnQ1h0ayY+3N77g7mNwWtB2lptUPBzbzZrv
D9kborKgbhx+EDMmWYSOEFqS1AXkfJ2vt5Z4T+qhIczB6tFAPZmrV3Z0/AOpgVwk
CerithxxboVVizqfDHQW1CQE9qMOOV1rJ/tyASJAgzkL4M7be80+gmOI9XKzm7Tg
8P+R4nJMHgUvS5LbeqHJajRfzw3XbzS4g5R1tpEOZREu+52Vo7T/GAPMdLNcsNQI
DvkDcHtzxRZ2PcNDB6W8MkYP22YnAWuLN3PdKhxEtNI795Qber7jXOhSc5pdkQYF
zhGrEYj7yUtVu35GIK5y1rSF2/+SatBVQGcu6jj4qQYd/v37zsUTsx6xfP4TGb7m
4a9iqRZyXTkWIfojoOiWY3/nRhEe/5OTYBLnZ5YlCxNAk4xwDAfAXhCHJcDnUV74
XsSso++sNWN3j8KiTn1OMe5qUYzk+BgGuloXlykebAbK1WlmDCiYIau6hblliK0/
TahNzoD2Njl9q7sycV4+ZQatmrOHlU9IFQxfOViWyMMpxIJZ1RDBEItzJjs5f5Xr
Sy5+FnuQ5yz26Imjihhi9mTGpDQdkzcPZVprqHuUVa+wYA93Mml+keAjYrXszlVY
sPnIjcgdEgIBbK4VP12h0vinQ37v2A0NB3VNa4HdUJO6qL0omAz7onOhDAy11ZYA
2JtBn3sluV21NtDjICDCkToz9lDE+PFqOAkj9xXUaxKnt/sad2F/Q1N98jUjoxSB
KL/juto57ZzPcHE0ePAMLk0jHzG2D2gAqMa/ko83yrKn9yK+2goWcbAMlym3JH10
mUbJqpeeH8FCInTuJftijyvkZoIpmr+mPBamXxvvNCmifC4QZwhI/qBsJq92Gj6B
Lc8TkAiP+x9sNUBauqKNL3j+9zeYmzrSLbucsA1IktUjEj9DgW6BUEwkAKop7D/E
4m/zxjqlpQWpPLlGKKINdo0QmWyMiSXKMNDOM0TVAujRvviOueCiuSn3XaV8+Agx
j3naSVrExOhHE7YUiPTfy/Mp5F0Wpu09x2su7V4cTcTtr/zxwIZB8fZQbi3aAIOp
Isr+i296zk10k4nS+a1DecbFVQThWlnmmpDPPId4cY9MyoNDGo28mVd9H9xt5Gsm
oPDImL0ZNA3eYsJVZL9N43YIcfXZWoIvVwHCBmUpfj82IpY1ChzhFwHjzX45uAsz
1NFp/bIJyWOtvGR2lauCaZZvPVIX/9Vb+m0IfP7Dyph30aL8u2AiRDYN6Zt7akdK
2TB3MefB4NmvfTIbcBxWlql+Zku2OIL0Y7uI3uHSvnHb5ZNdrq2jt2eHLaZIxnFD
ywYD1r1+2dYmelprHrdaVFMeMX+Wu98h6UUWYoyrZg6ilNbzrsuQgueIjSAsQAmd
vP44v2uI9E+fonoeDpnRgexBEcYVea3jF4RoUO+CwT9rJm92UK7DUSNgMKjKYt0x
akVnDchPqSMND4QNqd1YtUwrFS30G9xuFR99zUyXmxzKP6Ij0fP7W9jH2D4SqDY9
/hkKVlCaMXFCp6U3l0H8bMdVak8zmIxuH5OtmbLPCp4Dxrdg7TjZqc+S8mIqeK+w
IT0jP3MjsN44iqCicNRkZGUqs2BcwOs7QTAvWQmp9ED0Z2j52VDk23o8XGXpbNHp
0eZc5OPyZhm2+PvYa6mFTgQhy1ojrKilHYxfvsJc3qWmQuetlD5PvcEtRz8q9Bfj
V9b+tGHGKXSCNJer1qKoUXrpkmXiVQyvVP1KbT8yfuvpFcMzsTFmPstYuXEHaA5Q
4giGxnXgs/EJZIQ3ppowH3fcVCZxnA1xT5FHj5Czo1eDW+4rmngavMEdacHr2xWV
07MeAFxixHHbPVjcmKlm1zyWXkUR0bAZsLc3Ch5NPMCDVRuls9cEk/ciFg4jSn8e
mnltQCwkwCiE0q7R8R+gCbNYtYQG4nldz2Hvvx/mnalXumPfucQBtPRLLh2Tg4PO
06KZY6qCTWIvKMBjfhTilW6nDoVFYWOOPiXt+9gKTdZoWexOg5EHAtdqespRTZE+
CS1jeFLlMRaKlqWrq5Vc/RyoTkfLe1NsUfObiPxQdD7nzdj+Em3VF5p0tF1MLcQ4
6gkMWJ5Vo49YzK5t7yq+70HQ5vBMieLtOmGqEz+bdybs+C1shmZmoGnmQI9h97I/
SLDs9wJSH8Nv/rfMSVhRMPws7a3GKfJ/lyjSA0lZMf3SQQDud+2pnmGyZYEy+poJ
8ixonGZLNzHQWT4Uc1YHOkQBzcUhbhykZix36Onxdnan11K59S9H1+5XdxIFrcfp
wrjYsCxegEaRoUjLOBklku8BElx8k8JbKlPdJTJVwC6MpRR/ZkdN+GI7I2pfVC3h
q8z7YR4AFMClvYaVwCeYEQJHFP/7hNCjovZyRP+UM15GxZHbV00g3w76asdbB/3z
MZnSBB2OjGuqycWMJWreU4MmFq5QsP27yRvCzQk55aqC7BKr6VLeCRDqldLmsSfl
kQXuIPzJp2Zm/24iLVWKpcNds4s9LdWTFq0MQXXvV6e0j+FuHANPD4VyYj9UgRXw
RVsQ2keL+8JMyO/nH/H9b4n7iWm8dzchKGSE9tIO2w+LTh5LAY67u256XaBlCdNh
7gH/6YqWEXDKqvzHlHuSrk5unxser8AGYlvUXUSTSYeW+Gs7+ubFG0pCMOmMw1QN
pjVbmMZ1Nlj3qdeVRvqNGyGBusTQgF7nMkWp1340syE3T1CrE9fQMYI08IWDct7j
2tlB1YqFtNMiRixMvklbRU8dr7mzlW7LMW831s3Jj/NcOFUvcPWZIFXhYGMqCtn4
L7B/XTrAawtBGkGXBOf/YRmn+UBvHD+2sCmBhCQSMqg8wANncRHc2wglhHQOXTaP
yLNRFEQY3riOm0kcG1LFaX2oV6GsFTj9Kp1lxOmOeiVIyapcjN+ripCNqPUqEruZ
epH0HwQGRjkZKBQWba+D1Dwn+5NtFcvx/6uwPExK1l04BOsqfrFTXzGHNKURKz5W
jkqVosBAyuOxaWJS7WC8QN+2/LADQInjVOO0aTYluX8FKL7EmEO7tG/b0IzJORs/
fC4uwopy/qYQ9ioheCxDRcFTn7SZlr//nIL4srz6kZd3iuNt4vIZHWth1o1UhHxU
`pragma protect end_protected
