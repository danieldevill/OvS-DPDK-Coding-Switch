// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:04 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jm1CKefjZ31SLv6wRPenS3NJqSD144nKZ7MHPLZ2uS21XNWIxZafPJxlSKh/LOHJ
47itSkBzDm+4NqHqzIazlmSCip6VJtCUBy5oJ5TnXd3+5ZlSOI7RrVzORrpjaNEU
qSdqVXk61wMeZR17zhpc1khwZTCiuRM2nucEM8D8LTQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13104)
2Jpd3wdFmG6l1f0wpw1XYYEf+X7IZKAMx8TCk27Lrkl5BIvOItKZ48it5X4rEcd9
mPNbvOHx40R99QmnOm/pqYjjcjQTr7sDwEQwpmdyrmLzeK8oVfT2dHhKpUJ9Wif4
KilwWVRx2HQPXuVo+ytMhQx/Ohgtor47YfbPcBspyv3UIh5XOhHqRYPRlPisnSvN
yWhz1b7h7PZVdJ2V+hJZRIq6BBCHiU10QiT3evLWHnlH2cSUiitesolB9qJjIyNj
nJhIDFtt2RoigWyrLZUN2iutAyI80yR7ap5IScVhpjNzRfpYiwTR5h1hQmZ0xhpW
39coN8/gAckK85VABCqJZUQvQDiTjL1q7/KWCIPx9lKXNd6V5vUCT3aNklLcmFLr
oCzWGKB6UdMUd8p0zUy9xg+TZUrxJkiG/fHxEeNsMu0sFCJ7wu56zjeRX1SppT7L
Gn/itICRsdZLXMwwqLe7A+m6MtVtI/hk7/A8TNfbt781s3zU4yppl9+oDILQDavG
xrq4BzXnX/xLc3Js2cSV2bp5R3TBEKKU4vU5gtAMmzbz5Eq/sFOTiv8xa0CoMYvN
LyRNW6TYMCE5vWVSbKBcuv7Up621lGepDlbS4A/G43/PULVnauyQn94IX7bLY0gG
c7+eNvAo4BE2JgaUsU0WsuXNHpWj5vsz7UTJIRbiQlK+8ZG+tgg589v2gugfm8dd
orS0Ez/Anv4ufGWb1BsmDiSvjdZtA14T6Rm/xDh/oxUZWadCo6G7YRSua7PcrZWt
QHvTOV0FytQhmZuzqA5lAS9etW5qMEQtLxsbfrzri6nV+0qT4bd/8mNIejaVR2Xj
PHpX95qnAfPnv7TEYvuNlCvC3JUSsFtY/1todYuEQfZW566wW9CA8hO2BfIExkqv
YtBgY3eOyK6vy+f9EmSckot+K6hxsAIv5yczUwIXJZ+0kpLCNRNyn73MRET51r+L
A5p9ibiPXIRbnx7DGqwtP4S0P1JJsOyhQ0uNlIbfqfv0ZlhJrjmvsP/xjwBvtPs8
pbm8r25l64Ztv0QPNaPf0prwzybhqCZ4ax/wMgtX0TzkZRjEaB1CH8aAgeXdIoWc
1U+ss4qSqgk2Da8tDROXrgkTTxkKZg3b1nVHVHqwvBTpU8x0FMKtLaNgsSiSeRyo
mLgQOBSC2eWpZGfZTwjmmV3gA6+KRV7XixvQW0ez4Pu6lDoEMbwvl/YP+Xqjy4H1
Swx6NrGtgGhNbg6yJEHyt+HxYNKIrCFQsGu+BcP5cYWLhDCqqT2Fy7rpoULhZp55
9lA6GHJiJTKMGYBI8XFz2DvaCB+sIx8ACnGX4Lrl7JOTBM5CloqBBc81QjFokEbM
0i9tIVUGhsNmyGa09oQaQXJ+i7RY2P6UJrqxDCu2BuJWIETmpcDwm/uH0BlpwhPx
ypZj2uYYQE7bHRzENYHlySq6E5aFRJiaOWlTsogd+MKoHg9YolX0rPFjljAX/2f5
yPoXJZKZXO+eSpSB9Kqczzh94/sAAg1jHFklmpyNQB8JKjrZAr+9/ibd35zWwUm6
IMsvItJY1V+cdGm2NHFI6/IfsSi5DqReip0g5FRYE8Zwfs/CBTAF+m59v1eAroPm
R/VNOztSxpOxFkU2r27I6aHYEzuxn8yVKUGvAFAtr+MvAUarLYCnPlheSCXEa9nt
gRAB5AuELOEWf6Jztj52i6njhzDIEBZjoR9GqNpD4AE/yM3hw0kX7y1zVYVD6Gxj
h2HAd78IsczDdVqZLPdB63+2m5WhcgvbnewES4gPoszlP9Dwg+6MKW2th+cgAD+z
tL8XUluLi3Z/fCPBOOw3NpmX6Ma9Z5I1k/6FRVRCIlr03cNyLSq8uDmFsAmdZP1y
cOpLxnQ+o29NxU9TooBN5m2pgCzFc8QKzHgzkJ31dMgoxKPoaawUgcXsPDAlcuB/
9qAVFACbyk0JcR+1bz64SNFzuCISL1BApBZvOQqRU+WaHAuJPJpfcVTt//orw5vH
wanUrxenP8N/iPG84pS8k2YHm1foeBEzvi6396a5OSn5C0gYVqlZjnDf0VpJEgUV
MNVqbB5CY8KyG2KtT3lwG6wE7O9ovnJd867QWVALjw3DaTdE0Bs6O3r1WtmUlZmi
UI7MuRIiz2y7s1tFSlluj7qC+r0VxpPjqNG56yScfGel7ALEFrpM0AxkP+A4XbTD
plpoBzBa5yEM/gEjtF4AR4Pbc98kcPDjnaxvLoftgIfRo5yBeOdPdMmW3b9eKcMc
6TnBTu4/uDX5IJFYUYVglcPJKn+NnSSODGUWydSiiI4c8XnIiQtrQjbpsVFR6ZLl
k3VAN/p4JZ/+njw3FmHhdj5LwmIs2BB61JwceegVG5zxzXj+qcJIn/S6lX1QBABv
EaMOIsBdZrYYFAzUDHNBd3fNnZGcPqAHS8NQTrK5IFMcBJkOFJxj7eq9T6cEE9XT
eCh/ukM5hNdiE4PfylYVAQXjpoLiSV+/7EfDmUT9ITbEuPUgBr7D/AshGJTcQsmo
GykgK26KwVxlsTFZuehiRiE9oc8x4/WH/I7+XW7/ygBhs7x2x9aSxCYQ65hNb5/f
iWqYoFdTpa8eIdi7axURM7h6AMzR9Fefs6VluMEQnfnvlY+nSieMScomyBRy1ikI
s6x6xXTwMKwdozXajE/vqjzfE0p0iY58qex0XUdPJv7BcxiWNpVzc8l+QWa6tO8w
MuW3WgaOquOvG0TpCG6Y4vs4iWWFL/0EbCxlNy59R7XVjQ+5/Awp2ZXB1ORkQZpx
oyfDyQzEezizOp/w7NtHhBK6VloRTp2OldK91jeRxq2vooMzcx6Vsco1zphgq0XU
zimHBKyF+wf7Yya/ern97I5haIsari7gHsB6VmUUAcruVOMGqHlsqMdk57mk14Cn
xOR0dUyYPF1kO94MJjVZPoQxDMch65hXZuVBQNRj5DdVVLsFDZq4N+CJdS2EkrHl
IYd0lA4W/gKmQKdnY4IDhVMCOdIDdK8PWLOyxncuxWdJeKNZEgaSECPMgoypwZ4E
8dAZW+Q9Y2qFSV3Ft9k2pnsFGX56cNLOmFQ6Zct0muzy2+Xcuxdv/oEVwDn5iWQk
L8yoDJddzJm6PdIDChExzf2RX6HDGf6awZ4ysvGCyeWC/XZPXfm7bEtetOBUywpe
70sXGJit2w+73+AEqDw2hIm/ypj43eIzW3O70iGGAb8bcMj1b4hYZobT9AwGVnEW
4NnaC9ii/M06PCjNAWV/tu5SHojFCOM34lynJMr2KFvCHCDzXrsHXmygDRQ9IP4L
pNu6zK4EnLC5mLMUYIRQI5l2RqMLSKjgDmsQyMKQ6TNjpmPXC9ul/mHEVHEATR5g
2xO3YeuAms2YRK4EjMlBuIAvWKsjSOHcRsOi7IkY1FB/8j3C9BtNC4N1iQibMVPG
jBQjhAKNWh3lgUND141LtkRvOH3wmRePl/wl1uDyli61fwBtxjqt4b2L8rM3rXJK
qv23+uurqvRbTZnCaPutBjjYNmS0b24bDYJsae4D3PfHI4us+Y2mRO73tzdlAGbs
uqyV/ppGBFPStyYC/xO9XPzoWWgtUmg0DYktjDkDzOUfk74Upt9Ki0xnO417GQgv
LzeH+Pu4lSlrwyd0+LMmJ4WR18QFw+dqlNvVFp/TSQIVf0Rc3dMM8fADBcCSUuJ4
yW7Mw7XEfS5rNfDaOOrXBzQIVRnYSN5nMXqnV2HOMv9Ami7adSHNyd1xnrYxSGwy
g+sfW3yzhnTWQC5gE0JahNOrQdJijO8TGB4mfZ1i3kKRwHcgiZcgMHClB5/5NVl/
+tiTmiTjKGLrQTpJLfTrmFMd40oLnMOK0VAvY7MdjmxeC5XfIt2vr/JyXCnMzd2D
NQQdKV3Y8BJBDGYN4+CyTU0uu3qZrKiaOy8lyrPqr621donUk3PuiwuJmMVYv3if
rYuGcj5Osp541/62V7wrvFZggeAI72W+TdcSa8TeqTwLm699mwFn7drweLLw2PLy
RHNJ94M0ADeWUNkAkjmRfm3gdg9PFlF+TZqIdSVLE0bH6f0XzGIPD0JDJ1LldPR6
D8XKWav1P9tI9L0bYzrSifaHXtDcB3aDcbqXlO8TnSXat5Y0thE9B4Q2IhX/nVBp
eD3MAyMbXHoJp0NR0eMWbvxjjRs+o1qhX6gYzXqhxXZRQzxUOe7F4VtcPKj7i7LE
VjkYKgVOuFmu3AcE+KYQ37/V7XpJ1xTuGAR/rkg74rwU3Cc/G7yKohKo3dWxQ2oC
yhE+VKQqT9VvOz7d+vYUVVLvx5MMb84YXilSVKizX4yrITGpnK6H7uA3XyXTfq7J
L1bADcScLPuAsEbuIUnG9lJp471ulFqIbbUiw/EFjB2Diqrmx9U13ovlam851LUu
tMu5zo/idNwGUD71lcc6B3cfTJEQ2aLWoXnBOMAUXQeSPM5hTQGVfEYl6htgVPVw
LqmpJ9xaAL3tUfpFkxaXET8wR1ZpEY3Jj1CbVfYoD43nVM+mxWUDkK2IYdDKmmAK
hwt+XFwoa4f4UGkVHvK/WcB73LIHq0ogul+NCkjaa3+UEx4pKcz+iatmfV+4AuQx
HNXHoeI3bJvmnWXyTd/ODe+wcRL6pZNKQ9syJFpMnGoIAJo+eWKF8UngxAFJfGjc
tytSo85rUcjEjlT2Xyg9JXdOfNXawxGVNP3ubiZ+PygVchC4szi6jFvd+8/s+MkE
Mw3+8uopib3ATw6mrzFmP9KpDzaWFHsXNQoWrnZzAbMJpWm6kdCo1VpXbtwSZSfQ
MF6cbSMbMm8DnFaYvanrs9OICjEjOETvr+ne6aEPRLBBcbRwmWkUmXeYwQcfCi1n
jAGC4EHtd6FpdHqbs5E8jSafxsmHlajLE7pzG3O4YCW9J0dLg/LlRJLGe9tls2fk
q0lj9S9M/lj26OnHOD14Ul7PyVtgU9zWqqDGVUNPE1l3a9pA51Cdu66ODVnZiCE7
+A3b5aa0Lz9Qn6gIT8Ab1khGAh50rIO6JfkSWm5oeVN2BH5zRvuygOlE3AZGsPB1
At54i71WV5woZ4mAVut2wjcN6Pej1kuFI7hVFCzcTYsQ2f548hWu0DZZdpzIInnV
YydqBDCHHu5P/GUkjZZUuV24IX7bfG3cSbW7MEmYOIzFfybqxkjr44w4jCbs4OAC
uFOGbFErW49Q7I3A2AuSdFhAeLF1kSz4VtjGnvvM/JWH6zeG/ftjqkEBSwG2/UrJ
LLNazizXEV/yL3O1Pvw156mw2aYvec3fcodnibmEZc01187zFlGF/ISVB/0pN3zn
1IPjX3WkL0OBKqAjmk5p4tFWZ4Dxh9ndotqR4izdzgecH7zL86vEnQLgzcS40sR7
QfmOmCRS0eKF6cjlTiT3rWGGVNxK5QAt4wMVJcZh9wZnunFHGDmeoWf7SetLSpt8
UKF6ul6KDgEoGplIaiX/xmckPZYKfMccCT+inzjSBbeweyJbgl52Tnd/W5NiTtcs
TTPCxF/5xCalEUkrP+UjRwT+Fecy8dOXvzwCRqkLnu031t5fc7rZ5y5I/rMo9Hwj
newZcUSveecFzjLnmWTBXr5bJBLm5JYuEzv3YhcTIdE0rMcg3WtghMwbgRC4Nftw
ozwla2Xdb+JTC3bBSQs736WiQ7q12bSVRMwIqSm0IiMEXa0z4wva78Yy60AE+g4n
FJg8fXly4mER5VXe9AS9Phwhebol0ebY7i8vpiNlEdrEvV3Vr09lezTPSb8hymu3
RPDTyeB1XVsutFO+A9VWjWRHP3kZ9aLQeWo6LbZxyXGLg0EEjl3Os3LRcVlapg3/
Qe2wCoKMUtjrpHhHSr4UTiecBzB8p8EmdN4m475bm9b3Kl79EwN3wah7ErwkB0Yb
zLYfblJYXFaQxTZXyJJIlfoDd8sAcMI7Igpwef8Ib88TOh+poFho08gCf3fE5g5a
E9wh2VL/AtXhX9M3OJqhfXf3LcK6+xzkJHitPHkQhAPsFByBsdWG34uuffzk1Lqv
/+2V348EZ3EuO295Rgc4jLnHVxSeFPFE5cAUlVUKuCap4RpViMCGyGbpxzej0M0i
ZUyeTvTfdUGpn+HM/7msRV6m7CNYqQ+32Owr6rYtfoaF3j/4alrKJ27G7f2LOk8a
dafyXjIruazpFL6maMrTc1qEoGB3WOiA3RcAYnRQuNzv7apWdtrBJeaYC2cudZt2
qbj1YF7joDh4T2aNglM4I8VlifocCHJ/rjncbZWxuy6qx52eEp2yBz0QmlmlLNni
FEa3vlWzY6+ECcji5PI+V+8Uioqhhc29QH0nt3GqdAtUo1Mk+lfWN14Z6oJI7Bh0
8pLsjn22IL6QLG2A6smIhslHJiDxO6zBtvHF69iD0guAXAr7//Hb2vBdUY0s+wL5
BNWwiZiiT9QJzIHUcdpu1TC0WEzP6h6ev/t9zouaEPDib7BEYZePOF8mg4zio8gn
CTwvV97HvOTntqwYPKEcTKx8S8MHeLEgWfNCzApYaX0arREhrsc2s4CKjQDGfZh8
1C9L6NVkiOZJNDiS4KxxKFZbMtsMKRnqkGDk9cc28oeyw5kZi0V3/vZYxTyrEuCc
umdT2h/irCF+t1EeK1CkVGfmnvm37TJjugRXTr51Yupi9Isg3Ycq9WCZywQhTuuQ
gEpE/rHtaIPd7vKj0RmhYCUlSr0NputtuaefHUOtzA4RVIqtii3TSWWp30NHoE7X
40yafx9MypU0l5uO/5nJPh80a73o5kCEI7BO/L7DJ0deXITEdO+y8VLOiGjI+Qxc
BPvogGnzBfw/yO5UUShsR2eLon2A+HPm4dsOJaTX+xKVpwmp6WWeQnn2mbgInTN7
ynPUr5RClI02djkyAMo11cFrkh7JmBhkHWUuMQy/77/4xxlkF1Q7YgZawOEyN313
iL+0/EiWd5VDZcMRY3k7Ht8/SY1Oq0Af8Wdi8PBpiNOM/JHsHZaJcoay8CIRn3rL
wRoyUcahYTEOk7ldxMx6j1WqO3jp18CEmAGV3Rr4Fp+R2p6npwXirjsMksw3ocPy
1FcLdZbL0LM+sRyd6VjXt97nX9Iz+Q82voCkRNYZG106XS8+s7vYm0j734JYiRra
Z4/IzbdxzcNl84oqRdqh1Aw/bew9HfiLAKujav50MHSvkEnsV5OwvcYh1k2G6sv4
UDfeqtD88Waf0VNbT52Sy44LL6ahzLXN7TUeOKs5eB4FVvNmHZ5QAYo9Yupfe9Bp
Kh26mxTD4OrJyKThbdHOjuNBFwGw6td0m+4hvVCpePgrTkvlQhhmjQcxFUbnH5Y2
PqbEODB7O2lKHDT6TpN+wpZClxRsaLOA2jLje5D9ak7aSmfd4VkHb0xtia/2ET/d
B/AIf8b+V50cB+HtUZHRCVj2oSLY8kl/L870sROQR7okt6/h7UXU4flcyxshjheH
ADUd0rFpunNZqsYSS5x7C/w2PaSG1sgDD4r5l3qnqN6s/o71oaZb24C2xbmEjDrU
fUbyMwwnLMJhSVgPc2Uo884zz+kJlDpS0nstJfY56RtMO2EwFO4KugN/iXx+emEc
JJ/6+wSD//a1H4EfckB3a1M1NBhuPDQYvkvHhD4S2LlIqgbi2VOLzBCju+8L5Q7d
DjD7Ca6fszkOy4imKGVlbHg1My4NvVUpexi6V3sIQ0qiaGcCVPX/0DmEx4Eu+xB9
sZiP8QsyR4LARZiob/VUXjawWFR+OedLFxLs6fLF11pu0mjJHKEZn8AV8kzjfjGP
EkFDPh1rez90kMwjOuKPUgVWZ81S46I99cUV9eORpsHNyu3y28GcI/6nukj8tb0C
qQg2hcZ46K3An4yxQ19LTTnmQSOPLzoDKJqORK4K460WesexMkBDjYVp5WENtxJ3
52cBw8d7lQL6jS+UgtuSKFnE50TcM9XaFEdNlHyhBwlLJBIv9glJAFbZWqAcjWI7
yE9/t6jFdHi0H+PJwF2vJLLhc2zHEikeirlMGKdv7aJ5rQLzq8S/A5qZc3Ebqjyo
TN2GN5FTaFu7+qazOA8n9Fev4nVbW8VZnlYkJknMRWLNxQtuWj7yzukwaWd9m/KA
Pc+A9Evb8J5NZNN53BiHRrIrzmA+TeAF4Q82MGmLNxc9lLiIg7tRCvmq3scZuDJe
e4ddrhbkiS01i9M6camx+MX35YEHdgRb28+JJSV3eNA4jwSyspBn46I4H/CegAoU
isgJDrgsC9IKAa8ek4N5Vm5mw1SNokVTgqxknY3vFI1+xZPB4gcyB9VbkDnBYgH+
H/EI14YS5KSVWsMfL3wPNpoLY+JrxfwI9VHQrSIGpzab2EK7H8rj7X+/pkqrlSBt
gTnagtXhVHpy4GmZVrFssoHnwFXghUi+V5icNQp1HF/yut6WiT4Yj/xPU1ZKG2K/
jFoXqPO3Af764Tvl4vRFxvJWjTzrDLRG2T77RTbiEGM1pb2HQfzq1/MqIXn9dF4d
8waZSXGlRzP/vOCIkS/zSLsxOEwKeTZX4F88Mimo1bA2VjvbqhHzCwS5jVMk1km/
KEpyLMWjkuwHs33h8s6VuZAKMuecMDuyituMJ2PYsb0FNEp0wjw41TYJq6IJuM58
M3fX1MQMUUEtiFShM9wTxjVxeksINDX7yPPfTvcTOJWRin2M0RT+x1tETQ9NNTvH
1qa30iErblfljGiWbfTFxq/PdkATaDVABAForUrzGvTQINcsw5W0XP/mhotvrFlb
VuZaf2dai0YdYRON4jvLw2wGEVRe3fXlpxU5hv3kW0sBd62TZCKInd5j3sQilfMd
B2cEp4a2NVUdWNFkN7gDg0HkkFcrXndRwHE+6Asl0U43+wdYstEBjkQrmxkjC8+1
5c8ALHBSk84wFwsg/mt+VqhBJouzR4t70JoS44yM/q1L0fllgYPojUlGucgemlbg
oVbwu/CSAmEzI6AhScHRJpA6WiC3RkBUWGiuPbU8xAFXb3qBXntd3WjT9cBpAkQ4
VpSBaCVK6G2PgLGx3xwu+uDXFkmeQSecP1Dty6FHbLpnky/j+vU16QBUiBHDzEPA
rWp1Rf0jnedLbyIpWc53f2TkuD7/nk9FzS06I9UqTj7O8eHiXvEQR1e0tjOoCNM9
v7AT6IWWdV3O5HpqCtOKQ3q2MIARPbXk6QPZRKzxLVj6dEjxfWRKdVmd27kD0v09
RpIcXzC+ZJ5XVuxT7z4/KB9GkP/oapWj4DwMI5WSMe95Un8GkdtyTZgeo5PdvhHq
bZAydrOp6bWcrtb+A2rzcMjhUx2hgBtI+BCu4Q2qk9xk0uYWSfsdg5vqwixWOT3Y
xrSfSwGJm+vlSPhfr4US/g3rca75tikVs0urCgcfkkmC+juzx232ObE+jgQA7GpT
iwehnhnrGv8Qlg8klx4xd4PH6Abrv3nM6JjyTPbqi+6Ctg94RxUXfWIKKZWXlP54
GBKaksKAx0OXoqt7MtDcOnPSWkrhCon/2Tdd0askq/mHfnkom2XNYZWQuQwU/ysg
UZUZzg8utuS/l3VZIACcwmd8R8iNwEshle29FyNMiO5eWE5+sk/oahpWEDn9j8Ei
RCc3quNUNjK6TDBtS3bUngHp0o6UbCrdWbmuWPmFjlAMPRI1+ccdcVWxNMMvtDn6
JUry8IJK/sSqAs5S7kpyowpUvzLSDC2H2U7DHVKTO+MZd2EalWCtSFpH//XwETFU
0yqaTKL1KD8Mtu5OpZXTNw3ywP/sXVQ0X4rClXnhAwbjF0uhqdtaCTcMVJFc6hWN
5UkDDmEwdSuJw3oZ2wiuvXLfX+jsk+q+X+KJOHvt1eUeJmrnlVeUS6LdRcYn0U72
DpKIxG9HravoyrN4zCYYFnqzfDNImnyf3BwTCWUvNuv6yWHrVDnH/M8v6ayco9+H
Vg4fb7FHQ0Ck2UId0Ba3I4LEz34KUS2nqwpw/9rRHbSZknf+rQK5+koisi5NExvM
Eo0SyrcY1OOnz06oCPQafd4dMZ+gTJf2TjcfEGUYZwjYJ/h28DhrSDrGuuwy71Tc
46FcMdvIKqOsZWNU76pj6wvjMbOqMUAy11HH0ad5+fDrb+lPAYrwQLIV9OEY8L0Y
AcHGh5LN5Nxayt3uostyfyLziURoCVsOUCyDNfi69IR5y4dks+UY4QOZLvipE0lC
41zjg5AZXwrvKtwpyj5mxBy3bCh7WRsi7YHaUZECMwv1UEKSr/7kKNVH1g92PxPF
RVbdC1Jc/rvU4x/POAvt2O8TAgD5JxhUxebJQrznx2TKiNUWnX7wqxOVMRgOuv3W
CRCQW1HcDGUlKdvRqeypXhUOazoqTr9ho8Iy7nvGSPnyatIitJTVQqP+K5AmeYUD
bPP0ZqHcwRR0RV8Cn8z0EzEB7bVByET+oL4uwMkNkPgDbDpNgQSaZI1fqzyH62qM
RVA6xty+mBnNGmAeNsnXC4bkQkaxapPHeiM1RQPfepEPc6q3IwfVrWERkdPi/p97
vNcLlAnZTZCWkzOCMC4C9m9Kh998jdwItxF3OcciA6DEpVZEllYjNv4K08U6Am9f
zdUhx9D7cdR0m0hrT9GUrvy5MmjD4TCxsCArpxqKxdAqGdkfcH6HRSUeZPIVbXWO
86QvTqlBkv5+yglz/UKVyVEgcDD1XCIF7ryf9mDD1xKYznS6BFN4r96+SODWmNU0
xFIImj3FCK1/u2HMVrgyhqggfc3etAre2bq6n7P1KLJKQXkMF2BR0ydekIi/h2qR
zyw6/id1hIf7x0RPzo1ZU82d/ZxO29wlxUwkJ1JhAFEN7nY+pGs4o3ZVe+Q46qrx
37HCMMjk3enKJuSbTUoZK+xCf1zRhdeXNBWDs34v86c1Hk3z5MIxvzxYoqlgkvKA
DpuXS3bx7fVvgeXRPB3f7IcS1iN9vlhAwObBMWtWFhCQcU3Q2b9mKlzwxNwLINhn
3Jr4oit06NYJ0AJfnC4tAT4D9fEP9UH1tsFrTWbmg9a7kQ03y140ai+lOavxUvTt
McUi6mP86I88UUbk1ZU6QNRuzL9+nSVlZLUImTOjdblMF5bdLedMYz41B+6x/p5f
H+Vb5bNYgaRuenJ2YKOBXwyMZRt/pgLfSOQCBLhnLVPeg6666T904xnZrl/H+GLJ
ZHLJ6/LWikbhusyWmHpSIBM0B7T+AX/oaY0N5b5fbKcx/njsj9+ph9ieGvTE/m1c
BcJK82syGz5waL5MdqEn2UKzNv2F6pqSO9XGeSJRQs7aSDruQ6Jn9U2KQLMCQMb9
NlDnWsZCF089t5AxoK3afkH4kkQTB0r4rzm8UJJKt8JvMiTAN9BYAZK+6JATNoX3
ra7P4ivaAWLYoXwJKjU0q8qJBKYyxRinF+wLxLyxbyrorFmzz23Gr9amwigkZKnA
GK2o7eH0BB1xvfcq42a7QYUDfgQrzagFZ1ttKTmr0AbX+KjbO0fy49o9vorjDPS0
/W9+QjKXkIhmF0UieeAPsV75A3+Q6I2s5D0ZIdQk3HtoFirlfGunNnPrupmDgvDZ
6tpj8hpDDKkxgjcUObctdc8a3uKPNdewXqNdQXtxJFyF8BcN3ikBOhnJm1VJyl3F
Sj6+ojnHhcso3gnZiT9JSsrOEUNLV6E6ZAniR8NIIh94TqOC7c44oEYfTx1mZifG
2zd//QQnjqzMhb5hS6T8IwcAxicUYyPGScPnIi40W8b6CsXj6miXwXySzBs+o8H3
euGloyY7Jf2Y/qc2eh0JqZuFVofmdnT4n7uIZbDI6o2cU3Pm/3bH1MYUupEmafJq
UAzep8HR/p2HMuiJSbZgtFPvLLQyTYxbcMxaQvDLbDSo4KtkphyT/zySUgwpKMDx
VYFep27HC1SbgNAr9mHsp4/moWdWj8rQtKcm07uzP580d+Z3OG0I1S96Lkvror1u
NzpfANHEpTdxxucnzkdZt2Zm+wgPhwWoPOii+aGKQZRiqCGkMk5HFO/KuFrNbg3N
6Gf2i+sq/3jlR19J3ryiZlvzBMv5Z7Js0dmDROctii5gPZx4FkAkCbUnD5YqSB8D
UxGtnJ3I2PH/pLNq7ftW089Ait1ZVRU5jZKfO1SmjoUhmejfHJUlEatHJNP9jFHg
PmUwCSBorqjAUtOqtrFGltnZkqnqVXnkkY1qwg40KchuURq+qMpIa5MOg28ZYjgH
Fzia8qJDCutJZlaZ99av5mEsBkvuKUB4b59dePM4Ux3XDTm+UV2yLGSpZdMMKK70
qbUpepZ/eF4e9yw7HDzPMf7rESZwI2SzaTmnVXwrt0EztfupUXEalbrFabiS1GoL
BYdyCFjGE2wV3m4gYnCxDe7xFHc3kQVxQxEqxDlVlKhX19QPPT+m+7FSCZHuWCP5
xlj7Es4GGwNSYPvdrn4WYYWbkcfuWxaF6O5SD98ionnBj4bNNonKr/RoU+Dea7dD
juSex6/lFn61AhJqQ/Q5al77qpJ6KppGKIbFmr9tn/pqWKzKktXR0LHhmFS9TG9g
jGEh254cBDUnVIESd+PVp83Wn72tw4ekYuLRw3pBlvVay7r75pCCXhMu20GbIO7D
o3soLrireylPwksAcn77krIYe5v9YYcF5owC8447k+H+2rXoZ4sidCjapOK0mlEz
ko57PBByYC/OfiLkPrqRyfA/1c8Nkfqeeph9PnNOrO2Qrmyw83TAztf1fk7t84x6
76XpJjMQN1fTS5ZK1RVxuass9ZNgGUVN0a4dKTwp7+k2Envr60pA+5jffHCL5Bij
mKimfeiQtOWchFKFSKbYs+/bshQuy+GpCRtkCtuqQrxM9+fvBlzniFJ/oo+G8Pb1
GrcKKVIvnFL0DyJrOaEkI9Su/leyKO0URnxsimP/WWx1f+qkqh4Pj803b207dcr5
B47cJ5flYUZr/4JO/lD7+tTuxrIb4csIHSiKraEnw3cYen3zc7uGj+vEV4VQ0AKg
SViJLU2gK2SDidQK0W9YVZ86V+fKVO+3uPcnH1FxwKbdXYvSyMXLx27/cLGV3N+Y
eGfKJo3x/PiLlGBiP5F8qyhFgzy2zjZ/fOW3z/RUMUffWKwZO6m1Dpo1vUrWLHg4
vG1/GbyKZaerKEpggFcN/jN/tcwVBljI2ZgIVDx65UgpPYG9IfDuFuYU5gqhPyB7
0CUZp39qwLh/qfoTBVFfas6TdbDtUYf/QHDNqiuZQjvPT3+wlkb+pJPod6u7Nc2/
DNVnSGHcINDtzjfMmSsF2pbuuRl8abuZWdb8TRHboTmVvwqwEIhLsM/+HBonIdHi
6NDbrX40/MawA+e5MpGqtX54L5NEQXWadEW3rjrTj6pBQKc3G2o4zvFbr8HQ8v1h
dvIiChf0mKKhiijWVKG3tOmIuOBN8dLB3kf2VFjT2dyJkKJU8twKoQX+kDSCWMcM
QigsARq42mcQ3XX4BPQ0VLrqbnjrf3136Slarky3ZKwHnh1knE7XrIrUfK02/cNH
RSjdkOrxUgdx3LwFCc6pttcprM/v0SRbbVlDzmLCQ+tP5XxmKjfwRJnlE44A7KAS
u4zF87ZQjFDffBwoG+KMqEN2hZnid7ywXqpEpwSEuaz3BlVKKAHzqRy6R0+Jr7um
noXdweR8p8gWYB87KAZBL5QLOxjnQ4tSoLAp2ZnZTqNTYs8B4tMpcC7h91m17JNv
xhO4M3dWig9ba+Ys/ydVqT+7wJMbNlQNCsGTEfnqP1FkPEFDZRmw0y7qASyRs+no
TtAypRiK1x0NF0ZiDmibleA1+W4k2mifWn8ufULk/oOppiIUAkjzvd32pnxZEHT/
adM0m0U3ICLNvlyH5nJiO7iZ4bTkzBWeZOdFSUj8IY1nVcEzKKRlA5e1SDLm6szD
4wBQo+fnFOJkkcX+UsYyCOTN3Ce03iz9LFjNsYcdhC751aiuH9MWmIayyVfThDIR
HcvGUn1iFhvJp4JQvmZPr6Tn3WnTrL53aWChNajLigHx7+boFOiW4Rmj5o5nIEYN
QI3I0CFyLz0w2OHK0l6cVoHb2cYg16OZzbqGO6yGpFwpsT+9ECFdtqEbNFvV8/C2
gW7ytahprlLkPHCaEVeS/zSCeXZ/GNe9ey0AqGSYFq08Frcx6K5TdpnPqQgzwsRf
1/jC3NLfSUSYfDQDSCBrmccEEpGao+ZI4W9J+Oi8scFlMUkurVmhYHd0vXDUeA9q
m0Fwvvmp3aZTdym+gn+7voet9duJ87ZWq7gbdvFf9F/Q5FkKvt5aubmZ5k7By75R
GA2g//dD4/Gs4RLh7owgDZdBA6VRtmNj1AthwodnBnk+9vXSWaWcLLUSjQdMcV9/
k14K6pi43hWSyqwXhvsRaqM90AHkBQWrsuyr/xx0lhQkLKd7X+EyMJMNJxzhkvnm
tuUE/2NBURNsaQVBRxYhwE578VF2Ns+NAkxyKejnXw/pjlew3AxDIFNXyYVgIY+H
Y8pOtlu4V3RWrkzm2N7TAXfjXAsLVrprXKyBZldX5H0zR/Mqz/v6a8LpAsVkBB35
GsFwk1frq5FZLbrIvOOE4Cujol+r3ByXlj5DsaAESlfWAi9GIBPxc+sxsxRuF5+k
u03Q+kWKyY5wV9TutCG0D1H6X9KI/tYZKKVHB9xUrWl8Kg3cYoe877xCeiXTctEp
YLwYtlWGv9Qmih3imvywWmAUdAl3qwM5dmtZ7WBBDPFXNm11NyUCFPDC6MgYBnv5
0M5wSRyX/aQGVs6DBLY27yjZV50+dq1mNMs/WCib3QdS15Jamf8iDh6kwVfWczY1
n0OQdir9Rs6lwmUse1e3xcSv8ipy0d9WObyQ0INLCJQX5HgOmq2fYsVLGQpSDtaL
pIy5PV6fP4wJaj7doLkB8YX7lHxsFdTMsG4DOqBO9Wf4EqMkxdj9meZu5l0Tmb/X
FNA51boNo9F1ums6vvMetd0IBVUq4NlxerOmdUsCo0iQdInRblWUNgCXnoBA+oN3
4Wn6AnZIfM0uYI8xvu6Lr5k+Mk/qhI4vz6Uw05OuqDiHSG/j8AWSOSDjpk90oE6p
8/QpBtjp2ZCtuh/rIjHRm8AeMlQ8/SVel2GpTa4ziq1br9qpoXUkslxzMncmWXnv
B4NOjCq7FQ6kYHtekIsENn4UXK8AiDgPrrIN2uofqlS3GJHh4wN/xJAOUI7yBFRD
FE4Ggl5zW/ZFgDai94JMXwbMdd0SCJiqsp5DAuLMXqiMfQjjUG0lAtXFFYR1ixp1
QZTvpJgi3lX5NChNe58Maysdi4dx0RsZlBWirH5OKWezZQd7JfKYQBdxifYkO42p
XZwC72ckeSsZGHhL4OXxzS46eQxe2vDmMrP5HudUwFPtqnz7dnLz0zHxH/atCcCL
x5jVVckvspGnKCMdS0IgQuC5BZ5rDrlb3CDmJDt9PNHl0gI/b5GGPOJZloNEcQmu
eL5nDn/yWNVVIWlccv0eWZ1ITZKawv0IVBuXsUN7RWEZwK/Q9x6rJxJKRMXcGZ7y
hN3aogE6JofX3N6wlWRVyFoIxcNbYShkTNfnmX0KjtLrOGzvVtleUwniYwRLUR4f
Zx58H2nLSnyoNQ8Ys3bEI6/rk4QI8Bz8U8suzljE4CCbl+cUfBiSxKNKZlcMml+M
z7Ajz+7GAJYWeEs6kV9uwR9XPitZ42TB2m15+l04uYlNBfWKVMd78fK5ab08E5EA
pDxB9ImEu06LWdvtSK/we7KbQsYvxeK+qZBhcV0HzrszCynqlLdGlu+LIXUPiYKa
6TowU50bSvRggW/h90MMv+JyX8QEeEZsHR03e/t/nYkHAW8aZHz1kiQROWpV6oJV
skLaP9v8z768OuSziEDvGKoHnO0CwleZ/QggIUcb6OBN0NELb5LV3X9P3uZK5X8s
ukVr+rvjGwivj1BGwjrdZrhpgp4pAAWS11Ix5J77aN/P8j0ppx3viFEKF0oeiGkV
EMQ+2MEtmiU6XJa0OuBhujcY40/0z0kf6E0iGL9zf9xmPq4FeRLFuHjzpyK07CYy
3wav8N1CZEizBicYjyrCapiQBch+irWrPAUEyh0UfHqLwbFcmolhjJ22NtsfMWoU
evq/DMyH5+Aghp1cxngbrZd0x0olMrEx5ig974JBslCqd5rxXQ8I3RRMkAAYB0EB
f0O58C9QWX4KE/iw4zP0ZdOtcAsEVTbD9KTY+DJ0FfpvG0q2HnFTGuutfoi5IRPN
aLRyiobbUje26hJtJiDJtmmOyzt2SsoRswH1klNswBAuBB7ReL+nG32q1/jfyaFN
B/SzGoAGVHkfTzQ3fiP5LU6cGvyADZbgVM48ixaI2k9U0H+NczhZOvzDKlBlxyc2
sUBYT7+X4LzOLaxzrrNuUZ1E2ExqUEJACik6XpHgrlHYDwMYx86FT5aIqBo4QpMR
n+qt/aFe0bI+36VQ5bzTDGuHxIDbo0hcMdgQMpoDLD59ooOJd8gZW2PKdSUpbzLL
JqYyCEcJHgAfuhvTA3MN67QZrW5EvRwV7C30SuXMbwsOXcPef9AyqwZpfC54FlzY
lXTPuZaCJ1YMerxFUKlg3XR6RuGF36iXlv1aZE94DmF8BE566eVsgQL0cUWNvGUf
8zc2+JkBIN/WxUjJLvRu9yI7xEI2CrOhpMlHF288m6PC3B3jq7GlPoQ80DluTsXY
u5UnTgtWh+sCtz7ohxyWlQ9c94TmdTlwqBLr1h++hiwvSSWBgQip2JQyZBQCVCwA
DgkZjB3tDUsF7m0y0wTvQKTHRa6jMMus6J/8PyLdZdmZUMvDbLy41ca15F84vnc0
xCohLe/aXkCtWitVr6jfM7MfhE4jf7oNg/BfZFo61tU88ORTAD7FTfsB587ntBbQ
cd8eyMvnFtISqe0lm2oO121Sm9loskaSOIWG/NeiljbhyueCt0BVBcxOYvB1lqv9
aX5V3voX6JYeIEHsXuGyvlLfy7kKaARw02tSnDObrDL8GjGmIcCp82dFoYUO+OYN
iIHSCjkIUuu1CQcrdBovM27mnA5hwb4U9fFWDKJkhukamPuOYHYHN9ZCUKFiS03+
G3XAghkmyxKH9N2scYizld5SFIod0IHhxUt+qyYDycgQl1nLgzH4opUFU9enhAvq
1NYcAagSh5LHZJXXWSkoDY4Fkipb0rfgcjI5Tx17yb/cOyKyC1rV88b+AY1ob9hg
AGV7fYlySqnBhjyFjkzzbA1EFyOr17b475GYX9uNochhxnnpFHbl2Md+yeQVqW54
hanZbgxrKxB3Kh4GlZz/fyfe2d7V6ovKbYDHK+fIzcimzJMLbasYueM/41x+fo3J
IzyTCCDUQjwNiGj53SiyCxUsniWbmwclAFjoAh1xCeEpaR5UtC9S7iTU2fw+lFn/
RJbGvSQczGPfe+iyy5Fw1AlXLUtw5LQfd6FXHr0pi7/nJV2gZCor24fvDUvmSb+S
5Y2s3o/wpxDYGmaSBifP9mTz9EdtHk+anXZgPqs3RL1aT9cyqAWQ+iVz2077iiMf
qJi4wr0skHLtDK3HEpdm4AbED12AZ+76jh1eXuA5wrFYpWoauoQrbQwq/gat3l9A
ZrDq9zu315x3onZ1LUhRdjCuijrwInPWaWwM/MENJvz1ipz9CVMFzHWZVa0nPc9/
VaCmZUEYyfsK8ka/cpZKLtRgg8TGvVMKCNL5hnS9BbZz0H0sMX4ntvEtg1GoRMXE
`pragma protect end_protected
