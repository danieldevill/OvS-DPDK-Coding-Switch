// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:34:47 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nhMB0cXtNoDw9Rhm3N6uhO2dW9tKwa/hnU9lBfmnMYYZ68nuZlRRB781+bWj2+rH
gsoRMoYq93K9f+XbOja1aEoG9h7l9WsxAfnX3aGGHnUwfHcr1yAOWt1fMMbDyQlX
j/PLlWnz/dCvitRCujBk8/ZA4hpjLyGNe5sjjQ5aUVg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3184)
UCkX3/ajV48t4Z14A6WzZMmJscTiv4tTTkZ98gbaTV912z3EB+RJvr1/CYqa88q1
MJx/RASHq73jji6w91E1H/LGWzu2Dw5czZOvvyNAa0UxBiulOHqqBEHBuH1atUdq
xoqTntMDnjH0xnHPH6fVoUnikyU4ep9tVRxSWTMrD3zzqRhBRguAp7YgtiEw07Qp
eEVgs04oGb8SutG7+EAF1nEeUyBAvZAJEc6d3NmpqGQ+cXnH9YadxeQGyz9G7V+g
kLiYQuOhvi6SgnsfZ6vAeMR9rnbSZbpKy2gvHvPXdSpKrQmP7MhTmG6eY/UteazJ
vtC1UAWrXfvKDYjwJnTLo8wzeMSq2XuozJ/2vsgmkqieZEWBFZIkS4VRG0vwnMhC
4ECc1ACKC03gJoJpSbS5GTSmPBjo5D+kuNkK1xtYOAbai90VU0264aVQBpfAqxEx
1u+26kJCGLKP6574VVeMw59JccmMKuMedrFbp6E6pMnZjouhk8LSg7rYgFE/rwVD
V02Gl5R3CJ8y9WLYfH966psN7pxW9YEKOpiAosQff5W4qg/BCeOWhTvXu/kJqSvA
JaY1rIMNYwXMmh9I43iQ66eLu0frDRcxTtGJrJd1+pHTyRYx/66cjr9DVGTcQ2t1
3CMhQrZKue1gpp+cEqhYSgcgDMnWyfCHm53PiHjjlIV1YYZsby/5Og5AsiMG3Uwu
dxEd7OwcJhIHfjsKKFxNM4V7cVpbSYpteBdF6yKCMhUp1yw2YzLzkVEk2Lc1icLG
cTkKeePoSaueLvm6k56CQslUQ+5HjIBzY+G3W5g0R8Q/rl3XXJsofyEj51MPSorJ
IaShp9Ok5t0KIGg0Z2etJJ/ndK+z1ykWT29aa6V+OSUCgygDpy0BaYPvzXNcPo0L
LOHyy5g1sLDGD0ag1tSFNlQCbqE1+gHSCKzsHj4+hFk1GXF4DYLXi2Il7w+GINgS
bG3S67XZoK5aesHxL6q1hhZN7FvLnsw0m5xFB7S4fIdwFzY7yDz07O8M6eQfcGNY
vRe5UUzdUD5v+ioQ5+PRv7z2lzFSimTqjprWL4uvajl+/vxpFOyjbNtdWLaxx2Gc
NARXVywBnDiHlztGkI0Ncw/2bK86GUjNONOW9q/PrQYkbqFbs1lGtfV9wuIaSU6b
ALYpGMoZUjcNpc6LFAzDYHJIJZUK7y+LxmMoMNZgF4r0IBPL0GASIGs0w/8kxzX8
/70rrNWNb7p7Aaf8IrBlhryXBnwQsxQOTN3bBm1eQ/BtVHXL9FxkUpPoQwGHUCC4
/+00lFyMGjtBk8pA6gdq9nDcT7MjF1zhUoYJSMfZ8SeD31lRhEyTvJsIa8OeLbwi
+XYkAhVu3aFI2qpCyMKXUnRCLzKToIq+bqZeMudwct2HJ0Ohtb/YN74DrooSjctL
M91mk82Q9kl6cTdo84+VawcTGUfQ6WSTi5TO3LThiw/bYNGZC93oQz9LO8WMhKa/
QW/d0879tlybUi3S/D0zTfhHzmhXodvVrlVHPLsSS2poHVBgegd8lymXIv8Lm0bZ
j1inEUzPix9AaYJcX1ZVM0DRrt9ESWDPV6TV+rFGyfzZRnplU2awQ6gO1y8h/Iyp
syquesuQpC3W67TfqgD5xbV1SGk1lbjgoEqRVTDIHrbA0WPU4J5oak6GoTsqRQhH
6F/eT3xBEOZXmTPsw97GfrFDHiQYUHgcobRAiEW02aoP8DNdGm6uQIsDlcnU7TSf
M4K7C3XCDJcHIvGlGMGuP19l/sN4c4iZ4lb/MTZcqy1jUFMZpkRC+dOM8Sp3ci6S
hKmKHsw2ffYLxyMalvyLVWjsW1T6g0LEy3zzzhMPpLXGrZcnBNU3oKk8LlGaMUQc
YEdKkIM+tUsj44MBZ3JYDOHEkfVgLj9KpMhLAMkwLIWKiCqqYlybP++AOQ0A4Z/0
uMxKFI4M4hcOnUeSTwMAWHv1QB5zJZPtC9QztzIFg+UWwFWYSurMzF0PK7Y8g6H0
zSAz1e4sah2GDmJ7elh6XvjyMCrtNQbmuSq9ZZPnc7IdMIQ8+j5TQ+oH8dJs+WBy
O6gxp8YtD2Wed+0y2LEbzrSmrC091WTceMk0u3VZCJZR8SZkrKVaki7zwf0OosBf
pERe/C7pJxEoA7BRWoIutd/KDizvQCXmigQgm1/Rw1AbndLoRy2B0clh68yDL39a
2AremOFH7oHxBWvwtK4DHLG+B20YvR2Yw9cuIUVyfwdV+84ia2rcursMZn2gUWDh
HEl2ThueWeiO+OBKMaaKXTVLxgIq89NchjWBIKD030I9RnZTnfyeCAsN6+QpapoZ
BqnQ9/ZurSZFPah92nQWoqrSCdTuKmrAE9VqBc7d4FNKImH05FSEBTSOYdJOEnoD
s2CCSrGD6aHbXHvVV8QTqsN3Eo3507XAmoaMlAZ2pMgv16EGTSK1OO03TJVNhnDu
Zu/iVnFlErQKQf+RqAu3XO/X7tWBh6+pfCi/yewTcRsop45PF8+/PLe+wZF9Pav6
0NtYWfSIVolKNPhmvKY0RNM9QwP3vykc5c2vl1F1ugkRCnOTZ5jmDzAkukWVFvRs
5oZhLU5R+5RvY1LwqFAKG/zETCpfjg+XLaor9t0y/d23gdWh9x/91iIPgmuqm0+J
4gEn2i29MOXxNcvEhTwO/TInZn+jTyQxmmVfuOW8i3R+OK0sO1nAEFfnfMwLEZkt
mzvhvTorQDOd/7EjzCqYI1ED2pfcyU3RSpuTQC6biiRC8JInyK7zkRN++UoQIIOr
jHKh8YYzNZCX0RnDL3KRyCWBqWtSBPBuV17ZdZaLdezLyyQ3DQq2a/h9qbFo8OS2
tw0GsU2uwNulXcTMcP+S+q22znaRhOXiULusugeSSn+ztDYc5aKF59aaw1/wgh61
nzvOGhLJrn3hR+AMRYr+rY4QGqy+4WnudqtfKZisOAOib41jwwbQFHbYT3zbPN7K
mWWLT44JRWCMTiyOF2e99jyF8ILciFWUqp4pXbikDfI2wOVrQKNV23/XD8yJJmIs
awQiGfU955jm0BCQnvxfGreXqxZgWSrmRKtqTr880Sny97flFbAj6kXHD5nfQ5v6
7g/I5k1quwvfclHbusnQ0A9HQFTUkNRjdlnlqSehkvaUrbRvkRvyYbAhnlGw/qec
1AMG/Ut4yOeRsr/tejd+o4UFHNHKpacNyIamQbKDr4dZSMGTNf/uKEppeoNTO6MW
SyIq+l2dJWnxoSn+8ER6YlyTejbDARLQSCuqhnFhMTC0PNkV2CBMr0YV81ym2GwC
9Uou85VhqIQ/KzMso2QGxNbUo0/i/ATgrWJcpef57zpA4WBSs3syabKPpbDJjNXL
kbE7s9qO7Mmll70JggWtKFwT7W43JlL2ivFZ4Fm039zx4WNk7s8FCUt7dSbhyJYD
rqmdxcioU5a3SZXnfODOEcQBIwjqAcT+JB9iI7VuBz/PV8F07CiMNGMZt56Kwv5J
hG0NS7oo2a/AwadiE4Z9fWn0TZcHAr6O06i+QCyEXzWh52alTUL6U3xiJL9SGqQU
n5+q1Ya0vgkI6OHxX94ZP1TvE15WYRe3KfCEZ4UegP2ZOyz934q2JuUaeZBQC0tk
oYEdBS1m7dF7vm0v1HEUt4PDYBieUMDYaLO+0yowUyHI82FrhzscprG/SwqTSXxG
ltnV/+NpgUJIeNbEPbTOtNhGVNr9OpqkapLNxl+fU0UKF3yhCfN4txCXscRwZ24w
nyqiBVz8MDTA4Cji+l93GubOIQepQDQ4aKZbXB3qzdGFon8+96VfytObOdOdnMPu
WM4LN9xcGmy0U0Z5gVXacCKOdPFUl9oB2Rdm93yGki2P/oGIokmmtTaTXlYvk/Sg
fq5StHbREjwFZayJG9N/yVfj3YYLwAk1pmJBhzD6cRfqkdLrXl7XGHbIpQpldn8u
MBx+582sfLHXPJN8K1IyMeRygeNmZRfXT/HyogZDMwA5NDQtjFyP+25COrdd4ciF
tKNttkljKSFKoAxMJtB82TzyKmelndenccYRp5GG+KSZL6r1XWFudvPnI75g7uX5
TnyO36Py618HKbAltV6vtiBMpXmmLDNxOhmS4VTlgJzsaBNjrNUVa4T5w8Y9l2Rx
RRy+XywOKk1xZ/9wGapqo1DQpu0HpWslufv7RCHWAXFOYl4ZcLjiRIWVEa6zduiQ
By8HYzrxhkeStrkoC6l6wgx3Ri0oYHYvNcNGGDD02FwPlEmbYhcIu6PfM6/3SHRM
sB439RxSKZSAIBxIh+rC5w==
`pragma protect end_protected
