// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:34:47 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A4YRfXmPsoqojwjxEiemNIt/Xid2K9a9797yyKQcIfPWDZ7NyL6nVzcmarimmTg+
bbToYB9o8GzHmgyNMlcOZ6RWz1zbz4veg8pLO4+S7DSv4E/kTrUvoesciHP3zROl
UnpKnYkn9f5Xci47DtPmZFU0ZnXv/KFN70qs+5tj8e4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7968)
qAB48VeTeT4Qoq6mSxN/fkHPn0p3+IYzwd5UWAwSafcpSX7epo6fBOYI7YoeaJtc
T1INnz924pC/ZWPTglO5VVliiP9uf5Dd+Vls8/yZMIROCJm0CWCVSMjVZbOiWEFG
TXs8fTqR9UchbJJOACOqX8/dZ3hWnjO6wFr0ev47Md+ft1fdYkdsIkfnrZjnNKJL
OfAyGPeLwa1rt4kDZC7/f7A5m3AZ/BV83ErG5/rAt08eS267ZjGDNTKe7qpyi9Z+
+TZeJw2kAHMWMU2y+k8LmcAIoK8u01Q21z0/AUb8m1KQphxbrECLLKCYl6F1CjZL
z0PG4CQrPefwb49wN8echrb2ZlcJKc04+pFtifhKK3csUa/P7Kl0E9ljppAuad0S
pgtKG26zfPXkvKg2tHPb4xOrayFfk2wRmVLaPiFA2rdmVw4jjF5gNwkhRqmVOaQA
Itwec1APq95PQK2h/HRBM4tFQ/OD6+5qIh3+vRJO9GuLC5Pcyd+1o9povGddo4UX
A5Rbj8q15ZVYzWZ5CEtpNDjbuZuLt5nYKdwaEU0qWa6NwJdUXW3h5I4M7v8ZvaIl
CLshKYJziImheYM8bZ8t0jsh3n5lq1SIWkBsbhCO4kuxaUvHnYl30cbb6c0n66lk
YXXB1G7lXn5Hvh5gWYPo5mCmyOK5pG3CAuFvQS3lfBB+QRWp1VZtixQO1KiURNrE
Hg/esrPFYw2SY777PJRijXYfuHcHUpkCwtJoBW7TbGhnVEb+XJl7plMCIheMhd0i
Yzec49UZNTXxpQZeOex6u8AIDFlrNfPGA2KJb3KRAPVD+0/c9SK07k1eArTALLu5
DFKYqhCV74JoO3IdrWBHVhazMAji+LTVkmF2/IPUBrieLjrtdZWPpudNCOxFM5qs
KenXMYxGldXbRcPbnnoVclwd104cmXCIvuxt7aicbdQvW08X91CfMlQoNHkkiFsS
CxqCyyJdADozKthq5c7E05PKJYZxNvuAnki/r/QwRi7iMNJOufnk+uAYYEgVESLB
aVdvmcpmyo4ElPB6Fg1OnLUbKXE8u4ABNUtrkNVvsGjQtGFNMGdqiKWJubJHhTJB
fgrjTpnWlyVYt6WqWHaSqWTxQ7J7z3AhNgobOD5zSf/GNb9ToNc5XKtls7E87C0m
cU1aI8fxPzHa046tOA4sx7H+7rVuyAu4QQhBZY81RDkrpl8/EAdF1Aryp4uWaVsr
uJMBVDC+BFZmKtuQelJnL+Tfg5dHIlkYruTsB5doBId5z7A9Q+/SJsILmMZ1vQXw
Yg2s25dvChebLUW+cd/o4BuYyCVcmeBPL/L4sfgI8AEqABhxTUDvUXPXOZ9xzdQN
yp1nXSPG9XdiSnCMcO0FU9oqvXuCon+B7CqbBPkEu6fAP9JTFsfFcOQqo/2lYPWZ
QlVUKZE64YmxdeE6VQyoKq7mICVUGLBaf6nU6N2+xQfIStjMEcI+d7g0IEJ7xCwh
3q6lc4ykrXFPA+UiZ+6lS1gK+OF8+1whkVEZszHOpvmZ0oknoPCjEsjByzi0GYzW
AA+oZHpnleQaAF6cquc8Sa++ywxERfjMepkuxxKHAkA1lRmWtc3MknSJsAbR1eIQ
buVc/+9vMmzFnVaVki+AP/NDAxJOwTQEFFVY/VyJcDpwZi3JrpOgDtQEjXc1ZAMu
iA70qo93GdtHXcraLcIPNykQjn53y/SUVqf9xqGQt5d9gIsqKL2VGEOGz33sV69v
l0tAOdUVOG/XpTDKnCICU9P2lkToFwY+Tswd8J2jLrxjBcOH+pr+0H7ypRcB75tq
Ponq8bGcAE61FJEe6U8vwiANP5KLAM5h6lVVRdoajOlCUh5mVnntbtbPbcMjqSwj
9/tZVBPBw84egIVpfit/tBo/gC2zs/ejz10W0ZDRkywMUD7s78jAZWsj/euscIys
Hj6fm6w2bvFqrzEcVQsSeiLxf+s7ZShSCZvhrwfCdqpNBgdkzXdv5TNnG5BF81Ih
5tEkV7Zto/990fo4v8tJPYmLYV+tMGNVrTYPaFuzGJVQdpyU+3AoLepAbEeHw3CR
RIV09zWFNeNLJS/eOsJ2Wu4UcftWF1ldNOCO/mihP1gRNpRaaj5ZAiOPPForsMGa
34u0XAe9jvCWvgRZgQWwdkrJDi8Fl1nNSHxoqlqcz2nX2pO+mLMn0YCorzn7SiB0
lt3LXQiYhz1yFTq2AaADS+U/MN+nHI4Tx6bLz2pjxYONKYzLMGN9s9W70LI25ixJ
k6bOSs4VYY7VnAbXrv46Wk+pqy7XJxBZc5oh3xPizqoGbW8p/VLMqWL5hGj7nAZA
tD5ESN885PCqajo/gJfeNceRMUdkOK4BlF0bCIIrjZACNXOz0k/MqiL2lAme/Rwr
W1y1Ugdj0ntoMeTNN4xHRsqNPI7QQnr4ctVWs03SOkUPhU53LgZ8JzP+eI06WC1c
uBEJBw5gh5wjPV+1JQ94BcXMHb2WQTpCx5Lk6hoEIkTw9Bjy7D5Jb5TNqBalHcdj
7ZEJMOVCuSgCIOlQRXun0S3TKhLQoy0BjS2AEUIiVBXN/1oxf9mph5fTJLxVDeH5
RTSPeJQAl1GU2ph/r6j6T9+YuZCTp78Awgtz0gjoxEGtLqp8xFwbPJ2+NfK9+AEm
2TKlyg5CwpLT4fsopUSdKhwrLjF3xZx3MAkqE6mAh9iIHbksWehZ6xhEwYmSjgdF
2i6I+N/5CLMdisxGeptuyL+ZJkE9O4DA8jKTBv1Mu2gnJZ1L8upFB8A78o1FzZoH
L+PCY3/d2082RbxxA56UpiATJywBuGRIJ72E3v+du9N7kApKQbzsUEUh6Gc+NThM
KpDrMgHURLi17jzm/C6obyAvCjDxNVvUi6v8DyXXl1XbQ/KLEv7AbOEJ3/KSEWdf
EB/HNNzy8GgLeGGezumFmKfIQYILuWH/kE3JItyw9GFZYx0HpcYrTxHQVbTqkPGo
OVthZaQsUabmt5nNejX/haxFULGrqPexYwTm8iFn+SVUZYUh6KPJ2UMHoevDq8fZ
zTyWuZ6e+dZ9gMJamDBB/t/KTZqg+60/98H+5O1XdA3d0HQo18Mib5J8xDBY6P+/
yUUf8O9VIwrm9LxEW86T12H7NSUEEuF+ZgERCXaxVy8eJ8N9pReJwezapuklubsw
X3XrbgOZiodyTbT3fjogEppVHTJlhCvJ8hzQkmG+J/kcxpnqRxCl6mARENdqdBAW
Jsx3X9vb1gxA6CDMOStJIHVN5/YRXfmlrzZnbLkTtVBTMBmPRER26Z/cTljwEa4X
P44J06/XDjMdnE5T++apx36TY1CN9ITt9fOmbrdq1cviehdUk/yVl0/sEk9V5mnu
/FwOkRSI4nLNT4AMJ9/QlnmCpfg9ECuR5mNh6VaCO15ggylouA7fNXp3NyQh8E1F
q506xuFJZRj6BB9rHHoTNy187QcpcEYOHEvDUg4E6vlnSkFFN/33M4H2HWIhX6Jw
0IwQJVZlTYlQuRWiK9vhHCkImoR9BTfrXkba72jwA9xxcw55qVEhSF5YS6UvGXmv
MqG5YuaqZ3dINJkKxjdBcEle9i9vBkXoXth41eKa1eE6VDIP7K5EkZUDXAV/gAY/
d3Z2GeU856wH2qDapqm6mylgDUVqZO1CriQble5WNDOvL7m1xwop/PhCCzJBumvs
TJs+xF/dr9jQtENsjOBNhJMx9FuhQteFEP5E2b7JnQlbPhrLhsNFlA6O25vB0ceT
KmBZxVNRxd+cAiQaZjKecQFEklvvm2cUGPyxEYA8PBPlikZ8rGoV6UmRUyd5Q/m0
8RR1G6inn/eZhcbH5ltdrj3Deq7m0CAJdQXpAWq/EHgcQY/VsL2AvYydnaS/gUQw
OfMWka1Ba0BScln+l47r+t+XgPWbxIk82wAtL8S6nKH0QDz58kXTDwJjk7tfEtb5
M/bYdEm4l6uVbThEGiCkGYZEY7cxBp5gbaf1nw/geNSeZ0uzoq239czeewTOCSbe
+kx0bGs3RiRZkHQ3uslCYQg9BUhI4xDu+mzPGIVAfm2FHzAdxyol+S3rwXdD97Bk
2ayFdemTHcXeNEz3QBp9XpAb6qShWbpn0vhCjHVFRtpKYXJow3hXdK7IkTIx/xQd
y7rb/K+bbaCMz8C+Vfz1CLtjJTYYcZ4hJAdT85g/f0OokGjihHzlo8ZRxAYKTX0t
GdBeQ9We3GutsOcMJClv9WGs0Cs8Sw3e9hOxWIxYbXigLyuiX3iLVv1Syc6RWHNx
3qbQ2iWfVe6ip5EjMpIuGJilGrZf+su2g0JY9Eb3UXZvzQjxuXd2bJ7Yc/ygkUqp
QRB7CymAjJa62M3QawD12PTpaCFlKpXbM85womJe2KjUTzlk/Km2CcsyTeraSpi0
ah5JGe5WM+Nh5iypycwXcyHMc7f60QyuT48Mztrfbag1I3kqb9LgQKlvsuz42t++
vT4ergzbdfFnX+NxAyggJFMZoMqS9xGUqLgxR/wrgDDu5l0fnOFt764dp6xDQQWt
lAQapqoKB49h1PicAu/ORKAwEgeH0gnFcq2qBn1/JCcfYNdsBtl/V3oMdefxNIlF
Eir30wT220ZgqPwQZkFDpvIYxiM792Tzam+up/2YMvVIXbqeLGbC63o1P5hEakgy
9JHYAhv1wFY2aRltGg6hLqnpx2WgsRGcnhY3qKdCDZIekh7Ghvpjsv6JX9tp2hto
7Ly3ty70ZuSAdtC08rsJxAknOK1CbOkjjOE1e82fJ3b1rK197TntoOfVl8bavWI8
HnX09nq8QsvXhOd0yQTRL+J77jcN4iuWTEUYDHUMBWds63ro2HqJEJ9GpWyWqLij
99qsQGYno/jIrxcHVXub3dCz9+E5YrBevZKYgxQrCraGSyxGW3g//Sr982jNvmjN
p5bZn8d2gWpI9cVLPkz7D48cwC8woqugQAV4FOWglAygHV9r5DdqNEnILCIxfwAE
eqG76cPJQ5f2FnhlKE1JKygwu8y6b+13uqr9VDVId1Dho0x6clH0C+3yD48ohh2J
2J8jbkw7ms83N0zW/Sfwg8xSS26jRD903wCRmO0BO2Q6H4wGHwL5H6P+kyd+WEwl
Z/2OU6+2dBYtOQspOI1XY8M/nIeeo90F3qLzObmolU4tCuvH1DZJ2Ft2LsS/Vmlt
ymMKv7kD2U6V4iiDM3NgdFl/2sDkByrc8yCbSVLt0zr+JhkF5A2hgmh8cMRiCNo6
2TRY84vR8og+rEseYoZLsaF5Cig9wVTCOlpQIDABMeJtxpVMB6XzxoAT2EshQDOI
K6vJbYIRqUEcuKp+mH0PfYxZi+dcMzhj71uwoIzwofYJD/bFLXormKzzRsdRtLGJ
QCUx8xhmIy9bWKouVrFoFH6kMTe06szCjp+ywMmCnxcewZ2VnjQnxUr6LI2O65CX
qFN7IMspVMppWmD8AiPKaEIn7x1WoTKuDM8B94o86GZZAm36WLWMH9s5pJmFIiN3
gerZ8RrGi0m5laKOSdTxyCoAP63YDVdIaZhTBOulQg1PngmahTieoofYeR9+vLt/
ZYQ2atinpqJpYk6Feii8qgunNZ1NxdXMd2VbhMK70G6gHz1krcy3f/TA4JOlwKg7
MU9Wul9LpBZtjDWC6arcp4o5J2G9KnUKwR1Y78PeuyRIY6qKm6MxsB7FizDPRRlM
ojPobJz4E4BCkJouyCAxgobyei0SnZtqG+w/8PUXEiC9HGb3c1kw0MW3q2cY7DzI
ys32lzrDTpkgJX35ZfDdYCde660OxI0OdGmQPqF6Xp5H0JmEiZ1HRozgaXIyOJ2m
aM6q7/sCHxl/NFm7t+Su/ArsytTOmZm8N9i7rtyFCO1i4MIQ2XDOE1wK27ISTrS8
xprjDvnxHEE7pV5XWQmh68wMxqSwBuEx5MNlUYJWWdFaCqAvo/be9DAw36nTTnUq
GzDcLfxgcJE2rNGW/X5td0CDEs4Lftkh0WNci+tH5pJVw6Ln3oaQHADOfsMvnd3l
7OTehFtPMLYWN2W3MnDT0vnzyM9TTIsyKKcwxGsg8HxzVE0GajzMmCAaPW98kmE4
xNG2qL1Yexark6NLDKoyhoSoeFrYWsoNaVDL6E0HumAX0/BG/t39Vk0o8pWeZqwM
uJe77j3RfrzXeizNLhxk0eInc6DFSzou7o2WyDj9fjoeIzX1RRu0JMk0tl3x5Gs8
6UTHhUDOa90wkU3lmC537LnFBmPWHBtNbJ6/kgK/PZxlKyRiEXfAxI7qY5lvUHIp
Z/JZNro4FrKAKvX3OGvhObp3DJ1uMclf6YKGp0f4pyjvsl5A3HCFxqvrUYdCyDQC
Cf7z53KpY5sFo71QE2EmMZi+5wRMMaDglyoXKZIKzGAM4PxeEge9IX8cMFwi1tbe
wvBZvX3+Wz3m0aPDLnJy/xNkHz2FkcldPTGA4Zjxm1TfghX5oLKxHD0JGNcLCJVX
61b9C40M5r1lcmrgv8TG2taEdDX+d24fPgRr3UQPwMSn3j1TBrCcYCJ20F61pNnw
ttY2BVnmBQptpTKX47nYTRCyyssyiv/OgOTPa+Bjk9KnfC06a4HhF93K06xHnlvn
2RPkLgzUr3/jiwvA16Jd++TAm1a0Yvb1MVoUA6jsUacQI+r6xXtCa6SdvM/ZqmHf
4ras4I5tgZ/HKcZjNxorgC6WHi3Tv9Ced/540L77MfMGYwncmnDaDPYPF8oT36jy
UsFd/5B8xbL4jrV/gqRECVYbakudfLpn9+NlnL8O9N0i6oxyV4SOFETt9kFtve4O
oBJm9NCyHgtLPvZx2ZV39XNcM6XrqGSjxUbFbxP7l9TK37hqJcpRNpRPpQ05CZ2P
uOpZDI63/ZgQ+rwnEFDeQkxILz0HvrkpMOEUmAZizgot1dN1iSrmwKPFSoJsbyzj
v1zUee/balOFJhuGuGuYMCKuJkSlGZwCYesppXmDLFSAzz8PfulFb+XqwP1uIxz9
kOd9QxbAuFEkG0JYIjxFNJDl/iX4w9qySE20IJlC8MPhgMMAP3BHYeTk8dyeqy+B
xRYcZZOG3hmvEqYCs3TNrHubvI2iyzq2silahbBBpy3VQPfRn+RfGLbhydfrQOLR
hrIBmEyx0vY3pBVdn0UATe2TCw7dNnAf/1glpBaMmZ7G6frE3gCVEw0fpiNaVXdu
XKDz6h3hAn36XCO4KUq+NOTNGJeTQOUHX7SwHxHWQ++ciSqSkPd5T4AXabCynzT1
XyFLhYqwHaItsUKPw0z468pHL9CULtaLVhFd2yb+VFPlwWgRcxr+cQnmT6LZ0iU7
KEMc27jr/2O3DG9HWfkTZ2iW1zTn2nnu0v0V8SipsVKlVrMIFqpDZIfiaFYmWyYF
zqKP7BNev/g6NtJXE3p13mz247K8Ey3/B3LOl0Y9kpn/cuGuL3UC2oQGtbSJyk4Z
JMaRyurNdqJ06N2DeF19bvUdMa0z+eRCjdn58bBDAWL1qi4Y5BgkTfhMl6ekqyo+
/C+tTsBxvQklw0+LhtkxxpBcUKArWs7OOAz6E+WOi/2WzCQ1zKiH+P1WBtVPP+Lm
rKTgy2wcCBAGr62zWMcLkyXOtx2frWWu5UtCFcE+3LnxJwQ9ivQ9U1EMfIOQNJNo
495jTMI3gwuyIcMjdz7AnlOuqNIaDI24XplEtErFRz7dpjUl/oTN8v1yOkVoZV1Y
Pm6DY0lb4UTKiwbmqTwNwRIcH6309eTUs27hQJnfrdmXtxMo1hVysjBwAGuLYbRZ
Vyws3XKuzbJ+upF/yTaGPb7Q6+EJlJLjg379uwZu52tP9nT3rOih5NwIF5Md6Hsn
wU4vs87Clbv32K9W8Qll0b4nxSUXhSK+0f0yVdhPwatL10SMNDHJAPD3MTPHfdh0
nKWXJwlM576tQnIBupYrKqE5ihLy/+3zK6V5B2W39o6FoRUpLUCPPCY2dtdV8L50
5Ft0qvih42Czv8MnnvsghrD9jJu2CqSmk0P8EhHgPIiaKqlBpGBYX/tVawB8YHuV
gvtzPPKz0/qS3UD3ZBV+Efmmfvh//QXqeFgAtV1UfU2pcKz01Dfb1s/na9+Mpo2f
wdsq3nC65d/aMKvoHFx61NH63DpLX/+Pg6NceLJ55II8mT2iX+iDLVSiwxwiE/W9
sR8q7LhEydgoj2qVVdnZKITRyJQuTXzg2HyNmKWGWAV6NwxZvpxfs4ykpbhZYLFo
iwh2LsmTR3mADpUZkvRBzTsUN+4CKO+vGlXufbodj1AWiyl2/rETdL3V2PWXEcNr
p7JBEypVzgPQ5SSgCckWwIcbyEvKA3rmXwMAxuVeslqS9pYKT/mZ21XPEPy240Cl
Pm5wruxwV2hqT2SWeacFwD6ezDa/mEJHNl88oPRD/B72gYm0vktIXctquq19fQgU
3HCwBEOCSghhxt/4lRk+h56ybNm9DG5nKqlIZTHIgrzDCHtMkWLerA8DXVi33swn
3V+7I+MKCmY4cjUd8U6AZUrRoxfUciRlBElVAUWGxoCk+lf4dOKKkPOl4u9uDPVV
zaxvQNp0tj/vVnJb59BctRDkVEyXxCf5tSk22hinaJKDL6saFmfrLIByO78d7y10
4q/CfffVTBA8bSzXkvE2wYCGKv1zO6rcaT17FKkcXNWKRReV1jlaQDyeTQOsF9bh
kYhjAUXQnTv7BPKfO2e6n5D2QFnI9EJ4Fp2dwOMWKrPWfqy0SR/KEpoBx0axkraB
Y4FdHrJHUB7pWJ5Tr4uj2qAMWLSIKnmqpK/Ktpv8yZl/dtHU/8A8gle6RVooz11L
pG17oGyCJ9okmfIhy1E+By9bcb1DYQLr5tXewtYP5cWSd0vDFxDQorTuOO5Ra43e
XfOBUZqo0H2SHSkfMVC8A4NBBMJW89L5Nf0D4iuutVP1N8UxkmBKZ0q/mS5yMU2V
uvWlW91EO2PztGpqCLtjvi8aRpPxxAJ301IvYMQGTn3gWgXN+LCnok1GOuEhA6yk
0blT9oTe5YH6lZvO2dE9gP2aBPAtqsKQxgAgSGv4OEv6bMtmfgMF/9MkVDOc2t2j
d2C3PCQTD2//ik0Saj5vUPUeYA91ro5fcLfclL5vp/UBbUlYGxIef1jdg6uAaPAS
ogN0CsVJfqLVHIeFc2ef7VpFOpB7FxFDs/eNmL+j9L4TUdVhvIFdeuflp4qMwY8o
0A4BGU2HPyhZtDOKTFjDHWuBDgPXsj80MFR/bFi7Rb/SVea5FQ3PzzNKn0G3g+1T
ju0Pep61rgEpkc8fnnV2X9fHhNsLly0dCBlV0XhdA/Azcsi/NzG1K6Qm8UhjRtx/
jzE/Cp10Y43YY53m2G9ulKUAtj//jeFrOye2hCp6fZeZIaA+FDnPdr2WkGubnmY6
gI3irGOXpFiYnTsLbf+HkpXhM8WGlgJC9HfOAlwE1ktBFyZOZa0PGfGrPb+sh3A8
YWeeTLAm9KnzEUZCtE68Jo2HZGAppuAizK0AVjyei1xoDNNHErydj6/LT0K4+lj7
sNxa7u7Z3rkCmWvRUUYoP6WqXXJNVNQzmsvGw6MG33DIfFclJv0LLN53PYrSNHaW
oOWc3zWCfZd5NhnAjskck7nWwgtelp3plVCTCcxoBTiSw8mCeSQO4d3jipRRVaUe
HDljabDincTMqVUfgTnf8jMdC9BGr9mRPWLkW7ChB3AbAj2IcRGX3JKdAm0sMiLn
X4IKVwufk45SlqxQ1TNQXYD8eFhEy7iiMcznrYCVzZOHSDh7P2MFL/91MUrj3qPT
qqJTBF9T5t25eSUYqmvYRGyFUU5BMFHjnuZf0nKi3PGIONPdB+kKGxyOrcpSquwf
hdlqBdhBAvUjHHUed/SvqUUUhVD7OILvH4CaTnjVkzrmkucc+xgotIiUqCwvF+eg
TJzuZkIEfloIEK0LPvNmmgQIzqkOaaGxeLoQS29BL4rYVNHo+/bFG3L1ZqwfXkgb
C5+sefL3fdH01JD3Bjywgc5kGJUfcP8EZZaMrOQ7+UdhTh/ilELIUh8KEuLcNSgb
Htz8qIPFFZphpXwtSLAKSp5VAz+G6WTS6dGIssu6lT/Nv91wc/RsA2wr2OAkfP00
8GA1+Q3UvLK/OHAhS+xy9Jijn1GjmUe9YPGqTIDOb52POAA+miBcQKLb9n75Jmnw
42J0BJjxHwgVXEYrypbgJGMUxtZZgMI++dgncMjQffg6g8geHu8mY9EdE8WY2Y1m
KlYnjQ8CHhtndVtReovcDDsEJAxcFefcGb2oRaP+1hd5/w1Mzgh4m4COav4XQRA/
hvWhxqLi6+snOAhU1fIUWlLKMSng+LdfQzlKx3fQT4DOLuzhSdh610IpxEEMEzAF
sGWtYyQ7N26h8ixQDq9Ivr9avxJO6emtnKj+/s8/XSb5Dzqffx1S5yzwi2tS42bK
bFVUVkcWWQdqv4sa0/rNm+CoCmvvwWkCOeDowiyWihxiIK/U3sg/kVEgAgPkcMpf
j5RVwiUEZPjWjOIJl1LxDbtAU7cqwEc4hA4ScgvMPGqWL5O7jTKlYCneclrUSBYE
9JXuU9bQAEufl266yObzUUWrRE2oYumlJGvXFGyLwwAE548zJituq0E6e39ku2vP
5xlTzJLbpCEDlnh07hqygaXULNrDv/+h7ua3BDpQ8Hl3K6VKitgPhVQh+o6W0lsQ
BIyKBsdcydzYwjWABgg5vZ/9WkZMDZY3HVX+jRo1u6kspgA4HBFqgwmzdEBgoYwd
`pragma protect end_protected
