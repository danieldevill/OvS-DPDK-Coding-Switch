// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
a/iFdiZ+6pOjoAniOIR0k0rpteMWlEatNi645n3manZ9jL3F+DWRuVaakzn3PwyY
b/KC1DUNsJ5QTfWYBnyELmXVuHygDpCdbqXtspXJE5D56k7PjVwHuAk9EPnO3/jW
9uWKaeVKxdqZ0b+b9v69PHze/evL3izir0NIZDn5za0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30144)
247ZaJn8+8mEUG+1X28z8JmMCjnhS36sCOgQcP96uGM3ZC7/PeJMKCMmRllMKMDH
ig0r4moUQJYyTlG2Ur8nxyvMquxpFUk7gTj5gAzvbWXUxeYMvOdBKuHjCFeC92NG
CaCyCHSV9XdwsWlY7AifgBO8PgzbeXH2L24vr4oAcJsWJioqVXARW7wo7xed5pDa
h6am2AbH4qpOy9Qv6sKNRJ5Brq+OcQ112tQq/yczYC7UZkuViRkSrDhnl5pOdgdn
/1PgwWDP1sQ3B8p07KKTwsOY3Ut7I2bldVUnEjJdxmouyxmmbV68y7JS/rttM+QV
mt6l3dxGVMj3zsCo0MIhP6XBq0Z/XNP7lV979CaEreSNWnUzIwJPdODXxnXhm7Qt
TYb0bZLp09Q7dKkbHIqR6av+R68r8A4qWhJldt/Ub1Bo8U4XVwoxzt15J7S/6KN6
SaTjNvGRRiMlaIAcARgQIF2c3hx2SIJCIBJ97xVCF1Zkz5M83y09NuEprZTI4CHN
HZe+MAsThBRX7shlslabnGk6zmrp8oTJo4+iUFNesJMRlVkT+QDzDr0Sljff0eFk
1jQLX4WzdTZQHd+1W2Zu/lrTHtBMgrF0gdq2UMGo6Obi8TbIyi43oz6T7LpGFcuR
dphLvfZtiKrUDYmYeE1+Op17cP4LnGoJsO6Wt2VyEEKnLXCoZCN974/vrGMzQaFl
KlmAqu2AK6EpAsERq+Pgr7W+T6hn2Yt7yNs/q6dUq9N4BwEOuh/RIAKCnFMEM2nF
S42HpRzeK0yopN3OPJSUuaDv9w3MZko2SMbW/LYU55uFVSb96Udb41EC4ohQ0Ev0
0TsF2QEBKRjH77lJq1UW9ToyQa0gO4oUdBNNjcL8as9T3d75JOtWD4Lc5Mbi6VaB
WUC1NJvVStr1CDbwGNXt5vTcbIooObkAV8AoAg8a8v6K2G30sGZvlunKHKNLQyDu
drbty8NwR0d5ZIs+jAJMFlO4Iz1x9p2cjlfHwCS5XCx0FFBQ9IL8cRHeCs/PkOl1
Q4hQEvSX6ZKrhkzip1fCFZ7iKr7khj9g67PTREZxF9/QxEoT3gWeJY0GERM5dzjr
h57jMOe28Zgqn3eRdLxgOqQEZW31OuD3uG0CR/inpx68UT1DJcv6PdkH/L8ahN5W
hB+OfKYwALDMjLTIjjGPBHPFFcPsSpKnub/u4rJjpzjRTt0OS371GsoC9gEx41ha
PKPxrtFN3y1TSyBRH38dSEQyrUA3Di5r8t/ZHTgMw8idbbcQRLtKiIYQiVovFCLu
3mNunv5WEM52ReDOA4F5Pm/CcE0MlZkd3NUP/o5K5J5VtZHj6A8kfsu1DqCYgp1e
wRDKBWo6adAO0LUAAXRfB3uUps2QHCqC9il2fllW6MAGHk1rHufBrpmsEzhQ60dM
zGYA4Zl9y7hORv+krpESkTHJqkV+BWP1EaH2k6XiKsYHHQx14/kKBV5b4uWCq//I
lTV/sgTLW2Ipn4PCASy2IUHIxUvhUdo+yg8jFcYdh0iSYHtvZlYUm26ykrTU0Qen
MmEPH8I8CjEOvtC5MDGvhEGGF6R8VMU+qdfu4rKDt2XLHBW1OYe9gBdtXuDZTfdZ
CS/VmqBMm6UHIS4YeRQ65CyEWfU/L4T+Fpm+LUZLx2yE3l4ZAnejuOIZaqffIJpN
KwE+X/Zc43gzZjp5bMDiZdfrCIn++kxcv2QBbiMg5/tVePffMGucUbTCcaHSe2LW
66WTjgDYzjkESqXza8P7lYzjkUuFswooYIHoIsdT7MqoWx+kZ2GEsSttfHHGmuja
7kPlMlk6M4FZZJKQJuy3gs4D0EZwWMH6mW8Y2iZw7tvAAjdoJLc1tDvITFrTu70V
AR7yaO/2L2Quh3S+thvP80eHf6obuB/UKZBmbH1C2o0ncI71jfFDJsFraisQquEv
v9kXStn+YQwm5wQq98Hc9IqJ2cBH3HCXGy3awHrLjqaY8sSXiu843V95Be3wQ5EZ
V1XmjkBSWiwjWOBsr0O+rgBLGCxoUt/2qxftk0u4NfldH65ZSE288fZvdpPSRwsC
d6O1A+Qn8pfQuK5yK++mxPMQGNXFDxPPksRtrd1GMC9/zOwURa8HXYlvnv+piU6i
hQGah/tiDmaWcH7McCRJsRPgxxbHFTGO9vJRDXJVVTYUU6/l/nJVpVr7OIZzqnWg
9Va8hNUWjMjmQyxDETWydh8EdbCkCgqQacSTZHh7RtYLZrSCSXy1P0JH7usM2VOH
mJBKbYF7yoKVJWQdIN0C/vrlUFSn12l1QxFme1nSVL1WwkgBCl3W7lzgg0fdLRLb
vujNi1ikxbTjeboodnoIk16yWpqGe5Oq3Pu9eKy1qWHx8CQmGCiCenhyNTlXLpcn
vFO6FctYzY/vz2zDaYbhpTZkMqyQDMxig16o5x1ltk5+CbOIBfCXeUFPKG4Uj4FQ
U9G5PMKE/aUx+PDyBi+uEmnJrmQNlHdaafNYjVrvK9XFIMyGuUeCVVNhjhfZa7yi
wvzKC2nNWUas2Q9V221WAFWB3H40rB/PToLJuzQh60t/Svk2VzhwCvf5RayoJx8f
3X6gJXWeDJGxmDZFBeiQL1MHJrAJ8bJ2VA8V4Mrh7+nVVgL04qEemLhoY8PSUa4c
6o83k8wcr0aTOs+9OkQRCJRvMTH6+G3NWCatyN1OBg2kgvejqWQVhTIJdGJY4Fig
Ntss8PQCNRZJrTafEzfWOWX7WICyZZHl3JSWb6lLjrvR/Zk1LKgsF9Y4Wsfd89/C
IvS13mexTRmzOtt43P+Lj888hHLyk/EbKWI0IPFO33OylliqdMLGSCncNmB8ovHb
KlYd+D6ixlyJXfuH3KparnVCWj/4yz2J4jyqxeZF8ECehjgu24at0Bjl4x7wx+EI
sYLgz14FYo4txV6w86qzQX/gMxyoRsnolWQvZ6aIgaFYlbc4Lj6j6JRvABYuL3PP
CgyXTMUB1N75vuyprgpg0QjtFojaGZexy1zTjUOBa8aMttTCckbkWXKzFDCN6mST
7+qQkdV4Gu5is+mNXtYuZI/1lOMzexLjGHQZ0fMKtu34hGZwBquycFRI0OTNc2XK
V9HvvRWR+Acr5Plh5acmauXUIPFUYTBX+lZQkhRmwjuFuNF3oX2mOrIF1pAfV40B
dzyQMSUudWpzuXO5DvN746Kv48XlOQE8l7P24a8K3HA4m9wimqZU+udmo/3pHx88
nbqLT49XnmskPEdRjSoG6HosWITL6H+G/FGQUrWKcSx53sof4m4Z1I3cpokjDnXz
Dh9iO5XIJ8Zs3FiVAATO8Dudspfcb2I4tonnSyWw0kuUIXiF5g6qkSFNEDudI9A3
CLGSMZhSW0bjHKb5KIgnOZd7iqJEXaLUWjFGrWLltawElEbDIb6qEJg6C1M8lOj4
WB6YVun3K6aR5RS3avI00q4bIchRrbnb9Ai/V61ZgHf92NPy8W+yrNwfmbic1RnY
Fe7C5ddzlcSWtjoZVtlWiUWNxIqc0mwONE7M021i2KZsL6/AO5dNRtELu0B33Iba
gkCM9cwW3Aaipu4zAt/QLMFlBLYbslnYBCXLag6EZcGUU6UniiTTpuhZJU/WkDV4
ZyQgog444cnk2IzhG3lBOSAyenRyXd4aBKGDJjdz/Rr48eWj1A6MSq3shoU3b6ye
8dIxBMQtta9BgTYWBERdVnHtV6W2QA7Osp4qiVIDxN38F52hg4N+5YFgP0UjNy6g
QulsvU/pPB+2MDa+bf2SuyGPXIhDyGEjCUYa93XXH1B2J+Tp1Ort6U00gceRwto/
c++Us5B9p8zpdAs2hthSAvc5LY/uqVpjOgEhmJlls5aGuAU/aV8zYaFPCfpyVOTG
F+jPXDJN0Ph0ZBxEpnIVoYiNlDSOZt3a9u6IQzwsY3+roh2nYf8c2bWjsCTDCPcJ
vStH6zcVT8K7Ip7gsf1YfK13g+dr4n+ZQYfC45q6+KIQd7sfwJN34nVr5j2Q9jDb
t9Dn0pwdqMOsVzjzGbF8+8vob52lD1vutB5HnNlfMJd+CYJzQ6UHUzZunhOe90LT
j/wTvOMLtCBqc/LFNIaEvoDkqszFrbBtUTfjKhtSYRWPP5NydaHZWDor/LdfnYz5
0x7A1fZB6xWF12hLU+NH16zLS6H4W0mysgDIJHbOIPE16ZFQyUu821W7OVu025tV
76yYm3/zOzwEki3gYBL7+qwIsC2I4LEphMftd29lW3na+l734AY923m0t7SBbSoJ
Irdh81c5P9RaewaabS8LLN9R/XHc+wy4/iqB1whYL/eivsvjqJAaiJn6FmCjqZHa
DHZxqCNoGd4UdnF08qdw5HM/tyudD9x+RE5SnuiT8YjWVO4gFms7P7UgwP4eaRDD
SWMo1uylgrtgiYZQkHWpWLSkX8nSnvD35zKgSatkZhxmJFi2hQiY4oR/6NUAucA2
jJTicbllng0pbDum8CdK4NEYEk54D6M3o9vrzDplpBZgYSYLT6QL7OsZ2Uay1kPD
phTXl8LzY3dkwP2XxjULTedvwLbdNWhSbgKyyZvRfbMvzAiVSKj/Gx7gWsXS0sa0
wVaVf4IpBqjNTdzs3zYKaxysEI4xdZAncazHZ1VoTnRPM0/vQC2TF5H+29QHsNLd
kfGlWy/brGqa2K+uWY1SYSJr9CSMvRJXBdhzXTR1NL6RVTKzxp32yWOZOFal7LYc
eaHRgrr8uQjyjNxi1Ep4Y9kwGQ/Fvo8IP/3KT+4es0g7CKrtPtrcT4orBwIQd08f
EF31snKboAMRDSGUWdhH7SVLIWnj1ZbZMOTOTp0DjRGbkxNa31h6xvoKxrX8DECt
63atrWXJAvY2CXocpiwSLNFISqLJnRSprtcLufeYTE1KKPLviHXakC6VJOwdWqxm
on+YavWeYLqpkzaVu6TdJd778BYD7KmJdud7ALoYARfEH1brSdUBWuFJbixMpCvd
YvHFj34hMbdVOhM1f0kLiA/laddxuTugnZRKk8SDo6yAx/Cy2aVGwRz3TV12pind
rZzt8GpnEefjU/NpW/112+Ze7MEGmyxaO12qnnHPDWeZvCK7E9sqNputB1l2rInj
S7RBGjAEfW9i/SxN8iI3yTolXJCCpCQ/v0jz98JtRptAwZJi/70wnvlcq1NhZW5D
zdsIN8+FSaqYmR/jhbNmoJu38dUPoVNfAK0LeMmdU/R0uRb8OKyHZXtU2zPNbhhY
3dIqLINBwwbLUHy6GDVLwhm/8VRX+JHacMR8x3fyBYbTnIlbAYEKqN8JT/3A73wP
BzqrsHQJb77rwP8xjbpe1GAu/d+fAjMfS6ltPg4gQfqdxe08NtNU7oeQy1p5QK41
38AIT7wleAunTgXs2S2ykQ0jQIWYr2pafmFc9XiDMNm81ZRH2iCaR6vSp9+TYBdR
34lJb9/Bem690O+pe2ovHD3CzI9lSy94od+vMvfFW/ScAxlJ2tqpqAebkG2TKOLr
emr82V+KnqScLOehbzpoyQof+vqy/6SMMcFzval26xsdUjLdcrSnNke5TxRMnEBd
kLbWkAZ19L7UiTZAYtChasJCg6U4JXbwo9+eQvk/rCoA88ll7bTeWbm7V8fosFxA
YhjaQvJtR3LbL+bowkqaHqizdzSX9PJCy+Lwy6LoFbRsCi3p5OP8pILxiBEztsox
/1HomQZ6BeeTMvg8xRLvug81dxrJ7r3A7UkIuE2KGnYBwSbA1rHN3AFm17pcdDKh
8BvBtncma9E0WqqnqjRMRX24e5dvRA2Nq/VyBNwLj+/XHBHbq0MSrkpX3onEF7/6
2v3TmeSHUATuIZKjdEdpOSFTPQdd1Kd8M3Jozic4JRimOQA3nzv9ansKWh77eiFp
DA/lOV0uiKoGHdw5966TrSDS0QRBsYsjY8xUuMoUOc1B9KSl5p7OtsgVRgN84wUn
288iPTPTRB9Iv6HBTeSVY9sWmg2KBb1C+6VS9yOuK8pZ7FGj+AGfgo2YmyRzxOTz
N7640AZp/oEzLbmCpDqJZxG54MRNIadwOL+f98MeFe0PCwcgTGM1cSdhoQhtZ9n8
mPzTXrU5n7+TQl02CnsBM2P9sWRxvms/2mVkYqz9nSzzliespz4O5CQYo/zE5c74
902Aihm/ta0X19lljLdAmPNPqhxfqhCEdm73qVZGPjiIQec/uC0FYx8Ap5aCBDU9
e7f2FAsF0yyzhK/lZoUNUUjLzmEpWIqUodIIk6JmNKBOs3leWptAC7nY4KDKBcQO
6fbwF+oppMLjVzKaEuRw6x5WTwOOYdrCt0YH1YkDQwAhjdyTzuUkqzA65Va8RPFO
k2mG2mO4P1GgO8lO9uawGw2PPNpyejjhiHs40GwUsJ4hfahbGUla6F/3VG7ilZJg
quVpDUrCudRyv8x0gQr1H9vGXo5rMb0nUQ2FtVM1u/YIkCa/kUSoXGi9pswQtSJO
tA5W3X33Z6AH3gO7aWsLbH+gB80EgGMe2UXPFFJyCF4XGxcP2f6b8undSqPa303q
GallKldFA9JRN9Px+3RjInV95/WOSO6XK0UVJjjt17xBi4ZnS2vgCQs8hA1TnSgl
9uPKgWJA718vXeyvA/TShsxQKK6JgtMUiKhYOf9Zsk0AUfMrMfoq2JwxWEEGyfUs
+XTvgmJ2s0hLIJXzXs6/fjYMMeg++DHuTvbxCMOd+2KSXXhVQe1I5lPm83NT1Yev
DXvgRHnR7Q5byU6jvveHHzVRe4vHyd7qjmgetkvYnU77UTnv3Uqa/c1VUlkxw2Nf
LL6kuinKH+ExpLJoGNTucoQaOlvXsexXdIuRoqtVRtHwUGmKdqsVcQLBV0bo20XU
dl1z9aALICPQ/GJmiUm32fHNdsho/2zM7XYGjnoHxTmpE+Arla/HGMJ74OULm2VU
CWIYUQbV5Z0mvSuKaNDGN0AcKctvXZxGQlrx7BPaun7SuKdEOOme37PTQNY3L6Cn
O1H3Y97nE/Ts3H67uuyXxfTKnIFbqzv2xPWFt4ZC6jPll4T6ocMIPvIPG1fnB6Ud
YAUJSNDSJgfVlIMwShvwBkbquCH57CY21Z8gfNfO4CXlq3awWsDPGeUoTrd5PL+Z
rSuGvpRenie/b4jDkVuZZJwQz2PIwGOntT2uS/SfOvszS9YSat4paFlAVr+w8QN3
jUJCRrgqjkIMDh/H2lUhGhATpDfpPzdyb6GocDa/tjx09MGGJ/3Llhj0kF1YnxzS
9XuB8DtB6llqI/OCfC1Fwx8sDLLdUW4+gHd1vBxkpVHpCn/YJELwcb/aTR4fDKbk
GqF2Ar/jgJ2t4GMPg0h0XnGXY5NL5fpCM7HkEmGeNjjs/mgMhdunRXwmJxZ6wl2b
EvwQLs8j0yWSoaT5zmuQ0vAjbW/H7N/mde3c2Jiwcmnz17DaWlIrmzUH2vs+FOJk
sJ7bmOHTdo/mDUjPJ7SroRLXp75muDRhgKyCn9Mlg8adbMRqH9vitlq6phu+ThKQ
6UCD2VW6zO08/NPYeZJ9Ab1vPtmEOxcTUr1ejwXcM5QWmNQYl09KIFEncEurGLKz
GNI2tEznAtrhlfeHDPywDl2JKYLFD3fJ9Dd0wwW0Hco443vmoZBoqsHYAS8mWBjT
aGRmOfd1CfxWwXIriUt6okw8U45T8QhdY0zCKXxd+OGaTw70dErqgGujOj7+pgqu
WyXbwFOiFip8VdsuRv9Fi6U55JCrO18SVPv8AxETxqzXTnRqkWiR/ezo2J5QFBhy
ioQo+1f80e2p4y0qC5c8JVCOy+lcdTKspiDQYTIV3fSKdOclamsPwgyekhgyTpnu
mnXfKmph/w9KhD3PmW885YvRcMVD3ARjVldmEB6t7V13PHjJqmJjLt9soCib4fhJ
PqOCexD6wKrThCVljFezBJs2DE1mT1jiQrzv21Z076xY2QzGeG55q9+GG8HdTrSY
aHLl5k94vJrH9dKuYI2znSSk+/LYUK8pZQEQMmwBhVlFwEcWDOH9SrYnK9wH8K7O
oPhdxhKravpNwoDtoLPSzXocZtu102VrPqwNx33fz9GU0kDkuf+Lrn9kfl7Ccylv
JIT7ZYOYW7QsdQfULUgEkQH6Tqp8avrcBiIkZzU0AJ3TbD1MJFlc2Zg4ArWIq4qj
xRcB3R3KgZgtxs2WTVWBuSwl48JrOKLC+WbdhGWj1fLqobIilevh20vWeM3e3SRt
7SHFNWu2iajEzBMBRA9oyZpWOChH3Z7ZZgB0sd586p8V556BlE81CglaPsWkOqRR
rxCEo8yEuixr6joOLGkHLvZlYBN4tSWwZPRyKgvFDG9VshSbiWu45YtrA4WBuqwL
Yd9lBOLt4rHVHoZQVxUul5i4mcDoN5os+YKCXYkix/pgojWBKJuckCrEl4ozWWcp
Dr/zxsHmxLGZEGkIkPE2J92VzJWc0BPmEbMIKuKcnZObxRGhnR/WaNR09OwccvHr
WzI7hZEHM0CDBYxpUWg0D5NpBzdBb3MSyldoBhv63YR3bY1xiWBfJrlmm2hC/YWq
hw1ovmsg5+H3vHylhIy5HnzxM5Tztjp+2JWrSI8r+0f3g1C+KIW6AKhZKE9/TM8i
32k20NGrVra/ms6vPvucaSCyqNjI9jke7Ov2kvtXGffBYRVWCMX4Ye4nmhdDZStg
BEzVCoHu1eDU6Sf2u47P/pHF8lU9We/kJDVsZIbc7kE+SrwxnrmA8QzYLpwPPIqX
9gN0fee7zhMOwXJDcbAmzQg6ZQG6Q9KoPh8ZdmMvHc10s3C/0O4FMxDWP++FXRhN
ryUtIWF6moEL1q6sO09IAoEXNN3559SGduzw+ihsXXmGc356hOuc9bPwDGVh+91+
cYtZa+io0QDWsmuf+MbpsvRxKMyj2cnVUhrtHcRQGZwyWCciDh6h9WtTfrjsH+2Q
xTRvffX8cVOKjh4tV1w9QCzybB1jdL0ngx69DkZzAc5FnPzJNxi7hQwROsh0nc0K
pon2AYuxbd7n6EadR1MwsnBVcTqGbapkf8v3plZlp6O/R6CE2x57Q8Yj3x1V1Zuq
o4GpZtlpTMN7/B9EJOb4lInEvKIP4/aN8DEPh+9OFVCicFEEZoOVpT2rq1DDe4d1
r3fYr3K+S1qkplWIoxWREVjtvs6tCWcNyOtkr2J6F8ksE/3KGi6PtuDfAn5tXi2b
1ikBZChKw0QB+XkvqnLoQM2IRAdlFAPK/Wa+QoXM6xdakjWEIZpb18NbuKDDbU99
mrX191d0W7vgGd9U3YmlEXxPIIXmnVpDU9ErJhdxWcSVsGfqRUe1d5hV1EJX9Jl6
5vcYs8d45k0SyAi4xNwG1XfB2n6eLbXjsK2fDFF5fox0mSYTMduHbg2k8TJ8ZU0x
weu0hHjvbULsJ7KY5BBGlV+BMVyClxWxunVhcHXT7efSsJVW15EkOcZt5UONxAA+
uOzltrHLD5vPG6F2DPJsN37Vho43hVehLMW0S/VFNt7MbjBjaBFOf4m7JD0/YipQ
P/8mZBA4gRplebFQQqzCn/T5iw4Xz3/uZfxXKJtScOjtTt3agoiRm2YKNy3EYgun
gdkOyn9wAX+ejaCbUmrOW3A/NU93enG/1LSZNcU+qnJc+qyGMMgWJ0k4pJ7l+xJ3
aAnJlaSK4wr+B2IyYgNBzf4MsU2GkQtduliWB50RjV2vtqPGbS09adjoEa2kccZ8
Gw0GxVSc9LtfgLuqOJgvEFvU1P30aLweNPyjOg12gkGr0PrQCJy1TZWypVpwc6bH
+NUYgXBrBnfZ17jj5n6ex18gBbEea4IcTxSBR4/eexTrP/jTVezcK9l6MwkJyZ4t
s6eZnNKR3MfyE8vyXaz3w4aQXtWDPiHPc8mcDvmIaRbZej0kbe57OisTSvWvCGOq
tPKFotLleRnxDVptiICId3v+akrCYX+MyB0nirQ2HMu+2+sQYTuO/QLjeXYzm8DY
7NyGtpY1+cbAwIZMkuj5tCeZmKF75kXrFZRu6rMVxVNP4pfpREAYnEni8hxC+zQS
XZxPBDrmNSGvbMJwHwwbMRyjPpaklMY0OHKriKpQ6M2+nYyJO4ASvrhNlSvb+xOb
/g/qRdrTqs+6ZdpVvAhpQHPXAb9/7CIL13fl3wvqmFhNZEeTW7dssgDROZNsFAos
4z9cKRM1cN0SNbZfQY2HfcKgu5tA7DAbC6V8HPqb7WO2pffLtnUA7rruqO1IScDG
5QHPBrxuOLrAy0bewuUyz2smvz5WiqtMWOJjQd3gR4nNWBSjqHFs8vHs2DB+Yd53
/ijz78sLSeI2UdJcapONig/U/Pojljs+6x9Nc7y5oOxbMDgidyFVAP7LDdIT0yNI
VxgidxF5WaqeWSN3OeGWrkPuzWYVhqixFe3KV2bER8IN8IrybXzdKPEfbO57d4Wd
P2HnYiSfbpck0r/s3AIMstvOUz1nIn+i0kRd+0afyl3tLQ0DVU5xU1s8MJKxQv7Y
0ouwnxDxgqM6nFHcn95cgcacIXwcjU69jtZmlC8ZxJe9c4BpGCywRCBA0hGAe+7W
jNnxTiRVyJM0v3ZJS4O7QgjK88WaCjSWHqO2NGAW7ZoJ2CFQrb+YTOsTO70h1LEd
3O8Bm5C1xKHa9G42e4bK3ZO5h1pmKO4LsuD9xRzRFCE60vJ8X8ZGqNV1dEtOfGFq
caEWVKeh92XHAVUM1Kr+9s3LqXD6zc+FZmHqEP2jyn4C2Ye6PbQnByVqx6NvxMPd
v08Ez630QHeXi6Da2en447h1+ZiIQ76PswvQIUR9rRhtJMcisz48+2oY57tKb14P
u6Xm6lA34Qu2d7H2W6gqxATwOqZUA7gCvRFRiUfR8GDVsmxFVkuuDAZ61I9vsaua
zeWoGRPxf8vn65gZi3kGluGa5LDtrPTOahwg4gq+EX0QC+zdSbSodEg9roBPRQyx
6nUZEPR1IWtUXiTC1dfYqi2vqfr+bLlMlibErT0MH8FhfDTTjqKyhwjVbM9B1I7D
2IzmVoQN3/9OWiDKcAjkXKdgbQEtWpeNeNqA6zTS7R1iWV431UadzjwhIvV5sxbw
SOCFFUJDGnzm0LtBcYri8Khyy8GT0ZAPUi8NwYaz9w8s5k5Q0u4tJ8ca9qQ/Ezp0
l6UmC4cy8P8fiFSqcKZyxdPYoNYPlYtQEQ83jFYZkgTeP4bep60DIPpYtUsquhFR
b0ul8eYpWywioNYgz5qloazulWs9b2+ylPrSwt7/fL5nmg6vMM7q34cnf1UEcIt3
93rxtRNpj0Y6+m0sew4Jy1Od3a/vpFTVt+GN2+CTtK0ox7e1xOUVc4Ni/XMe0DmX
yu2O8tDy0Z6aeuMtCVnMnwgRfzOLKAqYE9BS0lyWX7/Lzw5hOGpAWipIQPisat9q
1+0HJAdJEqibMYucJT34okHN5kqALKu9PMiWjGz5OAqkB1D2X1uz1lOFy5AV6/se
k3kSo6vZ4Uc4p6ZWCFyiKg880hyUWt+Y6VBPwysNOFB6TxOw7ezB7iZdlDNi28s2
eW9tN+18OcSqbI7uQQM9yPE5EaxZxMvNPrWRdZ3H+SwFzZLcykrwB9hl5WGyZPe4
+1ADg5Q+sYy3ABjg6XHUBFjZwiFnZsXJo/1XEmS3eTl3bHEi7tRHwI6SRrNhv1Uf
wXG6oSe5+FcGFIpflfVhABCg0nfu7E7cYiWmNN/cw6nzhfMu5C64vhwl46ryg1+H
jOiU1kZCOFJ/FUmvggR+8TGNV4eVMkVuVrmCKhtXnLNgvyN/1Gv3r9DOibZGsRHr
z08iUKUU0vHXC0iB3K7hP/GYfmalv0ndJjOyfaZ9c3AewjOGxUyQsDPxNPkDu4Cw
PoqKvh5WwhuCYZfDm6PhdovyX5MVCI3i+0Em2NK8jkWpnf22BSyBKprGOaNmWOeF
gIud+/x3/EhfPA8KHfdYZWmnl3xxXbAAEtp/I9MlvG7eiL0+chlpm7cRMdvzTCJA
PSlzml5bzbFwmur+xl5rXS4/DwM/HDT7iWgt78wC+IXlBALPRbEz2ict/Kw0dYPv
n6a8V3jEq72e7d9v50x8jSjGbttOAVru4So225VgFFL+zx3PRU6klnIaeHvFu3xx
N8RQzIKmcx1FKpw5DMJKR5Uo2aGlvkfEiGj0Eb1omKwMsIMN6S5qQ4UWhyMbogFI
SQPjp00TbS5XCRcOFttQPFQRYrQDzn4znlHmNv5JmMzTyYpTjDP4TQ6F/8dvZRvn
JrIPSsIcG7WSmrFRwjcl3/0wEvkHwFVAetgpr+evg3onVVp87WINNUfTaLy5t7Mv
/n7WWYUjx96T0u9xhiT1Vr1aqWqTMm3zGCTbMZQ2OFcOlwTYJbSR38kLhnq78sub
odNG9F9CYXBarIr/Jkt8BB4/GoSUh89haCCmxUZVi8I7rieH5iji08Fxprh9Gmea
UDmYlJpDjWDKYF9JRJQ6QLSTEirP2dmbfXRNIksRpOdMTm5RZw64V6myaqVv+KHh
9gfBQXZJEeNmHrDrETtb8Ux/s0AQkbSamWKW/DpCoTMriuyykfzGwd/Ll4O9p8BR
Zbo82V8x6cinaQ7rqkZEn4+vKqH15kDZqMRpPWJyIh+q/9083PhAQVoowhbL2OMw
nwvv3NVYj4XdMsG/VjfqwMIMIbF5cw9TZlHpgGSxd82B7lE/3YJ7L0V1bxhxeITL
34JCuy7u1xLceVmLHGXO77AUnh2jgVS1s6ggcUyQyhLyUj1fYchhtPQ79ngXtCUv
k0mQEkx1cP0coqrthPs2FGhMdsiXFR1P+NhkxcCe0Z8GAYP3wuN/q2vCLpz5TGbm
AteQJltEGkcwJVFBPGCHsp9EaCN3apwO5uAY9QkP7uQdSdKS2fKwx9F6TOtQiYES
PM/mjie98HiRCN7rXy3ykrp2kDqGdtkhBRWFiJC85d3vD5kT5yiW5BfzpSj3JpYh
WwMkK+7l5VKk4eKI8rBwbXyCID2pTvIou/hbgMZrjL8khjSKsFa4Nc7yzNg50xv1
qI/AXVxNLlldrwuLLWViBxeiSE2Yen+AjSeqfJ72zJdXj/AGde6ciX1XFYNc8ejZ
c317u4x4c6aIvNLu5xbq/nyVshD2HeJr8Fyd0uilucqq5XkT+KMfzGPOgnO8uZDB
pUadEIUYRfGrZJRSNSHqpAvOrkwcqoJ3WimcEFPsjNHOfL0RYibOJdPl0rthdSI5
x7hpA4RBp6WXunKMMR7Vt5NNf7jdP4Yjzd4aQgjvae+RgXcKgj1jGYa96/Z0dJ6a
5/AwBMxUVIJXZWaX8Miqp+WTDkkWml2pWEwburcQ/4LLKJ/Phb8T+oNP13QBCaci
s3o6yGbEN77awUxG2e8M6PXSfzQJEakQgbfcRNEn8fCRj25P81fk8m3+c3OVJgrz
U6C/KI562jYdY3Oz7wmLRP999HaoMOMy0Kzf0Z3sB3cTgAFb6rGtiMTthbteh69H
D5EHEfuoYrSiGQBrpgueRGRvti8B57RbpdVLsWz8u6dqiIyHl82ihGXV6hJ4DBvZ
kX7/vV98X9PFlI6wJE6Q/2FPqec//uw9S6kk0nW5t8/THmaVTvXJDW0B45DiFuVt
MXytuVQBKMD7XHqx+atkjmvUGdFVXwkExUMtEkiFYBNLVqWC+3lT1ztmxlggdjo6
OJtuiXVhiO8MI3bxa6M1CDFk8J7CHjT20HHKgBr31mFg2+VzdoYDTTfQH7ImTJR6
GfKRrn6oq2jV5lxerBmrOFChAzZMkHKec71GVMeclLTOMtN4O0/YKqRwy0ypf20i
aObdKt9nvOSsROTl0v+2J3pzllogM/n2LWYoD3Y6g75zQcl0xi1qN/cwqR+X188+
JzbaNE+dF6IOM1eS7yU+V+bGWEaUlJMck7vBchfb3gUiWTKFoWaAMVoKdGvOa1KV
XYucsXKcBA9S/4gQeM0eW+VwBiA1hb2k3kYJNDru6Dt0o7RbxapSyqN/lulGppRK
UeLwP+yzkFusIoutRyTOjH1f0I1WTRp0KWPMvx3RHxJ8VbX/XulENnQFzLobZubk
dEB7LJX8vdycAz7LdAtS0FTmmiYHxii02QUyqpxCYpZnu2ZS8u3c5yX1f3MI5BCE
sgF0uMJ3M/FRu52CM3nfCzN3KcldNBy1ED8idbUr1gZFGnKDdRumENWqUhI3UZ5s
NgOmRtRw7xEmdipa6AzGcaoU7xNkt6eK1CBqAe+yI/Zy61SWpowdknvtItCiZpGO
N8sECUOw4Ovj/X5eYPJYp8Coee+T50rvfOMFjD74BsB5MxB1TJXOl89DZB8iAVU7
d0+zukXRq9AU258xHJVvMpOZ06A0dnVUnriSgDt3dxfPkRYalBzKEv1IxWPkF6SX
8uTou18u9ViOYUyhnvbGPSyJmuHbLAuYuIJOgLWmvkdm7uQQDN3Howq4Y/vE7RRH
YXDHYXk9fK0/MMzkaQcxfrhP+2xqhuUaZ5QgmAbtXM3ENkutSd4/sL3WA1GkeJvI
ker22dfEXefJuhksqOz/50RWCl95wpHI60B0Ie6Y7rrzJ+YxEQKg5Kc0TLv4eE2r
yjOkmuQFNPi8GWW87bVvN2EbA+IY5PhNzefA9gkEQQwikRLqx8OtbYI0p4SWF6hQ
9vSDEA83mWhf0tRtBdzEyDddNEsrwpjXG70YH9tQWsGMVi+RJ2DUDhXEnZEropdO
z/iOm/Jt6lyefKGRCFRDtIRaz9vABor1cxqYwHZDEVFw351/g4ZLMaBlTPBOwb8s
Ug2kXFqYdLTyYn6RevNeAhSfnBiFJFYrtmdyCKgAvFd3LJRp1pSKSt5gPKgohxFt
mguKSA0siQpHg4iL8a56tOsxarAp2PqMw0OYNY7i2EURfHeI8s7r8O8ctGCS+wHN
FiIPFYIueFcpxz33CBm58XTR8FfrcJj05Oh+GCSzDlkKgO4WY8dJteeIhy9HLazo
9l783nbL3WFjEK4Hbn2UXY8ggAJRS46f4ObB4IcPxgvI+qfBWYgbzxOiFxeAVeRk
V4rBGBPsVq2+kbnU2vyWUOu2vOfjFRUHwtqLzUfhvXrEIMsogLlFTNwJLxrpav/0
thYXcmckuAQoWVMV1lywq+9xsR/6eC90oBQQ0pqmyi/YohXb3FPyBAqsjdQsZ112
q7cqSJdAqKRoGV2JW9DokxVYKPWw5W1PRdLBLYq4qhWZCCJ8tJ/xdo74xCKNu8RP
jIbRxwA3JAeIBHWqLTkq3or/Uo19vISru3rJD+5tEYCJfrSX0uW9xnfRo7xDurFz
zhwDSjRHlLpsDoUUUS/MqqQP5W9D7Kh03dxbiEEVP3BGz5mHoaCfMER1ZKpUKNj0
7i2D9M1I1BaUKJanlVAfL377tF1ojYWynQMM1Pr6R4J75A3UAjYJzrPcUbSylIqP
mQc79hL0PKjlXdD46EuAhOKkIoqywD5PfunL/SnUQ0e+L2TR87bI2DzaeBUslaSB
GzmBYcXkuGZgkF1IYHBnhoBfSd9IgBRy4cYBNXpE/ZQmOhtQ699Htqf9lvOizdWM
gkqCEdpV23KdYiLZVvph5OFZttZm3jflqi3uPDHdissBdaVs2VT23HzjAV4J/H6p
xR1OrY8bCLoTQNEpwTO0Jtbh5QQaQA7s1WckEkbFBtOgMWiKGOuncxjF4I3H/BzR
UeCyAUb2XhtjgpX2J2mpi/nCvWDaDy6351Mo6SSqIMPQZ41kvP6+1DZCNz6cIRGv
zwaEcQedtX+cQynJ3prLkenawUt2zLeCzJSNheOkDrHlz9i3P2IQOOpRjLbNvykS
ym3aIzfvr+gZvTE/m00h70tCvNVDQ9fSf8wD/qucS8JVnp7jvJR4xeLEihDKIe5A
JdCNYg5Rd2diMh78MOAxwRynVODBEoy3U7/I9+Mge1RN6J7dM2FH/STZGOqNMGAD
u76sFpBDzn/6DP24q7Ee8J7fTeHXbodvMt/pwAh7nzB053Rtg9gX9cv1Hj48Otj0
bBt7/RXvWox3kH2o0vPE8W6sWUvHyxgBVmGMXskuLOXiGPv0cwWTVcdBdq490O0a
rVbBau7yYD2XX9IlEwpGcEX/dXisUtFBBgAJ5Vz/TZuGQvVPB+sWWHI10n9bFHP/
yHsg98V8/vtqIuS97wjV/IUOKLog5UxTgDVd3YcwAzzEG1N1Yye+ueyHDyfqLO40
h4qgT13gTig+RwIC3otZ/E+VqymhEb9zmqBT9DsmbgvJPNfQH2kfmD2btAv9FFDU
0N6W+MmDz+LJ5/KDx94SI3Fc+RIGIWOvHFkYUw8iRjeY05rvGMX2J8tnCVLB9inD
5rdiCDNDEXxJvV19pAdBwyngCzKTxU3vu6QiqRVqEkegKHKrBT7wrCcKgc+wK0PY
LBwXX/IeNp57G/jOTA+1TiVuBe/4sjJTaGB+0x7it2Unn0COToLBE5Xw1CV/w6dN
9Y3ilQMTY9Xh8GsX/FEfz1iff7Av2c9czJTGpksfSFWrnQNzQP3BpZtEYJghmfbX
n8pLgo/nGuYLEZkD0q7AuVMvHHsHm/g66c5yn1TJ6AoTTwp6TdlTaOJoZm5l6+q8
HTLIEQS0FnAyuRbYHOrDhrft2CLdYkcxlekbtOQqUmJf5VN8QMb06sqa7H6aZgbo
lXze3khuiEitjap6W7HSYYK9TpVERyxo5P+0XQNEYyC8TfVkAizSUsgSJwDNww7d
VWSL6SuOxpXQ4XqZfSs8ZUuw5LwWvjrzw+3P+AS8HOdl2Y98HbgutIIP0f7i0WKT
rPTRHxGbPPpeeCF2JdcPDm963Tz7P5oWywYqqLQs+TgZUYe4LFn5OEXAPDFgNJnj
2xr5TSFzjg7t3ZCk9sHcMt3GAtqqQPt7RAZ8iwEkxi5/vOzcJNn64DvDPEUPSWt5
AdCv6hOyN3h7PV80CS8orytQkSukHlSfFkja6emgALYKVTnvQlXQEhtjbdqbC5mU
6hFnS54DF1+t+/km5AKp97zq/1aWSNj8QlMhnjTIrb++VjkfTeulkdTiR/+0k3Kz
FseUH0hTzlks04NhmENrUUqVWarolVdUf1XzWk33LJHC2DIk/lVMGfo7+1P3P26E
9W7hPTBK05x9gqCPnRKmVt7y8C/na/uovQK4Kk7Xhu2B7d+/Nw/8hjV2O4D5hFa4
Y3POyC7V8/XpJoiDNQzJi29cE4uoFk3CkV5mf0dxOMI1dQgENK+1V4Irsv1qi1qA
qtk7KETi2CYf1xvVGQ4CeW4MvDIIlxrfXTDwe3wYkoST4Z4OxKEMu8FFAwIt7VQ+
96319JXCP9eTtkUiDghxdfrUw63XrQQyiJPEt0tau5KSmk4DB4q4JYYDwCQmoBd5
OnY23jmjWnW6S/J8Rn+lxuT4MZ0xUWjDl1IJtXXTyxr35w2HoeWfYeHJqOjZS344
zrh7lIOd6rYymn/fFbhHLSqCeGX7Y6d2YtkalTVCkaL9GvHdnKdGD+4neR5ambTq
hic58WhE0T6bI/ZIPB8uEeLT8WTeT+7PxeGbmSAHlUEIZGVkeSvWlJ1AliXAeEJc
5hRa7I2GAnz6iGSVdSOIyRXvEEZP43/mZMGke8NjwEUy0awFTKPng+oYBBL/GTzX
KhmsQHoS3vfh1IZH/bo/bLSfWpF39Gru7RyZfgy+xGtZ7zktglpb/xVbWOSfrs+G
uMGbp5K5mbjhVBwwE9x93KLyL/5s5EIyyiORVWeVGGFvtCflHA4vQDFKSPWcF4/l
AjrK3MivMBIHbz61nzhMOBxXPbCPOCtq13Q8BJi8UVUpijeLBT4miKuqrVF/W7Kz
jU/ykTYG0SvctFhek6ZzP+HtKDF1Qbc9e3MpguUzDsELHW55j1XISf7ZUjGJUE1t
UAXnE04MaedcuMNcT7cFCr3mrYe97f3rzhUHanynSPWgP4IaEDH2Xqhu5Dlsq4fE
TGQWiXHwrbQ4b87b15+lAV6K6LnYst0Gg+uYaMFAkS1UUwjVxn1FmH8frQ8yEBvN
h4Z3Tev4y9nbNrQzf2P+EdwsZ9x2Ttael5quwh7jPDlkGYJOZuXHCtowzK+pGTRs
+99h3jWvE0uPE5iwuBM/RWdUzx8iWi506d8sYJUGvI/SkRg8UfPtcU3o/IwdBE7U
alk0MMvmwAzm//jnX/kpW7UCVj/5Un7BAY3Ett6Ex6wr9XdAl+vikGRSEmyDlzwv
Pw/uAzkdXBkfEAODOyOopiSpmWmVwOi3+1mXHsEvnDV+lYxwIGZeAte9xXfu3d8p
qaJSHsacCAyO7PtBZ2KISzJYPQYzXb2AJhsMDt4UmZgQEzWvsrcnd9CbRu4dVhIs
cQyBbdR8/RT3wu4fc9K/y1NBYAjwlHSjC63T6VSqKX2dJOJ9HNSMmU5GTosNGlUr
36OQIxuL5mKuELZg1wphxO9jV/I6l+7IiN+jkhkjBCunL6Oa2RqiWUc0mBxWM4hX
E69NIf/a1iJLl7AV+NvWYOt4fI/L/Y3VeC+z2SzzvUelm2ojgxel9WLToWt2vkwJ
N7ZIXV37SVOsevrROoGa5ixBJovuwXvosGbsc1eXdth6EPwzIsER8Cs/nZPGHVai
q0n/6poWvPr1ZsAQQGOhVmb6OGDuZnu+TKldSg6bxIt8fuXd+JtNg49e1bBP6/23
2fLjytWqst4359xai116PwaPfbTUuWiX/IaQXC/169edX0TtRU62+q/b3PnGaER4
0QS1Gg8AavGu2tg6bly0hVFTMEyrUGrj6KA1SmPkxRCC4ZYRYZ8lyAxzV909tVHh
VR5vXU5pWcJgaow9TlCNhKKJXS5rMcpK5JOAU1EAzb0BZ9dDZ1P1cBstPf+SH6qh
gIPXOJcM1FeRzgF/Z5UaRyFR01iI+yH+IsaoBiU7FCs9YmwDo1lKRLjNh1KDLgcc
R/+97EiJXxzXSA6SQtn5psHkKliPIgJzWiajYentvFJTe0L03HHetSkF6Es5p7Xy
ZrzP9uEmzRMcksqWnyC6GJGa5u2cpe/AXVg535qVe2Ra8tbotANPXGr3Sga3nsW1
va5RWDVGbH5y2jzpxGX6FXwvSBwWHPzTNJKajKqLTmzyKByNHt+7oBAlSgtDhWUv
eYEuh+es4uKYtGdWswa+63EpqyCuKJV0zckF6t+s9MhNOFMGB7M39fWO/wfPcTR4
U3Mbo+fp2kfX5lndfb9X8qAFXwQZDySYJo5Z858eveQzg2ypYsKnTcPE9SPnlNAR
tjk1YuN2xUkiUymI7pd0t2VK1Bhy5Ad9fL4vCkZuopIHnfZXtdUrNtIed3OMmBwN
M3qMyLdE0wQ71JMqPb4RIzID2QVm8T8ban7dmMx5wd80HXQO5fCGtytoN3XReJ4P
IRHyPT4uiDl0vbqK14KMk1c4LGTLMwd7sN5DD7yGLtkhGP4ZhkwSncEtwaXGV0rr
kSZdKobwoXaTpmsbEvfjefRASeG0Q3zvlOWNh/jzTy1ZsrG6/WXLEdppEY0JUi2A
Nrqj23CLdZwKP02dVexERcwm0mnydBYjxea25kYmWSNgDOL1Xz75hXfBdu3JbxrP
LTYHRBGXeAhxVLsr4Rs+rf6Lqb+icYZ+c4D/D3ab2wwC8eWBGobPkUGqJwUGhAdG
tg21DWpkICOX6jQd+rJi2HzLgHcuxPD3s7xQDsrr3oZe9mjFx/1oU1U7aJ4ZkRAW
7AyhodcAeU/I6SaJ8J+z4tA8d+d45AcSex+OyYe9Wgotakn8TvIVOqpPyHW2Skr7
UOLw9xZeL7wmo67t9wIB+/Xfwz30PdGJa3G4zbAJmG8gf4QGExt2+wV+Sph15D1k
oLZYfp//laU7cefWTpC5od9LZ6/7IjnO4Q6KcPUGx72bYDXuOdxO2YufdoXxaamD
YmCuR9Cmf+oYRHtgZc86ev14jr0k0uVpJw40MLUpzkbT2qtD9IDtlhAzK8NF16Z5
Em4Hs0DJ9nusY5GO3AQv8dqOx7X2TJwmMQxl0G74jWQdmNrB76R9AUo4iIwVVyZm
EXhf8F1fjICEYrORtxJcjjfKNxVMB6FPdEkp/Jk+lOWZBDBp9nh+3sBoSE3QV6Mt
+YeAi8283I2L6Oh7zzx3OzVbqYXnyje1kOa/HTJp54KDjNdYi2kzdZnreHupxddq
8l0IH/VJIBUEf3KEPGrNHAbm90BW1NnhA/Qw5r0YZ2qODDNWc1Zwq+d6FpYmUve9
cNuLSN1HqLKTDqcNPGd5OLyWA4P5jk5jh93SoQfOSxqVy6OOdpiA4JIY6DwlJpRf
wvwXs5hpZuAQ30Nn7pbPFXhGnPj/0E3OI5UgYcchXvp0tJVDFhqxsf0pOnB84YkI
p7LRtfu2/1c0w34Zi7HajFhkSVBbwde7jd5PDxCH7vJWtYNvCJyVrzhdeiI1haAv
tIVBYxffKwqKXeaxXY9s01xBrd1uqn952J8/Ke5PBk91snsvkEPFdbQUdz1p4L2o
zX66iSFDudpZNbOZX48nLH0nj+d43O9DYZ90x8SPkfHQFIr1joNiYGj6tUmbc9fx
RkgFZUeWuu+FBKOouBuTHzrRvmy3/71+Ocn84NAHG3v5Gm3HVM88MH9uDcjjCdE2
FUJY1EWk94y+/DCjAO6pEstpuUMvQ02TdBlOSAa05Z4MX/FhxOD4HmCNzytmT0UP
tHqIK2JhWKoHg7hLd3ThE8IDQV02Wnu0DTItjI5t0tyFML3c2V/aw/QGlh2QzlxS
QD4meeSo1qykGHouLREUVDVjC4708KatCnRuv7k7R1Hc9sMTpS0AxuRy13NkMB34
JO1IZy5CPF/UYoQQR2x7krcARSmVsx/fu4t6WeU2yPQSfzbTTz7U0PtMdbcMhy0j
9+Y6x7stkOBWHu7fclZcdCZlY+645shp4BF6YsWaW+sGebn03FdKZ5QRb/6BX3go
lM8HbJUwO/jJnDvSl48FIxQHHX1PIeQGac8mwFnRAnnsos8Q1tUvBRYE2Vub/lrC
tLZEFX5uSCjlPHVF79n8YxugbZeffg5YgAYx8IkIeLYcWkfhHDD4azzpalJAuqU8
jgRppib6HWwXpc/UBQCwAtJkoMVMNizEPDBgLvn85y6BHRadr6PCqUA8kc5NrGcO
oewOS/lnRGKlsA/b2ghamWjXtTSFx7mHSXqTY5eabht2LJ3vsROB9HV1wpTz+fRB
mQkVVSFNzorSWnGfGluCop3rkc7I+TVsNwTm3mmczgIzdytJRjh4qpoAlY3Bga42
G/5qXwe4AuFtFXVCe6uqTGWlbqX9iS8klmY4v3x8RMj/NYEIQu2nh9wlrDQb7PJ3
SS1VXq/luKr+FF8P7Q5m+m07ZIaCL8Sw0o1Ic21s/SPk0JHyIJh79PWA5DnrNPCK
YtAjIheWo5I2oN4wkLpPmimeeMQ/LHWmTupAiqAf82UYY/eFr9nJiHH3J7PKcBDw
MVop/tVOu3wW947oDj0g+M3neoXDBtL40zqOkYjw7+xELvFcy45ApdTH3JOKgqTK
tCAx6wZp5JEiCPuTdANGCH2siBhzC+e95Cg7Ht9dhFGvDp1OJ+EwdmqUt8UOShRV
HaARdttXHFgoQlqenQHJdDMdUJMCvGCVYV0KoYvH0ETqtavXx68/ejefB9ISDalV
J3N1JKfKA+CWOUdAvvWNoNyJboNyLLfcTnqBPeU8pH/BfsfxGg2HECyvg+lzVinb
d1bOZDa2GbVZd5YayLIw9Or4vCFyXpWfup7rX+6ChuiH06dadWNJA13bw7i46SzR
kQkWdTC9lqqTzfaAoFqiF1abtofinkCzLTbG/Ku9pnMAPy6FFiHSGgulrHX1alb1
ToMzCwbx8MborICZuctZlfFWMmu8J/Gm2GZ5Kx1F+8Bm0UMROXSqWyifYoVpTrrZ
2J8Mp1JikHSinp6Kq1LcWEmE2Fg161TqI9wzlu+D1mkTjWl1HmxAvZuI5PlWV5N3
3zMSlqEMNeIj0B6ILc0Iy7fkvXFH4CGtcyofYfLuYZzeQ3h+TerCSgT/1q5befFd
hXrvKkO1rl7xIOHhghIjbnHIsynPi5Wg3SBZqu9fUNCTkNBZM6uN/cBs20KOULiS
mebIZgd3iJBxPlE+A8AqFfZOlMJW8DT3dKlxolsT8OuEsk7eJt2NbfDkK1pVaagW
mcDrHFTsF7cqB5dQEp3OYjNJZ3fDHKhCLe9UG05Ch9Jpy9KIWijhicIURcPfgxgu
DJh58HoiKv/RHDJvo+gfQHx+sAWZFvhUPcLApFfPc3vmRqIXeKOyozD9lMybbRT3
NQr4K+03p3ycVnFih8ajAK4y734ihM3M6uNpjOUOKHqTLxQO9hGdg6BjUqkY8LRz
hE8GQwv6+qlPfQqYrtGrxYIsV8p2a42Azgtbp5mhjWIMUvjsP6XOcPfcRD7TKDaV
vWFRNygi8rx6wWtSjcZp3Lu2zdlCctZHarFSvOIV+lxSPOoH07ex75nKR8//JpXh
t2pCO+lWnb7luX1Sya8zBgZwgHCVFHORHxFt/AG2TTEIS1KlPcpqS14w+KuH7xXO
fkwuvazHc/Cb0ARerQw8dmxgrVl3KrEOTLqYPeWfbWg+P//YiEHi19G7RSYkrnDx
6GSLoKMwqgqoTSLsxVQi33PZ5SMVFOS4JEU/SZ8VRX96V2Agr78M1b+Giukp6V9J
y2cvKqCuK+0zApcAUVM5l89quUcT2KcCY7x/kXnnANQwweON+O8Qm5QKnhZ/UbBk
mjMAKv80OxWOVFlFlA005yhhy1VkK1de0ktwEnULYhiTofFJdhb5tqFTO8fUkLJA
4yfyhhMOz998L+wNIYdfByvQbAdo1qiIB1nXl0v+vAAtBfsl6tMMCa3qiMfeZoyO
gRqzSJ3H136LBzwgXZJuDbNcTX3E0Yw4oKFZBu9PE6PX9fS+pupGxNyS7cWlRiaO
oNuHqjx2x446j9u5ZJdmw8JGN48kwb/BGX3c1sW9PInXFlPWG+v3tBAG1oANfJex
3PfSb8591RFo37i944fJGUXYEtI4teD/88luJZDmBwSNfyMhmh1xaHf71iToWFzf
CWsUA3LmZFCSnaHtArT0Gzp28oRw59d81FGG24goNowYKoxVvpMFVmMbHlEWP+eG
O9k5xG+PUQJwlZNlLOOVAsmFKdo5Cn1Zk/b1XuumklI1nEMDwM49Fl9dPFySn+bw
nyfSn14yAAM0LzJgVm6rZrvmrJeLF8gueRSmpn/zB9z/TAZv1/KmPe6SjNSniBcf
X1w4LKhj/tlZxqgV5Zo6eWkbMq0KfGlgxmhlNshdMR4yWFYqtTQKWDtiyFxzXqoX
K+LAefsE3zQNXvzx7fYXinvaDk8fPu2NmzqokS3FVLg6EvT22wdoI9gHaXvSrQSH
nAUfWKcmUTCHXoCgXSAltJd63AgY8KEEuX4nuUo49jn8ZNL6QAK0GwKrZCJe0cg5
87U6A2/UwK9VaFUVISxOlsgRuZ5/ldPHk54xz4B+evG5e8lw9h0y85XcGlfxPBpG
IDkEQ5n2WL46I6uTzPuhCaKvM6x784pMYCrtYbvH9Ep73QGyIm5bhuMDxuiTa30T
nzhse2ONS1AvAVMpVUo5/x5NuxH2MyXVzv0yUkvUyWNsQvgBkL9J4lcHHyURdqvy
Ct0zi7DPpFSOb47Fj2vhyW9uEqJWBpYgqWjj00AGPmqakbS9+BnOF72aO+fV3dHm
SatvIeHysjCkpb/mFTat1Jwx7hV2N0cxInbLU/p6kN6/jA5QtP6D4OHMaGxfM6je
45aWne07ksCBR4yNWjreM6VLVdPvfqTy6vYzLiRISD3v7F/kh4VGedvRzawFPtyp
u6g9ivE3d6Olh9e4Fi7XTMfUAH51Pz4pTJr93QrQo0FQE1QiH5kSPQDFrK01Styu
sTw+fN0/BL87E7UG7s1jna9IcTcqIvULr9zEubZsJYzU6mKeG59Tz04wTdu+E8pz
aeGTAfTbmaBfWoWZmGDdSi/hZeKy4TB2sJBwVc0fgITjmK2U/YiwtZAotWqzB0T3
8JEGIT0vZ9Dx0gScAyaPdPalAOu2cyQrrrbbFB3tK0Uqr80rFfturRXccVL2+DTf
2z2rXr4ACy24PAInmgsrH2AfxlFaliHwLEfchohI1Mgk14vpgAxFdbOlKmlYRguM
ms50Rd24e+AQJ5+s+O+zCAleJV+ut7bsAfC9M/kEXeRTbeNN+Q4VnVGeNZt5D6EC
NG4E9VrNvyd94Gpopj8/GEGCWfl2419oQ5qztb2uUlR7t1zuxB9sSxKF5j9zKUA5
3ZFfkkKMeEP52hgPYflsNqMtR/GUle5h9R/PrMI9zLMI9OHPkezQa0fJo0k4XAXY
8+I4qP3d8KTKgrx6Gh6EWXk/MSgmIShH0o92BDIAJu8TH07lfCzhh9f89IHR91sD
CHVcxXQjFd6sqXU8XxCv76gkhPOwp/Fo+1pVPLQz5i98d7GPQLGui8J+0Xo/taRE
1aXmDy5VcvNT3VQLvR8cngGU5ZGUwnLga/K1oiz8kKb7kcn6D/HiggHwrqvFvlXU
96IvU48ysTNygmuCJk+SSNca0wJoxPxq3uZ14SCJknL9jhbxdPyj292XjfnOO9Z0
m0nar4xkDPaO2LhCiyQ/g0+Xwh4CsPkLUTp8TZbopLYlCuMzcPUwMQndRCj36ef1
D2/qxrU9yudiRUHx44B29j7McDOO7u+3bwr75aRcmXo/hnQ27KS97oGywpqa0hiA
bI5t0W0laDZAk68k8X5pQ2VYzK1Gd7zGX4kqHQYVVPteRxQptrGfUuCGVUYiM7hd
JdH5tdGGEMxc49J/+D1h1ONZZ6iKskDWx7qcTWGyUDsTQy/d2hbmgKfwMzpSFojv
N/YKLtEbwY+kNSiOFVkeF5XmaaCysm5AxbHqDtsdHzKFArU4Zb4N3VBdErdcV0bT
LAg8WyW6VEyI79OuJq9BcQr/PNyjceDvF5kBWLdoWf4TQ3Sexiez4uT8OMDBig0h
y5VhiBhZO8/gJiBck9puaQ5wfk2E5E+BGy36hX0Uzk/KXbksCWbUb37qoIpfr5/O
YYlXicOjRTbk/AKlJBu/Z3qqWFNXmSynK8R/ErLfM9Au5sBWgyfxijAbo49XNg5P
IVnOTIyafu6AaucRKe0QPd5C+tR2/WelJF0aiKNV5unipHCI0+L5CsDLe+jgM7op
8Z80xpIug7TKhy4xBcd+W9iSwjgYEycRVJtPLjzArIbzDJ3nPea84CCRgUL0EAlK
C3UwvN6+kiPuPXKD1N4+O7tqnGVIVS98n3oz849a8NcJ+QU2uwR8rct3ldUz/mBP
WRCEQF04e5onMwboYJZATR13EAc8J14uXDQmLkH+8/Xb+Mx4c9kme3+NA2T49P8M
VPiMeNLTkKsn0jipU3zyi7sONDtfDKCbsYicQ0OGfXn8Lm1LRiWX4SuC7rwjQw7P
ssKHKMvjTEI/rTK5+sj83LgHJp82IhyRlDp9AG74d8jZ2TAnHIqr6PDILRK2rVv/
7MqKLOWAUbIunWUigsBsEKJGFXwVKVlcEGm6Y5S0EQlo8Soz51Jl2jqYZ+Ow+7xt
3y/VDXAOPNkImFrceOQIErUUDipEUbHv6a9EkiuJFqNoyYncX4zrSn+3f8z+LWKO
wcf007mUSILOeMHOcgE8GUjuRmlfvng83Bs9SMdVCJCA6wVSi+IFZxaKWi9PX1uH
0xi2Pr3len0giRTMiiTalgqbAQaSTilK6qK8B3LJWzezeDFu/b960we1e+Zg2Lrg
Q7q2fY9qHFYzMcb6p5J0ciW11ubxlod22HeqWg+R+f5oFweLiaNEYopHn0Ghdnbv
UkpfEiPNmeXLb+XvjpEVvZfifIS2lnBkgz5e5HoDTdxdRWjTKySuk1rYhrcyRWb3
ld9vGwUwwQmTv+bsJ3gE670/rNqEE4bE/yx98yKSbnhCOHjAILBbiq0198jE3pzY
gD7RFG8jGfeyUAqYoZjKEdDWJTOmPvYHjH89tPREnDNLNhYetJsIOnjdKJ0hAY+n
+stEEoHs64Jsmn5vt5XE9oV94ZhenoUmS3KDHa+/dvz8X4NIfPfmb5be8uKLZ54R
JThHCfxSe8P21D0pl3IhoSsxj3Aa+PEQuHmCw+JFeSaBO5/0pLVvEOt7u11vWgTI
11lMqHnVrDwMqdZiPzY4qMe+PoQ5ZhhfcD9EfC5XLa2UE7vQX5iKcRjS7zwStghw
//QZOoWHdRYwZdB2uvf0w4cJH6R2UAN0S1QvTJ4z/8jeJWMfFPte/0CXhRhrfgrX
7YvZJlAyqLEseOyAireEbWN1iszYlxHXMXXc4ltTZSQvd8xbQoKkaR2JwN9VV56O
XmZ36gfs9xju0bcSaJCQjWQ6rTvYSx86qzr41jK+9uQLPHzstT57brNjLJjbOxk5
WtZ2qeJ+28H1fPAE3uxUaR0R/BVAhMbphK+Oo2bbAoT/nxTJ70mPdu91nVlkX0T6
Mm1lOjlCg49tkJq3uQav/l4Wdm0nrm3dykz1veDiXzRZeq9I0Tiu1qb0VnCJ2Hsy
STntoU1APUT+b6PBK6hsIjQ1QiBAgQVA6QZUCnoZ81n7Q47TDetsmRn+IWEESA5/
bp3unpzqT84kDJRP/xXT8M+5mjBsXV0d2O2Bz61pCNiBOIpiPB8M6WL/kcF6B3XE
wkuaeR55lVwxtAcDwIA7FlKFhoZlw059o0GjSjXlBxsYTIrncNMMfQXiupyAhzEa
S09GZQI8tWu6RDP7MrVFuD2ZP3f/jPhLXv4AHO4TTLjOH5gyosiBGga1YwlIn4Lp
LNgig5DVL80mmf/kzCX1OPvr88XMMLvswCrjO/KKcO0RiKvnX0J8rWDu05dSrIER
B7Y52+45xi+yPKm007e/fV23e4qcLWusL3wnQcwbM9hW+ZT/gh+9Jh+8CPjsPiod
stMDGYXYwpiKAFHKlTEOV7tQkkZ2UWzSm6C8/gXELEygyxDyJDzP5+yUm3iiPL0W
pm2z4doZ+MIBU0pPZiqM2QckzUU1hT8TiOzFtDMPJwZfqV7Bi9wuoTan5dAN+0m8
gR4ZZTYOLqH3/4m5uq4yecgl4/jkjiwse5d+nW/HPJgtIj9DuiBZr3A1/hpJEiSe
EORaGDmJG1Xprrt9lmO9HA+tleNEmyohl8FRhBEqY3oRE97yJJ2LgkXz4ggFtiNT
2lBU53ktNAew4bR8pL+120YPz+AhOph/6WtmaFUwxBStsH1iuyBVVyNfoF90QDqF
h3sbV8e+auaL1tm3dZ/Lnvgnrd1TRG4EAnLsGfgWrO0TqNt0HvDiDUYsICB3xZXs
5aze4ZKAL8taEkHNjII6epumcf4+Gv/S0yAk/syJlunGGRL4tZyxAWpYWjFouoRU
HyeMbw4tm2Mb/q6Py62rGyYNETYKyf+gXCQyBzyWCg5xFUVdyfyAfWUD1kXDGVt4
Jvf4Mhsn+yNh4URnkMtjyLF+JbFn3qg4qnPPXmDUlbj1O4fK1DWL+uIWoC2zfRd8
ccZYEFjCe20Da/4yHg/YdZhIXWgUdHb5vgAXEtOY4H57zj73NJcppV2ICVxJls5O
EZre82/JHdvPRE6J3aaIfrO8eyfmcGeDLWYd8ymo/z8zMYCjBK3tlENQ2jlcoRfo
vUfN7oXY/rzOg+uQDjUrCtWEfQ6Hbo+zeeiNxTRZUOJ8YB5Fbta1Ri2oqgH1sTQa
TspJ02Hcm+ozl3h9S3Bo7+HHUw+Vi01/Ja4WIoo7p/v3eW+N7fTermm40jIcaU2u
ZK7GoAko38PDki40X3OvxmtLjg+ck0czvR9gvt9T2Sp9+kyFw56rPIWeGZt0dMjP
cLLJ/v81totIHCA3mBKo4QLFCrrSMBCxjosFDUgmvSkpc8fO5mMnhXrcJtOQ9pGs
xQ6FUs02kwspzYE/N0mnkHjn9Xgdy92QJnzymBRiKYeUiMsel7abqQuyRsPNlX6Q
iNiA05m3NgPORVjsx5P/UCrq6tqB2KvdjxpL2TO1sBU5cBEVkbHkWBpJnOn/i0AZ
ByhSoi1KzdJ1k475NxX/ufo2KqPcqUk6UzA3ZnZqWf0kryESGJtbsGwitL8YFR5G
hWPfPdsiTG5isQgZfX8rvktpvooG1ayEnn0u2tRhydaH/H4jLs00w6QHce8Cxnql
P0C/4QS9RVDm2mYmONF9+66PjFe+LX71F3pq+E8OBsDjpQa1lwylT9FQcwKwT1ll
lcWd8cPimP8063gamaatJP/vckTLRBJOSV/3ZGYlPDO/3cMUe/S8G6PYuhuBOvbD
SIgxqJ2UqqNu12M1wIDf2mqdOj/2M8HOw1kNNz2lHM2zLACkTGCMqdDzD77tzz8D
4lMZmS2vAWqIKHuSvjAegzpOuw+8NyIB21FB+zYAT+m7kuJWiH5sCwqWySA3Lfy6
Q4YalcIpqxIMrRlZZCLN5sg4xkllIlWuXkiua4CtObFARzbNxCnHXxn5EzxtsSkp
ovHuSddl7WO1ZwN02EzjSP+e7qiAKVqbkAvKft+YFViEFYkqnmzw8SwUQN+CCP+J
uYr/GCXsAIDLDrct6bHBqKNoCN+0PI3K9gWFNJE4b/McScWrIBJlIBxG3NfoKztr
zBGDH4S1YRTGUYnWd+I4c9g5sSiU0eI5ZcjMLC6kL+vX70m6vBh3v5B8lG2TWPhF
aai/iGiqF9z63aQAm8BYlOZmI/nAgM/6Yeu0BqM9GgSTK2MwtZxf2FNmokrUa9Im
h4TMg+WMU/R4S4xokm2kmIIinphUK/RGe1pYXtHltb4UjCm7JRHdUXscy+mVl/FG
NPP2nb9sU5qkxPYRvBAd53z8YEK20WQnVqH6TX6LJ/uGZiUpf+PCTdutlmLMDEil
Mpz6/iIKBFR60kGF2kDcKQstMWsXVrfIsV4SXVaoNwZ+huQf2jpqnbFcOOvrVNsC
WOnHxcPFG2c69kXgw8vcReRUcDr0CdJx6NQgouaBI5/knZrpYHJnhR4meiaQ8amo
3AjmCDl41xQsRsO/SyN2pGmZvL1dpuY/B2Th5b2lFrQ+DXiU21/JUjltQmpDOVk4
1ImnnnXt5yc/7IodOLaJKAECKlRU+hGdRLc7lN+M70o0kXDd1qGa2UmYtUGNeVj4
LZfTK3SLDj2r2fz+U2h2k0G+zkqs6/BjUY7wT5kQetp7ctKaDxUdYc3qPOCgWakA
9WBJI1nZBJIxuQX2Bkj3jsuQJHFsGv9vDLGhJishd8I3KEKNk/UA1MNjq+NI6tsj
1m6qOdfQb5aECMHBQaDoP6KA6J9DfS0cRyu9stgl2X0v85Ipcc3RBE+q2Av1gFS+
8DTq67AIU3JAznzvmWFVwv9IaaMACHdwEkQrLufEAOZbKo37v6JhTut4wc//xRwU
m/vK0iIpvI32LJnI9a0fZsC1p/lK7bPeHdcQhlZGoLn6d87QWSTgvW4kgTlR950B
+Ie/l6LlPMmDF7osgYRIVoaQ11e+NVI36S9drsQsjtVjs7hy8qN2X+KEivW6Uzks
F39iYxaXyfPgoWk8Uk04fJ9vmENoR/xhRyzVKbHsCBWhBxUHLP5ttnrHz5AnIkSi
MXyvNU0wB9fOzIVLNTTa8F4VttvqX3WBdHTm97qkqOcRcFFq9v+86rJtB84DQMM3
7RgLDH5x4E8dMULjBRGx2rla4cBsk80oSrnJM45PpR01prpybyqzzpL9aId7eocD
V4QlhCDEqAD2p6hNMkFnjylfE+TOw7YRvdo8gdnCHhOvoc0fHglxUdsws9cPzKlf
/m6KEH4Yn3Rzq9QALaAzmLkXTAlRuZw8/SIZ1epyhC9ol5LB8qTCKHAluspMyp6C
RADOywpxjJD10+Sncry8Jn7vIE531JxOZSM2hZ4A6kNLpJ/q6oMsby3VFTfiX6Dl
FznI6Cxm4NwasvLHMsAFuK4yxbXfbT3Ux5mn4dkxvelHcqE91+nV/HyFqeT2/Jip
eHaGXnkM/Y/EQBqka2QvUw5H06rJAP9DxLeKlnsL5uNJXFk6yGX1KyZ1P61nrbFT
x0zsZDKHa2iychZ+C7K2D7SjYR07JMes1bBtfLyRFJL+RDguYxdLzqQV+p7lHbWM
ujkrLvwnkJA/ZCnw0dMjP1HG6R0S6VMZo5CB3mMXuyi2G07vW31DeBlEa8sLzSjB
0+daH8C24QnKLKMCoGnDDBgesgcsLO/zyEv32ORH4ShPXf5WyiRil0ft2X0r86tN
Ez9rSp9wSRH48iFYa1Fq3GN++NzJwV1//9qs/5BRlWIkY/fwaMSfQoOEd4SvZExq
PD6HnpW3ZB8l7bkohTT6T+uyDigx/Fb3/vqyn5IPqyTN0FIA/SzxHtAy871Nbsna
ACNSc+9bbaKtuRYufWhoDXu1PJ4xifv6cH7Vwik7Wn5zThFw/iOkaOk9FpM/nARp
2p3ThL6yDFmNo0SpvSDbupG3vm0Xsk6qumqCsnIuOywBtLyABTxzKh4abyWLzDnL
uY31wqyeNgksZ7PoZIWDr0MU/HLSFpDwxFzafP6Ia8dLkpg2+uxSYARCzo0hbCIV
JstiE2HDgoZVtg3iUndm6XyP0zNq6Aea71W2J0vgocfbBmXAf5yX/NoY6q7cgIJZ
ytnVJMsvdlQH45F/+wbJZzGOaYL9eJzqY1G2MLpR8wLgskZPHpDOBh6fIVQbixGu
ybUVJU7gHvvAGfiff67mPkMgRTV+pT4yv5v60OeHnmAnrPRpu5X6KjgMjSaSETnx
9sQqT6u1Uom0HOY6TvQW1MLXyer2v0YCX1tzOGaGba2o5C2cXI9bNbL30OZ/y1m5
Cv9Eba5Xc43ziQC5AR+8qbSKdQc/C7WX6nRI0YhM5mSKMP4jK/mKKs8OGT/tMSEO
ovooT+sQxfC/H+P9hNJ+JvcpYvPZ2+zQlsD0IaTtJdUfx0QVigiT/Ftw+qZSeUGv
DnM0jw5nnIlbFXYZjSlTrlvz/DxEEpXF+NMKr88QRmkTR4x/sFC2NO8PbOePZD8x
DZn+hdk+boqE/KFwEIHyBZXzgRLjcCwuae6X2ln7XpYfyWIc4XoaR5W1do2rkHYm
Ib982DmpBazzK/VVslQ9ZatJ26Xfir8YPp9BncGLKyMPVjLj4QD5u9uXU8pj3QI+
YYMmFJBrWIJ9jaYcvV/uaHF+xXWx+KLpZqjHCmtQdIlZHOoFntRN67lIQL8oo0Ef
Gp9GZzo5YNYSD78l7KBj4vnbCAVN5juns3of6KFCQ6kf12mQLSgGzIVX3eBBWKAJ
DD8Mc57SDplKA2Yhd05HHWcDscg38hcxOx9kyolOzjMZHzpISnpmhLa9Fahv+XEX
/B5MOORj70QkNfL0SZt3CqFd3qjG1mhvjulqgkQmdfN/M7Z/J/zxzji9gRpeKRsr
QNAigINfzfruE3Q4Wq/ljOFL/nAaP8MMI4NaCqfMVl1qHrDRwR7GrQNFaqdUqJuh
cAhPBzATaORgwi1714GZOK7Rs0OTs+bR7/CV8qWJghHNMw4x9cpEqK/8VwqIAw2V
lXECNyTpn4hxpQTOORTYbYzzhJytRI+pF5SPqBFP5ULNncAakjQ7r3WqxdzpG/Q3
ZHlSPt70egSIQsyGDFx+OYb2I//NtZWV5clEJkd/XmRcyMvzVpMpiHW780mVbQ9Q
uLzbpGZU5arW4mFCeRCFU3WpxVXpbLXVV73Jrarsc1Xwe2jPFFgRIOl76EqzZ4uU
lnBIzyqqz2zzu2MQeNkCf25OC1k3lBN7jTc2jVoPXEUR+dkZsXp773Kr0S7CkkLZ
bfWsTrK1DVQWJobqWthcWaxI0PUSWli5hj01S7HNeeWSWe/LM5XTjjUQE2mYYe6g
6CMJVhKrG/s1YRzPMldPTm7lyBDF2WXfGuMIjqCQeR0m7ZLu4kz0q97fSdxAHeFD
ACRy9+VtSfcPTVql/piv8S6IAUTc4uQkxm8TYcRzDGzQ78UAWy/D8GWiDrX1y/ap
IoVeemkHQFHq9ORhhh+4UoXdI0kirvKbofHcNK1OSrmlFa0/TKQr2OAOsxB2sfVM
WRI/YdYgyzN1KUrTM+emSUWvy8yYq9Pmea7Z82S4iXUP9q13DrQAYYl1EHS4bZ+q
7q9fHhjJbMaUB2j/W1NMPOsnIRuIJ980q26ZijGP/q7OaeNWKx0rkg7Ah9oqS3ey
I6/9Zia3jwc4s5/CdGghu3Kj0Ci6uuJcIcW32UTnZuZT4ykMZ+srJJWPmTcQRXvP
LgIa8YTmHzCKdyIFwe5MdNQFlAAVv3FVTdDOr98SA9oMg4UfQdOx0IfTExvVORV5
6lg7vCD8aGgf4Y4zsR+yMLpjiSyg+9xZTkQvh8olfNhBFF5f3TMgl8YXaNOi6Z5q
vavIo2UpWBpMX+gesPEIlXOlurar1xKGRr7Ieye6qF7uTbYc11ZdIE06VdH4vWDl
6swrfAAwjFOSlkKnKdARFqc4B//npiOkPNnT3468wCy3WkfGQfg8FHCr5LJbX+j9
Vg0n0CNrWLnVkPwUktCAhqOP7FaOz6wFnP9Aib3TRNLHH7xaZwKTEko3/mKQgdJ2
qb5NQjbdpXUkNHCPLmMP+FshNv+OpT6CS2mppQQq3c7N72Asa7hrr1/1rb1fcWQZ
Vvk9me6WiAfin9sBJ34Vn6vQ3Kua/KFc6GSt1bv6luHpYLCfCnHR5U5rHFUT3p42
l1EyeWtslEugVU2NCmW/OSqVNzmIF3ACfZF69U59sFy2KquAl7waFyMKTTYc4ADl
9AkOFR3RkXbaYG4BBYvwyslOMOPsK8bMbujzBC/T17Hn+asLmEIFFPNeGXatyukb
GziVh+Mjwm8ia6RZLLQqIh6vVcIzfysP1LUfHD7a3hotJHUgR4BKm+I+EV66IgXX
PBusM2axaw5B52OCCKiFuBYkbsXoSssc91JyptFeyvMrjYgYXEjc+spbTKJOTWs5
BnBbXa9X+zRDcRlYzRTXL2dHA8U/I1zP9lzw1oze/lMGTNl5AOc4Ad+rlxbstWm9
VQJncChEPA9+zylYRexQW4uo6+kid5uU63B0B+xwumml+ezXMcTMXj4nhWjJTr8O
WBV3PC/inmDzF1cIGc6omd48EgglltkG2hCTrlMvcbuo2kedtWG7DXiIMxv0udcP
q8X9byEVJjnEq96C4BZaBGDEojFr+gckSFA64lZzh9f2P6+6nmM7vC6z4BTBW330
L13tHz30+8lv7RmXfj+kUl8h1PR8fbImsfhXouxJNaKTka98IE+UD85BJYlf3s7K
nbL9UM0VpnqvQoZCkqxp59cjb43NVeB2qS2yySf+IlAH/ecpOq7wCWc2lX2fm2xX
RunhM7YpLHThw5mJwO0YP1vPfzn5yGL5xPuW0K7AR0GisUZMWIvFr+S0NomJAJr9
AgY6Sda8rjYXxq/n5GUB13QG3IwHA06yiG4AdMGpA0r3X0oWrQz7mFdV1D+yUI0h
bC4zDvoVahFBdnb96nx5lo675ATJuvs30uj0jqluP7bsF/2lKarMvWFGOMqneHNf
aPcZdnPETJYCfIJ61fQlplHrnNq4PQKc4fDsA7x9HDlUXrawbgDKbQqB/6wSZXxt
tpEgcTCjiAgk3oTYQ51A70kGPJU+sk4AHpK6uLO+xZkY3ZqEJh3F9EzB/0+2ZXTx
gao6Hp63SmCq9BTfvL1Dvn6r8lKSgTJie7FsmWP2SmD7rOtooE5CX3DFuw2WdWpr
8aSdd/3OHYhgLs7mH1Zdm1BhYIFNaW4mTGT/GvObusSkZmsC5NjOfWWHKY8g440p
fNn1ULU276f3BsOC4iSV3kEoOT++zRIK4YjLEM2ZRX0jqBxRITSov6Awr1Rtwgff
QgaymTEObVMHS9Y9Vgw97yXudv8EEsaGMHruNMUw8HyWXE2+fp/i0j/rzQZCJkNJ
7M8KhfSVqUN9Pj+SnC+o45/lksLCEntyggTQtYiaGzHUaSK4QcbDJ1Fzecqa9M6u
CMrmWHuSmh2KHWhncIWpqERLitjt3BOwm77xfDBF0EVQuqs0pqNuzXF4rKKlvlkL
Jpciz0CW1hw1Qx6lUJUEWVobyUVzY6MjamQ8qPGJ2UdiItdo+U9NRtCg7OACyVWc
mW06TWw4g4DfgwKNDkxtMy3/BV0UkC2WE1LCkcMo3tj/nVNzd4Nl8W9ba6tzEoSg
EpkQKIMid964itRU1XqtzlM86Tq6/OjFuf+bJMuzqRFfaYX1BDpL/IjRdjurfYPK
m3GlmOlu28KJ6qURLknvd0erXar18mDoR5X37oyI02/8G3p2teFH5b6mwfzr5eZv
495MgOMaftwxQB77KiEamZnf2NH2vd/dFEYmkBQCiDZa58XEvX5MfTTC187kVgUg
G8S3xoHAtg9axML5AlDi/EhvowQPHIwOsU3lgds6LoLxzRTFQwNETVhAZ9XxPP0X
h6BqJ9ty/FEr2GiuUVVlG/hoiVBHBCRl3ZVuU9UGWjbeErF7MpbxdMBIOM9VVxy8
6wHBvk0XMRG3Dgy1O7IkBn6PBuTwBtb1QUJWcLCmuQxdiMrYoMe7uK5IT2hOh3Cm
C3f+JrOLRlv5BamxnUmXrDg54i7ERD0AS8861tM20zjGWxi8hlpl7j6BJv+P186T
+q15Qtg4cAqVe88DvSyTuUuE/u4KYSu/KEX1KfvBcjMRofIhhna4lG0GWSqnQQ2n
NNezpxzrql5F/RV3QUhsLeVN1OwnSNy/G/6wmSGcVxKxvDv+2FS4fwYmcHQO671K
cwqaMCcGisIlkIZMb7BhcM/QobS/QdFortdKaXZPbomm+9Ouono0qM1JdWpqiznL
91bIGqCPEseM5/AwKOQIJILOf58mOqXB3aciAZCtiPVQszrNCFpvxCMvBGd38un+
bfvAZKD0uRHtG/Yg4mFEGSTfkeJ0jT8JxEvMXCjRhWGq5oz3vIDzIz8Pfc3KnhG2
uPfYhw0WVIrtUv1e07QJhmd4AnGze6AkSYVt6iDTFw15sJMdg8m38I6CWSl1auNO
oE331+CXacievE0lETKWP+6F6OayNz/FnHh5fUV9vPp/ufSkT67GaFOOxQtJa5Al
XOfZYOYsn0hgt0lNSFu+mXMdz4QVbH41PTTf4l4GUE6eKpxKupwudzD9npWNZhkY
Py0U+qmvUz7KSryFQSg6Cy+zeCP8qzl6GRnZ0kd6tqkvaJ/g/UPhttituCXUwDG9
sbsDJ0gIdwu2a5yk/VbMIVV6+B8wHoBt7c4ui9WJVoYotiC7reW37lANODNKbdF2
5kznHfCQhDHIVmKV0z8HWP8dDPCmB4OQF6pXGNpjy8YLTbRpuDD4YnIjsR8XMDAc
E0lkMSQpzS39DPjRZia+ozyEblu6H3HgXpJEgUmXhQDQ+vDe+2/eUIQsgA4MM//Y
CeYoVf2IE1sgAvu0b3AK/AO+EPlKUV1t1xVFbRHFiv3ma2i7ui6XcWQGmJjs+S58
8/I7spC7OoqriRZL3BkAUJNiyN55ojETfuymofWnlnDBXeCgx46QN4nQauWFAhoq
z30cSST571HeYfWwlXLvzFyo8vOvN3HlZEy/FNKXQ9T1CtTBj+j7F/jMoN4zqqVF
XIZueqNmmAjuQliF2raIGwJ/4b+w+bLy7ZluCkvWugNhAEUG8fOwT+MOUdlY7mu2
MoIYMJs40fizYlDgxQd3s/FFMJy3BKQya5VgsVeSg5IarnkPJ0dAb/dZnWPBkBLw
anUb5c3Jh/Vx7ypMvL/+pBviyGZxKoFd4ahzAsLVntrFd3Pw3Pzd6DoEmVfpJhAY
y1f0F1uHdloTcqmKlPgappoDMz9Ozw36NzUIc+mCZoxYdPqzl20uwuMd2sdje77g
cA85Uf9NstBxvJcRvB2//ObEunVNcRYVTNTRX3k6OgNbacU6j5yIcYuQc8ZRUdWe
tdONnJmGZ8wOR0JxyCgXC0sIEGTEgPmK+I2zXLbLoZFahngPeTewVOAVZ094pHBU
9WW6gIJW9I0H/0RbNwtZiPghBGtFRV9gmpFwZnr1D1TMu+YboLr2IND2EDnwp0sq
li1nPs3rkmc8LZvSqjpzZj3LzKuia2PiC3TMwyTdOr2TzeBngQB1IqKlKsVpvG2G
DAbWo0V55xAZM8HrqX7PIEPCBv6Y6G0fPMyOLKQZ/hwkH2muIvMz0nJrFe0gxOPY
Yq6vJbbuQ+MUQzjrWGkgc+6KDJA1PDddRJRuIUFr83J5n5akQcnVtBn9CkQlC0s2
m1Wegv2OEMHXl87HQobxT9KDgmgol7l7G2lsQIOqs/D2UerzrgRR416BxAONkMGn
JR/MT92jPJED20BA6V0CWUPBJQciHADI7NkG1hpM1kdC9a/wyYYwUKCH0h/VhxCd
94/kWH4348yrad7KmPit1E66eZudk7Oy+tmH54+1ifbspzaFuIxWuEOoFrT+3qaD
TtodyMN43fnAsRZ5BO4X/hAROvzr8hErL1Aan74VcOJUtlV0AihA1toFJbwhlSfA
p8G0+zUorQ6JPIb2QCduLTE+MeoUqKui7/auCkA+xdTRBkowQNm6762HIHvnPbSg
vYxg80xvQCV5AGCN6w3Ox12nlfgN3FOksEzdldJT03QXZ6wULsoMeRq+cLTV7kzc
BuqoBGy5oOzEBYgquCmASD2aOfhgpaVVxyr8UnFpj7rFD13rG7StBvo5JoRBhBv2
u2QMIPKysNSAMaMocasmfnmpsxo/RzJkjxLfnowzUsryRiOez9Xk0ZWXyReV6EJq
1a6P9QwKK3k31dQ5KusSudCDTSf28Mg3PkvD/DmaNma8C7j71lczywKo/tSU81I1
4skexRmR9L3eFTAcgXAVYHyKPh7ZogtKJhuTHJWF8CZYKFv/N3dSoNfSna1HWvKl
siFNoTjJtFBXKnMv7hH2lQ54WzmvvmQeT/l6cinLsa/pBNf1nZnf+89T/vDl0cYh
sF3WdRZZt7b36IU1Z/Yy4CORgvUuFRg5cGsQqIYVpHKEd0lK2LEzUjW9gnX7Y/Yi
M8e51DMHa6WFmfpTN8KWrQMJ1jn9iyab/YcV8hnJBMPvfkjmFok+WLM3P9Q/HCzm
bP70xFn34Xf0LWWsG38ElfplKyq0yplo8CJ/1NQOkpe2481gXiJ5jHK8Z9bSenXX
IOZfipMmbdSuC8YF/dIqrWyJnXBGdlcIVZmydF83je1Ks7lIOiJQu67tXZquZ0Oq
k3DlPrmQ4J+63E8lTFu4kOKeo9bpkHbmSSY9PE+LMLbtVnskEYGqXFKmdzscXUiS
nv0UQuyGAhWP3mFVskLwmvngZGGwweMMn7EybXxDUig5+2DRm9dCGhFBR2tkkgcK
OjLAafghCDRIHJciH7Gmmd/Ec4XpaT8pEJa9lGZKyDYW9NLNNXxss3FW6Y0gafOX
Q1X2oCZyD8gPsId+YoRuFjKy4Qj+qwzXiEaQRWbaUBPd2cft54+EB20wHuxz4FX2
DfBDMofKjexO7Cm3lTHgMJyLeX1xABcSetZ9kQu6THW0mvaOEzPaVx0sZwe31HEx
KO67LFh7YtfsgRbuo+qOaqfjWqWJ/k5Kpoi9Qya+8qfbzkLmN/Zw325WgMa2BYRv
DFZC+Zf+MUiQX39JG06ULi9zrr24icHA+diZj2oc/K2nUeZJsIZ8h+EXqJzlu/r3
TcwlSfG2iPHLoTtXf2/Li42acZEN4dFP5qOs4q0Mxl/nJjBdUHbHuwlPQec08XFF
0Ot95vCjJMcOOgqR77JTSzJYCTtd265U+jncQxSQRTKdroMP83n6WZ1NwlQcrYF4
JnYRSwJfDl0gsVnzADHQuYKeY2043Ed+mtjX5CoxghMY3ZZMt59i2CavUzj2/PhG
Kp7Ub4ec6F021G+Vtcm0FvJFV1V6j7wiZVSsan2CeVhER3y9ZcNFoncYHwYj+oMZ
O9UTnhu1R9u+8Q0TJHoTiLj2Rv3CT2Cg8iYPUWeWcoQncjHGY96M5yU4jCJq/lH6
n/kz8dz8dWQ7I7CDrH8SLlbt2gRmTCLWIagUkkT9TnRUVNwGCvNQdYlRDK8aLsVp
+4vVzni6bTI78J52jfy3u3C7+EuGekJWR0oXQnK7Pd/+IEYak+FptnLG2sh5OFF3
UFhZg85Plbthd/7Ad/iYlvGW7668wsjUezuukSEMt3RumYKUoI3gaH0yBtzEGRsw
3+jF7yqpxjnK5jAKgg7wzTx0AU47NRQ0QvIH+oHYiYmMOV3B5D+sNVEcoOriuVfl
nJPJOBFjb7elfui1mkCNEIP6CqUZIzGzGOPpGkS6iik2s1nQZBgzANJ/wnj48V/Z
3j5i4zqZU4cj9QIvQhWXB4bNysKY+BZUqcJGbiAMSit471WeESXQbnvWFo/u08rc
/sjvkp4vLxNkF/xgozoy2ZGFbllj7WvFdWQJTEFEFmP9Ke+KftSktVH0NdiyCUAw
FybKuBvcLuAevr0xVdCrH1aXsPl4NnyVT1HCS7K5M9dKXCP81/lpe+HhLocUUPDJ
Y0YAlfMCQsvK2zaegt3pQ8xkyYcgZQe7z5zL6hMjR/eMKVwm4Hxj3VUBhPFplWXp
VccVHKYmOdAYAKX56cIYRjGL1oqXlQv0JlCrkjQmS0rPfV41CZQ11CCWtm+kH8iV
73xmEmWGoPeLUkRdCqPlCXMOLMXRjQ21WFtZqAgC5hlgR9Su5rqU3brmmBjin/7E
xsAUtLtiNSRdnsXIxP7UFmcjr2KYhrx/rQiOdolrUxnvgLgdklpe7UZcpoqSaHdH
cmPLcXr394rUie+fmM2KV1sox2THthuSVDdufYQgfhAN3K0o2IfU7PtHGE5tbAnO
KMNiM0AnnUYLY+grvDpJWdASGUfKry/Itf3rD4KwBpXryadkrHRkR7NNdrU/mXPA
9KDsZVqdxqDvrWEpSn6oDp2U5eqyT8+K/dj6twLeFVbyK9YyIcJP94cvy+mNJ80q
sr4dpSMdhBzhumnnMe3ehVqCjfX6+YiGymJKq21P2Nz//+DZYa+7IPxJehmgKGqd
cgMiB06N/KooJfgYeuwHi4st7qEDlUHGRwAfGxZ6GDWLBMnmxeXZGy4Awb6Anqee
ULj32r+gcuzY0JYvaof5DxxA8xr6kzK3aiRE3FHsmnHArlCHcDBPSgA0V33PrurF
q85Ful8kV3cnevzH1x32Hq3QwZxvH7KuyHoLPz3PV/DsYdcrANwTYZ/s10iqOAyx
n2DWxRGtpn8lf29bAiF1rP+5Kzm9HhLUq+xIWvzgadQdJxz+KtwRY6qz7VryBw5y
vJiVdPaKFk7npwm9dTMabexJ5ltGhg2/fUG4dm2fw2UvNd2ZJCfOZn2LFUlCrMM9
SeOYLVOCnauOgSWb6Ya2cfOC1ZOLW+hwEhddY6Qzg+LjB6uD0rK1sP1r4SUF4XNn
EpkxMUYtRbkuZjETKvCooB6PXPeKxjaFOZWds3B1jrGMvYzGi0zjD1E1onJjJOxy
RxDgRBION+fKgzsF4jr6aAnqsLCV+lK5G3kEP6V2r1MQ7LLLkMFvJ/RaqmE51Hj9
eSRy4im4tPG7AkC3fuJiuOVx/jcGTudjBBTL92EAYevDn0bUYNbM35/0r13ZlU0u
xU3rz4z2u6Bizff9hqtvlyH5y6m8CmqiUNX3w8xY8odZsrs2WgnOvQ6SICvbAMxA
dLM/uoQ/3NMKNig7vg9UlBW5DeggeioQ5cO9QA5zB/+6gqYrTYDRlamrQlJXKkj3
qZ/2gMETg9xg+fgPJDY4DJTwm6sHmJZC7pdK+HAJugYh472qehfWjULDNYqP/ATB
+GHeEIkbK5wfnHmcCDZAjAWPPIIyg+sN+9/7HjBfryfA3aGyQTablDJJB0rzly9x
mULS/Kg6meE2HmQIqRdv/00Tau/HV8NHEoBekIZdme9edVMFTzFoTbMxSm8RWmT0
IO44tFNR/ABg5RLnqKoafrpQFQY2IgJuRx2ymPh5SnLONBNDokM+DDSmbcCvQwe6
HUjwXSgR+oHe9568zHyCv71oh1aL5iQ4bgsnk7CcL3rzFOL9PNyi6pW/nV3l4OU4
d9Dx6lQL2M4xZ69TkiGRLdOWdfmU+6VgP4HYgwHUw4SWwOt7HYFIknBOkuar2Q8I
RT13IRGk/QzSUShMzMXBOzSKxcvvCgZo6e7w15lYQHhJkAdZIHgSs4EMbmp9cuCY
tlj2QM1T2bscn3g4RKZM0rykYWBhK6kUkHf7JgyQ+fesYRRKOjNzTjxN6D1UbgG8
9GcEnBQiX/cBx+hKTo6LpBmYMHsSvdc+hUBzrlOgJ+v1GSC89lfuNLwO5AFM6L01
2vo0VE8ED7foaF9wxn0QbIGwxbYCGu2ofyIasMzr3wMQSWrnmVRD9JDG07mYZXyV
pzsVucoQfYabYB+GC/RlZRXCdAoRttI5pZCgcsNhprW+d9xSVWKb8WhqqOlYqoBg
CFeihdDthrAiCLKjWJ8DGt19cCW5kOWPoIGw6iP1asr1Xm+I8bjGpIptFS4r2K4B
mFQORwcwWBxpwx458oo5qE/BFrfIU93iSqKOGy26D4+2lb/Du8r57b7eot/oxYmg
miJDzFCMwV5mGajxqleL/6fK6jAnBx1+pYTZsL4YCfNUUWNnUWbMUZ5ZJBugTb3p
`pragma protect end_protected
