// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FJHD7ZjQaP1HA9udhdgMrF+dx/h7R0uVvECfIN0cNDioYsn1TnF2e2hTSGZB2Kzh
kn23JKrR1q2nrdqjwwbVR3Nqa1eKZbFWeHgri1DxRb7rzvN5rnLEVYd6HwGDecNv
J21liABLFEyGS6DKpq6lGroPXvI9JDKmXD2b+xc0WBQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70000)
JKjb3ssIdNJce3EVjkpYRSDE+capdYsIIXfSVHnh3zQoy5eUY3X9Uk23U6dKMpBq
zWO9PiQy1x1Erua4zft1V2sut8jfdyzugca7wZ8A0ji6zjITrAClm1reZWn58/r9
99DQOdrfYalH3GZgLOt/ejKrnbI+rZ3h+1XbXETE93mbVng4HoPqnvrE8UoebzTT
iaE8hRaPs4dXY4MmypaMSx5pb0gY+EGz08aLBQUUbqylscJQAkvNdR8IW3j04BdV
JLEcCpWAtxhAUpcUV8pkdcemliYdYj7VIBqf3t1BVzo14XZMKw9wctNRGuuJKtI0
HKk2jV70LmLJ0M8SndpDY8twwsYCZPCOHpd1Uh2EGHwN9LDQzmue2/U6KZYycn+7
joaPVJ7youjaRU8h50UByv7GPgkGKJZww1u4lyUbBCzUqK1Bg5r8AHm05pyCNXYN
b/eBG+6WuD1YP+dG8JGZHah85JFs2q16qCgrv51CLKK2eC1oM1EVT49Mi8dyxtRp
tcqRXN6YYM+4DKqiqgJn8gvR3gWZFRnK93t4YEMMMAXjkyxZaN9N9yN+KZVMNQfq
Hxwm0SS4l8aKIdKut+Dyy30qc/RbtWuagQNJVPXwqTH4VbOuZqUPJNzz7jpuouR8
jjhHwUBYLyHvpPlxxY9xAT/Mr5lJemTWmAixno9dtSZdvuQ0Yd9vLTmEOeY0cOrp
e9lOA804VYXBaIQytH29EnX/0xqT8S1FxGxMbhtO9NLdhNBe5UKxpbwi5yu7bx6V
GJZ9NXSJPRD65jP7Dfw8Ci4sNkoSzzRjpNyMdqJN+fo70ghqkJb4MZrsezKusl+l
ee17arGwXvACPjfIyiamNef9JDZhUqJQ5lg8sXpmk7u9ndIIiGOjn0bGUe3Dsu0P
d/QRJ/hD9Rk4NJgoMAgTzkAwEhQlM9w+kb7axGoyP8w4b1lAteWbxPGHyySz6WO9
AdxMSlGZh4OTGuLqlW2ej5wKj5+u5yqNyqCHMO/eQ8Wch0HkY5U9JLvBwACBVHA1
gI/49dN4O+jtEfB9o8GKFuOSRZIkHVH1UVyoW0hW9afYYVhT75A8h8Dipdlxj+G5
jYMPTDgUXBb852Y9Qa79oTsT/vVfyJygDbjQz9ezpTRsbYss4HtSdBP9psfZO/cN
3xdR/LNXeX39sW889Sv6JTBNfwICc5bWXH6xAj7jTkD7FdITfQyEMVFxuPMmoM7f
NzlerIpyml4FulIaZpygLXncaUtL427S6a1b94MrsuVz7oawx5oHjr+TgKtq+wYG
JLsQQek1DBJyOdlXwbyexeIN+qtUZGvPB4IZCPlUiBCmkypHFd+g0XAFoz35GqC+
PXmB9yTBtbiRF3hZX+lSlpmbdSBcxt5GqB3mU88+QmSSnAZu06rDqcwJsLszboHA
44MmKaNhynpLOKIMzBRvfLnnGDcTwV9DHs3WbBWdrnUzv9lEtUhrGZwPDk7xchvD
B4gM6vrKk5PU3+5wSksjFPgcTtDnvNWQYFgarnKxXc0cFWU/TbGJ58JKha+2HA4Y
7AxfrsPQtJM8q3ABOwFHQwA7O8PZqCrzNIKlr+b4mIPiJG/A3qwSsAJE6k0azSZ3
MyvIx9exKUvMAhgEBATCeCDKBGc9T3CL2e/Y9ADSg2jsgjEfZ9Z8wJ4y4hadgLsi
4KDPx1pm2MV0/IshnjQvZP9TTma+LK3KVzHcN0kgti5A/GB1teV26KYRBVDeRmhP
26XAB10vdi7v17pJ+hKtcmKZWp8vPWD//ulBZ4xcTCtO72lP/kQ5lGsHIAz7inZI
biWfjCuglR4yU+c58/l2zK35Q4Pzk3D/KiMl7VrvePavRN0rdkui6vzWR+eCJnb8
9glLDueSE5dHXeF34JinQk6PaLKCqQ0bgCqVLfdS+IruOyuCxHGWI8zp6C9VGrN8
nNYvN/jLIWe3T8+3RuVZd/ldfmgBjg+L1S+pMv3wjhcpj5w3V3hgr7QJtErSIEMU
gYMSLH0BVjkvp7BYtSmV7hmKDstoIkCD3vgliuXacw6o8tHyquHsqmW8cSKstWWv
Hc5B+YFUEV4qxMUihy3x5aY+LCCXYlPKSlo7mAlICNLzr25zLqwqqV0ptR2ot/B/
yy9WFNtUQeWQwKhAuGIWMP0jX+25xnbzKbWvMZgx2k0drBTveascoInuy/C5bu6v
o2t8n9cVpZUrO8tJ4HLiGq6ZESbG38yN0vnOXXiAyTwVG00982E/9hxnYkBhUbTN
rlDdDRnf6SO1XFJyQAXsAtmy3pi+GWnu2G9hVtALdNU/+q++nUQ0WrzhbCpFGV7e
r6pLzkthZ6qIiQCRE5GlCf5l18pwQC6Lhtg2MPyiHMFTG5aN/KVenrgLPO5gCcQ0
Gv04lb/BQ5P8C4x+Y4B2vT67biwgQl/K4duQk7H/87NarfWXiOLEi2jXP+Y4/noY
HNqnmosD2jgFCxcxTZEoYJs9IqTdrJqlFCUxCpqNObjcDD1vMbk7FvANI5Hct3X8
ZR+anWDcQgnQn+zUFq0gQZmyeRtcXGLRTIIM9hHS8wwdmGyKdCY5JdC30lcNpTHK
Aa0q0ht2B50Q4/8oVum3z0xgIommPKFVBb24vCLl1X+srh3gbxW5FghiVRaLXoDn
ruqTFqG8Zh8PRYlG1HhNL+xI2IUOphvXd0aJgkVktSL7Yfpt+MIlv+os7pVmnT1u
Lf6QnXhCsuYQVt1HGPVatkhZYuKMmcB0tAjjYgzfilsnxUZ+stPD90DcQg/KXGBf
KPp4KYgEWi2KE2Dp5VrckPoQo7Earp/JuV/5Yd41+vDQ8uCWK8TeVW3ja09jrGmN
T8hcK6H8NtUNFMvEZWnURPUx78rCelPhgU+oSVs5PJJlvQN+PPLDucMLcgkUa//n
vT05F2rSZj+gAske9IIVe2/azDw9Y/20sli3CZ1q+1I0ubKvVPBGhTfovh2UN8/l
vrChgYPMUXdZHMclWnoygR6EuCKY6eSLUFJKMiaxpTtM+R26B9vNQaI+uorSUrfF
nqy9n8G2IzC51pvL2R+/ZXaU75ioGCSLwBYrjHVkd+RlzdWYL8KrBy/tCKvEGIGO
+9nuza7h8QBqMCHiAikAFy76sjGi6ObKZ1rLhLHSITmyKDYPJzus+dSLb5KdOHwp
EO9B2JySZLpsTTMOxs/QA/qZrKqpXg2RZ/40dVsj8x3zElLTjoGSa6E/e8PtgiO4
/P4Qv9TNom+n3Ir0+J1lt/4kIaHzS1nBbByD5VoEgmOUUb+ZNo/lOeVBGmx8Ygxr
YaLvDQeVqAmN41AILjcZgeJOSLQZbVmNZZAfRwcsAf+Hs0qu0jFr9aWXBb/ma7yD
FHAYQGf+4H2W9bW/alGokE0BmD5FPMPYimxx+kZk9B086jNBVmyo53x+DEkTq/PU
Gdi2ES1lV9huogkWlbgExe9m39aYaBa/LuFWKQfqZrXhcLNQbAEaO3n/Wj57ErV/
3WeJatCqRH4AXyeCdLqfCoxvUffuiw1+QNMnItvtuf1x767p6f0gLW/bcCJzLf0N
oUA5oV4pIPO1hhlmCc18G2KL7CMjk8Qu52jPITzyObn9re64zWFW7VM7o+vSrkaV
RyJaZajLxexRHxh7WusBvbx6Wmup/HoRKUswY6zS9YT31RSbY11fyzRSUT3A24XD
7KuwUXLA6elF+YITZytMLdgJtGX73pf2PlEi58RRrTcAESWd3qdi4Gt9f41yX32b
YgDnDwvL7IHKY82OyN7alHQcocq0UkiE9QR4DI8Pjv8AqCyKPsTBPWRZctYQrEJl
X41ruoQ998NQOkAsPyvpgLH1Ec+FlFZ/q8s7wofzXkijxq1Xc5dszEKdm/7YD1bY
iIOpP2sRAdkPq9Cp5ReJ2dUEBXHwiuf1T2r1UWK8HKvOT72B3zp6cVyFLbpCNN19
EsMKRHgfxtjCX/Ho3Zv75aJo0Pa0QrROCwnW9IcR0UN7uKTC3BVpgSoa1Yp/tul5
bulkFOaO9GlisfQ2i8teBWp2sgWAHjQXNsgyhytAp79XeCD/rjJrZq4AcLjQRyF0
x3NAtto0MJDkniev43xyaXx+aGEhOSkBLOh5MN5uOIRM/tRqO92Z0mo57r6YuWz9
Omqtspn6AQXiyM0F6KRAtiPM6XLrfSBR41bCqzTalZAIO82qDN9dST2tXXhKIhwJ
sO38aGTBz1UBAl5SJRejEkSZ5y24W8lSQYkywRyEzrWC3dz/dK64e/1QisYKIylt
cYovIOAQgmlh0kbOPzvqsibKxi58wJplGE3TsJagUgh3d4huyeNaZv0g7ZLR/CBp
1gZaDuud/fzoj3X6uh5KerikBDBZOvQSUKciuFRKlw4lpfQiU7+VW2koMtOVmayi
xnXT3MuvRMU+WUB5578odxcn7Bjf9ZBOL+3lvbMYVod5/XygzQPiHgDn55YsnBGT
umtd4fjMhQLV3M1AWPJJkfq9pHj5rd86pPUWh2ORFUrCQA90dk3hBIHwvf3vlGKC
CgPNxR2bO/Gcx34D8FFnHkwypev6rXbBQXJXLkRP6wWGYgQTTEQpS2ep/Ut/zrM7
n+Vf6Vy7vHxgMp8lxn6RAEJ5SA/FIe8yu+R1QTVO5Q1WjWqTcsONwBqAig3Bet9X
cFiN93SPWIGLfhG66SUJbNmfJWxNZvvUN2n21R929PVjbPalj+JK0yc6vp0WFQBk
ISb/W6wRNvZOllYgLrxMkyfKv0jFcUVUzzbQp56lQyGJZcpOSHiHzSa918jpWAyv
RuMhE7MfT1nX7TCvv0xtxeseiap0EugLiVZPPRADARfvpi2tyu63GjUu4rZtZmqK
AtXWmF2kg+TVGUnQBCXao0tzYF4iqTTHOX8URWGT8Vv/rrmOgh3uBGaahIlPB9jI
P2/758LQcB1RRXIRXHcavHWkp18CW+kwdCEUnrOfp46Zg36w1Ld1yRDHvx4ByGsU
h+swSrPHuYWTS3zzJJePYqxiuJlPMXEKjwn81oFaAf05dNwLoC0u7OGH+iAW5KTR
c1re3t39uSStUc8dBi8JEUcrtSmf2X+r/DxG+J05Q+LyBEIcs8aH7Kt2Pnu+QuVA
+HB9SkEqbanFZ81P+Hy0oSqsVwhy8BvuksG6GA4Spf9+hw7iFivmldqCJtnjkvfm
n8GePfvt45XL1ITNcFBal9Ky98wXMuzd3L3ecmg7Gya2UJfDP6DGCH0QoU+Ykjrl
Mxa43G//ADVnHXwP4uyp3Bsn/qdf/jj1CArohrESXrses0HGAmvJtEWnQizR0Io7
mWKbcQ73/EAbu+Ttfyev4MEZ5pu2t40MlXlrDMrvAL7aaL7BpfYYwHnj7CjVBn/6
i3UNjuvoJxByUoCac/LdL588yOuveGiYMOtrF2GmnvQuBdXxdxmMZKubpV6M+7v0
yZfpjmc+wwXkvD9IfHd7b7BTqinNw4BvukPOljEOR/Ymbqg1ZwUayQa3zNMWUbYq
An9lEWkdh4x6eWK3YEHzPK3lnfd6H3BjDMhvdfVlDiG9N46FeeNGaTH8ePJQUpfU
/X9apA+nWzDF+MfcpLTuYSVOfOpVYmfxrpD8KRHRV1rOK5fsefQ7PZau8l7HdIo6
UxyIMOkIrB4YYE70wJp7DlqHWcRCbuO/hTPDbFgkgWze8Gg0GDS9oc1PkaMVqGYo
Gcsxqr7XrPzSyZvksUMKJ8MmB2AuzEtYsX5OlMTrz3TfMh04RSmCIsSjUw3Aq045
B0E9sURBPhTarSXl9x7UuMW0H7u8x6n5lcxXYXkhwH+ovNKhTszJ+LM7ZHM25RHo
5Ue+QL+rYA2rJNodEs3ZjqkuCY2iyKseorwnisCY9XhIAE943sCML8gXWAO+bUL+
S9C8LIlUgvvlCkz+hggLtXyy0+TZluW9neuaiTwfI2VbEgXwKvA4xeZE85z7njc3
DnJNu+scU76oJdUc4lw/oDsyHohAQ8Q3AJHGsqwSKC6Z/p2BRlBzJh3xo1lo4k//
oA+Z71/uWHyHOeLULHtHXcrvuLl112yYdscuDNdAqHwLM1mUqyIbo6BeUn+4ugdB
4/ogEITM4/5tJ8MyjOcPWbioBt5dAG6WfZ1sPMlGanr6aUrMAbS2taG6++Mjjn7T
F8InmieioYqW/Jj6tzs2yKL9s1ubxyCy0cLrB78kXzJw4fqiddFwbBPhXtzGLqUj
1d82G2uMEeXXA5KWh33y4G3SRIuZcGpSAywP4VX1Nyu/8rzuUzjc5yoDyL6MrTMm
V9WTp5rsMM1zfStz/YiBwO8reTd36WHMvgojY9ZQDUjW8yAp4nFziYh699owW1Qk
PaEAz8wePetPeSMnrIrzJVzCGu2kXoEeMNGLklVaVhaCfd4QUKRRzjjZLzc0hpEl
b3+CHP72jPcIH68Ve0TuIvSSSedwWugXRO/Rzkjxp5XsDnBsian721PTmsd1IqFg
B5yUFc5xNmBiG4TwuJTZa3gaG3C3ekpNv4v6ipuMifZ9v0uaJ1m4pxWL/j+bTTDr
Pz0zGgGBmV53IfpRRIbOTnGWP3bMst6Xk5p/FZDjxXpHpKm9l/uaBHQG6b0y6rK8
kf4uW/j83MQl9WPlkUw7j+Je3vt27eHq75SIxffIHjAuiwYebCViCk9SEFTwFWfW
sXtd/WI8xTHg2MAc9WzaBi+uflcvyH421ChXkdavnaIvGZKbFaVuHyIEGrDZy8Es
plYsF69FMwryvRD2dzDEyAKnH8kGKohh5yFEsSvVntCYjmIMYIRnRvo8v/IGq5W3
dWEvPuVy9LPiE4qVWHvGJQx2tqrWI5/zZtuuAyzkLoVVoow3srhZCM3o0hGDlC7P
77hxD/X6FsLiLsyk2Zw61paZDfPTBtjHo1tIjbPKRQNx2OpOopFsujk4+mgf1G1m
HImJlR5Bgd5JgKhdb7VBBHzVjpDB8DKZTLQ4c0MJgree8DCksQGQpA7nDBh1h3lu
GUoYZW9s7mVNhqS6srRE54SZ8r+L4WQ2pghzX46ebVl3/D0B5ba6a0e4MPpyJ8cx
45g3+bNQURz1QWiL+2xDEcPo4jWqe06/RdyG4YRKNzvDb33M4qD0Q0ctcCNi4PlM
F7EZyhK8s8fx8nEKP7G19PhAWGCumUGw9pQNkqJnoWyaogq5w80eMwO4gJTaegI6
vIsQwb+xtLhOeDvqjZbzcOggoTMcyQGfrDYZt/RtWAnaDDlpsO4qEiS2hW60pumF
qdDOpKisjCuzksxqEuKgVOVrFmikGMF8nzi24eMDvowkupj86eWU1ep02NVhppzX
AW17TfvyN+SnmzK4JEGBBFS06kpjalWE16Hte1Ts4m9YXa6vViuFjkkRk1nPZqZt
VkXJliiMWlC9qfk94IBeTYisx7FYHqNUqUOPU5CkpdQj4dUziOCX3avTnNXssY+N
RilhFWCSu9xzAY0CM2lUJwndZXWgwGzN5YVXzYIesIFvtF9v7uHzhUXpbOzJtyXi
+Acl7lM7WP2gaMxvFDXyGdZcQX1txy8yqAKPzhGrBxCQnf5fNXZLIjURlyxCssNg
EQV89qsPrL1UP1iX20HFX0ZQr8eu2nJWDvP6DyLiQqWBYpt3E9kO2IEa0CpaWBjf
LK0kxOXa8KhHeAP0ogv40b02HqKl0KePoc8xW3SgnFdzT9rnItDgCPtJfC1B6c1q
PYoF7CDt1W69VTmnYu1EAaU3Viobhpnp7DnnVnz+Kh12N499DAgT2IrUVg6Aoluz
tQr/gDNPEh/wJdNo8H52aWfBXIxQgQimm4+PSHHiJG3c0o/SPQ5Z7i5Bh5h4UrVk
JMgZG6CaRWmc9c7EEBf+dfVV+aHoZkU3SETZAlxmCL6QsL+nNscWP4QRvmkPxNqx
v00rk8AuDtWfVv1En8MxKUzBbLlcP7bes93ELTm0F9XCzfE1qrWni9tA0XjEKDmV
1QgVEIKlJCmNnyi20XLCytArO6JmJFhXrMFQD3rF0e1TWAsZ5Q7oo39vbWHgqCvu
uwvOFUuZ0eWOlSmGk9yrybBZRajHvQBA5+1CgBqdYC0aWT8DhfH4ax7ZZ6/cCpA8
NQLoIafUsEExFTsA2SS99kD0s6FZAUxrLzkED4/jT9v1QXw6XtK3V2EsyMzyp1N4
EyneSbqsD0DGH3M1mu7MAXqhQEbTATLF6YFPst1w7e0ozMiqyKZQxR2hWpueBlWh
Iz3wYc5va6TFkEtMORTfL4t6kYxNbmV26IH8DIuH2GAB5nGtqYdxmM3FPQoF9gYb
rI1R6JfC3XBnE3mcf3fHXOLnKWS1QhsgBADe+tKETfT46rURam5g6DdwGHSOMwry
/xoRrE7jjY9i9CKgkpl6z1/HPauf/lNsVIVVnekKdud7/g6qZJdd+oXP5Lcz5hyj
lSFtHV01BA3iRj5Ne8JIk0++ywso6hH3J85Wm14zEGmt6sl2f/QtGxtcILpX+f47
vr22inbUsnVf9eZy3M5Xjb3WC1lShNDDPy/b/tO702Yml4nr/zbvUBIh1OqzjJy6
dkqVLnY+jPybX8MvYfbbKoCLv5lLFM9ceNGIeHaBVCCYx3PxsJPScejYMQeX/wlX
FVJ9f2aac1Wkkf0R1WbuWNTLhcG2F1SgzJW6Z/0XvcSJBKXiKPjnFJMbjGe9mGw9
ksQKIOALGss/yRrxYaNyO/eRI0MDn9t2pi6j1LOuNfPkxomuKPf2dhSoxVRH7ml4
MWe5KJH49v9pIuUgH6J8rSuDiC3wdoeD1kdx3OwRgPhHulECPA3YHrGV/sQPb+X0
Js/H2QgJXgwwtUhCfanVoG/2kIuLQ+yimGDmdK0WpXMezx4knZbJNJhKHZpIcO6p
Bk17a7TQV+OoWq7g7ehkaWqLh5vPzN8nx/gnh3OhJPJ7P0DSKZOBGox1q1+4dJ0b
nZrWr1RL9GeGXcSCSvHHVXw4LYJ5nSeNfZ0c12YGSh8mDqd83DFxfn26/DQiJ5oS
buxUPfen8SYJvKvUo084vV49s1oHT+z8WS2yQu3WITICMg+izQHOvAY2F1BGfP1W
o0rRTQeUaa2iQuXApS1oT0KG2EH9b53xQgF4s5ohsog2v6xkb9H4AavyoQruLcaa
eBfKL1gVf2OWz+DwS48O4QjIwfbFm2SQ8tsFlRhY3zI4VoAD0yX84DVYpSc+Ztyv
/sMH1tSBwHCMjJwkVDmHqFOeKI9u1/mdDzrkl6k4fglPWuCqdtYO15eN8cmZJ+Ga
2hrx7BB5kRxMNvJPzwN5TTDX4VeUM13W1lFSNw5idN4BHP9izjT5nY0Wcl2M2VUr
lca5PXvyDFbaIHiYIFGIqYaRNhDFLHdurhuWTuFabiDRkfFHcqy8cQo4BqecncgE
gPkDXWxh2l69HjgXT02LKUq7/D6EdUOY28nJrNmVvsxL2fU6weg5pWVmEhxtpi68
x/dfXLkrM4XvsqYPQ5OaCC/Uj/Jqh6eg4igPyUVNUl/Huahpha+kDZo+s1Aytb1/
7MPoxPAJlHa58496MRKTxgKSlBg6Powq41Zh1StRsqPvAc8RBumdm9aUVDMdus0O
eWD+mfSOpMbECvMIFCLyh4bhLF8Id1imZTx0doMhTt1X5YszjEY8ALHwLg7veOe8
K/94BQAas6ZH4UmWTEdBe/8nrKm5d+oW9WhxD4Q1UYub3gbTW++y9pNg8Pz+5r6p
2miWPInt39QQxqhf3hKVJfLd4eq5u/iZ3vswMFW4Vh4s3GVk+UfaaSO0gFh5RcBx
UrST9DkZsn9n7huVIxactPqSeh5DQn0UCaQ94kpGYj4Zm72hcPCx/WBNVrwqDGQH
HdQxLS+BANDczrtVGjNGhFY1vF4ZpWXEcSEr2ZZedEn1JHvaeRvr7Ln5/VVUeowQ
I7GL7rhNFY3jCwzuCSNmRCc1MdEiafQivj1BDCa9CTTBexg2Oestr3cw32v8ouf5
fe0FbGJHi8nJ6fC+i0WBbpsIe72dsIaDq38S68Syc4WCjPuN/X1l6pb9T2TlxZVd
nTTuN4ZottXOKw015488HGJQv3XUcNRq1XMru5zi9qccYM4oyf1dZxbeZa6+roiv
UB+vPOis3tBztvSLcc2ELz+qbM/jTm2OOz4+C4LEgWP9sn+JbMdJ/PA1FfuULbpz
4YSVnHJO7aeADsHfTX5E6qfyHXXa2tiQ7uuSPUBZfFnFK46Q89BkjyMzQgAgnUFL
2FFue3R8sss3dOXrbX8ckEwbeSFLQcqn2cJKMfjx34J7Avue/YIM5j+WkiJRwihg
vkcDwUetZoRZF6hQncB7Z+Tsvuj+65AgnStbI2BTWAExTsjSGuYXpN/YwK8Ew0oP
17OOVzl8RQ7IxsAEjPJu+s13+D0Oum1bkFWBGn9dST8XOi1XYDHLFw7QTXi2sMG/
L2qdhhkyugGOkccRW1wHR5uKk8d4vNiBfFIGm14IJDkjFuBG49nBc1hJvnYbgGRz
l8lV6B42qABaFKueHyJgvpIhwxJLfOus+2OsaXSvNETs07ew3X6whp4BAEr+2mfo
gXB3jmNs39si2rcVAzsigkWjjtpKJuSt9HPBEyzxBqgr1IQSMVweMNJCbL080LY5
CidCC85t+NXUN/eTY5eBVJf/LWA4/NwTjJ4mPpKAbllLDyqsejK/tRLi3wWSW5zf
4BYEigKo6Z7VITuV0icnzGQNB7ekFwhFJBQ7cdszHRmhXGIyLyRki01Ucg4TU4v4
+zRhdAWxBXE6T+BZNxA2DUS40LH3dSCXsH51i2BxJxd/1Kqmn+djTA6njlmkntLl
f2W6ADqBUPwTxwKhNw1Wl0ighSdR/LTu6DtYsAdZzcjrEwn1DPY0robxB3SK8jUF
vAYNMnZCJIvLF8UKdF4BkCjnbVncBu6QoEvF/i757ecCg83j+tQEQ3erhgskJcrG
nAJ/Xg2u12F2VeLUSzTT1uryVaslfYCdjSKusw6hPfXthEq7ahkZPtzMnfnK3JbP
Py8cjo7z+ilm+UL86bw1ZayWkCkEYz8jIalhlZptHP2cYbHDiwRlo1bpTbHh6CpB
bPwm6R9IsYMUElAl++1jHrgZxsbivbZMFAqh/Tgp0qpVwm0thgqxozmroL/tE0Ce
FG7U5/2ZExtaf5f2ev0XR64gTodqWGQqIjavLKrj9l8KbrbfUfM17q8sN41PyB+7
sGGH+nF6TDGWh9Y+xCPS3Qiu6l+dav6JApHE7zqLNEWHw83USokspqB6NBMe8Bbb
1rTh3agYABTGZlMFMtP5ak4zLjKEHY43Tvonk90UkNOdytRe4uooowbtlWDrHmCi
YeFIHZAX+0fBSP1d+MIGNchrYZuVBERqKtY1FspCfWqHlQiq+4RUgwVzxfmwBX+O
mUdJ/X/EZKjh+kmJtbN1az9y9RWHcF72Ec/VniizIA4ZMw329+089lP7Lg11CDz4
XE6Wf7RGQeirDAeQV/ZZ9KkrTe7zsMh6j+V/LQxcAN8LpAAsVoxo1V6+ogmDS5pe
3y6eCGnGkAim4ObV1qnxrkOF8+EPlpMa1piLaHW9aEWTr6IJIyjXhymmxpndW10i
pUsoweHsPdz8fHXGHA6Fzq9vD0xGfQvO15mwrRmhMybc91kfGB7gokC/PRioTeXH
BMHmDek3UvA7j8PZmSDTWEdzk0MB6i4/AYebYd4uv5afsCtoxYWLrKQuSWFYKtpl
c7S6AC1MBHxV38acEc8cYYCPfVlh0eUI777j0qNOgJE7oQuyXmhvwWGp/rPdBjYn
V3ozqFRCJTQztIVcWUac5ZPak1RKkPYTYupCFNu9j4DCHfKwVGwvKZ5rJ3rJEAFe
lM+cAq7jO4TB3Rd570imMyUALm80DthKiGOVATZXHIMatXIWXyU6QUZD2GVL7i1+
rMDSK8zpd3PgPliJbwVl5//xwJ39vVE/rN4xfMds5oe2tEFkq9ORpQs5rhyxbEb7
QIe99AHipNqMwt8XvaxAkxXujavMXJbUZPHXK9GINKym4qfdYtdpzcS77XXkp1XA
JQHd368J9NqOqrUS1tXEPvs0Or7N83cRLHEnfXOIkdkOrEzEYFYPKEXNL/QwX2CU
B3f2om1cIPmwt7yHDpkSwiiA/KPG4im6vC/QaWgs3mCCh8yaXqav0vXE3T133IKQ
EmHYZxxfJPlTiaCbvZZ6af03ccVmcoJYYOw9vnqRHoxFHaAg284YFw2O2jghbuq3
kmZ49whKsdx/vtsenON8s0nkCfyZRwnIvNTHXu11bDU3m/Shnn7TmrAQWCPHWs+f
Ce8aTubC8uiQIJbycc2/RmkSsvJg9VUjYwJ+jtbs3PK0+QwuIW/8GfqDerlnJN8c
B/mg7F19q+UhOM/tpfPQ/QgCxnSItwqOGt6UQozz0+gqaTOC9iFhn8mBsk+HTw5y
D5jvKRvAJIo3lXJI0poeuN6eHnvNtFwIv+0TZIXmEYhc1qzG9/gc3nY1Lg/paf8g
hKNELf5f8pU2E50YiFPqDw+cYiukXM5nwdgqalrjpPa3hfNPWa1JjiZZCTmF2GYS
3rSoCd3e04Kxg2DUfaPm3hFYAZ0gzLXGjIuRN1gnwy17FVrBPMtEbWxJl0UUqxqh
CEfc5FL3F1H8JM+tLWsTq+JCIsQQtNAQzfnXr8BW/0Fal/QsHkKzoUdDf6rBLuYz
j9GtdZHU4fjLxGZrU8NxjIvzh9FQ/d3zfhVCrKLq+LEd24yxqJwMBlYbwyk/Obbc
BBYolCnrhnDcpp26mF/3Y0UTbOz6QO/lKOYohxbKyZX1BbVBIrlBjaDEakRAkvfa
YlAoYv5JqwwizGhmfg8Rluq4Cf0xx+ND6qYjutirRNfNAbUM7MaBjTweClilwU0S
vC5pssLQld5Nv63Z4vl8GUz2WwtIhDyfy0uPNXn8UPoVUKfTxrQCN/d0XgnMQwq8
z/j82SHJv97MzUBVMoPa3DSgcANfMrU1QQaTIQogej1mWtAQHGynV7aP4dKKYrL0
A9dsxPqi2xJA2EXziMolUEIpIjsQdGInPsLsvUU8RyC8tqfXya2TFDlLcwQiJggz
pEAlxODNxZJjzpX5YyUG6KduX3hAfbrhuHslOKw8FDSzM61gBOF4ANbG0wtYCPwX
1Q4LGLoy7MLwU8sZ5WZ5kqraJwCRowpJDrN36DpVJtIWS3z4PdoI13RTC6Cv5Ekm
FdcpXxpvU8b33BAHowoQuZD3s9ine2MN+gniXDELy0ybkP+LwuTWGZev6VpLzJ1b
DB7P84eSiL09LMYKfUwKEPvbPyM3qdaSrWXXax/S7QO2Z7Q8aeWoqqwF7/J497CO
0jufl0+y8rK9+rvQDNjan/yBO37yEQ3diekPw5olYgNh6NVwLQ1VFvAUInIQrx0l
oMNLFLMhPb0PT4yHEcFZQtxU2w+NxpTazrJTa0BJLuQBnAxFvPw6EeSb6rteLFlE
L5RkLUi1gF4XBbBmxoUL16YeWczPnrfprEb5aXv4rt1hOXqNbfC6Bz908tO/NFxt
mWZYA1/FskYRtyObyO3wCRsF08u7S17x4xVx7Wwax7HKf2IE0RlMouh7pkrRd38r
dGNAeMqX13dfpob2md4RKhBBCfOU/vpAA3ReRAd9FOYO8I1xspb2ISfHopKB9zq/
NOI4nTbWy1MYU9D6ExezUToMIl9Xvczjkxyzmu3+LA+aF152FUn6WxZKXemayxm5
+9L97W0k2jJFBDJKHT5gtAOHTAowsCUSM4HSterb6roouuMWLjGPwPRTToYaYWo6
wBGZXopZYvpFlYxCBdkCU9R7Nq/Uly5ggduCywcE5P6ez9nCic6eeLBeQbb2hcnG
WjoCJoRVK5UFoXkyH4j++KzGcS7NVVFOVzGOK9LHmu0UvMS3eiLxd+RR5pzyTczO
U1Ekm06sr+90YkQAPQWZhrl65Pc8mIIi7g6Hmq/6SOM0JV/4JEyALnbV1P7cF2lW
c4Wu0RisWvNfXYd1H5YlhHU33/Ihw4KDYRPnaZKdHWOBlBL0mXwItfmCbr2+KHvX
wNgFjIOQG6FTv8zibE0sh6bKzS1uvwlFljpjCo+Xg6bgATYFT8UznryYAarZcE6C
keSP7lNUDodu2RdFfinP0Nr/0BtTzHjAMj6W1taKGi9gBLeZXwmc58HlNFMLh18F
yz6BX/i4qa4xs53D0zVfujnyZGsqodrqCRTU0xs70xxiOidpeZmW2Nh67UW+KPVi
FiVeR11CHyVVkIHTsSGx5jCAV3k7SbyX67+v/M7XHFrUbyCNcUY+rVM3pY35hYUb
8nbweI8Qdsj2Hs/Wr0Xptk07XRqS0rkmkSAfXFs70lLq4Hs04Q82nQnZ/BAmoEug
GPJOTvGeXp8t4ca2eFP6hqKEq+HzSG5yukrXFN96p5ZOuang4ISIvvDPhRPN4Emg
PVEoxLpSvtsHzUo7ZxPivgpYrNYyzMcPooKbHfLgcaZCO0ZciPIyymAgF1hzc1BF
wfgAAhwOh1dld3qXfg4ZiMzvI9VLUThwBdWPLV06aI+HvaszLE1G9JnaalQiegxu
k7Voy5a/L9ob/lWNBtCAUEpyStBgBQn1M+99HjywLwgUIEQ5bxuTG5MEII5n1Zz3
fVpgMQW9l7Z13JyBcCRcRRTaQV2WuCLsX/BM/DziouGwLzaZc9oXVRDUX6D5r0op
EEcpVgh/1wPo0QIGH5Lg2yQrA/u37x9kB2DNu1P+abAhwj5j9Z8j9YFqGcVdkAgB
KI6D3m1vtGuG6OOjkxhlDB5EFatPQIVPHYVhNE09c226CRNccyIfK1ONsnxZG4lL
DRwqNinWzI1w1FjYOGvfdpQJ2+S0byGKbsoql04RPuMedtdubfj0FWu9nBaXpZtF
xYClcJ/JxKUVPsFgndYrP9VuLUAHSacbVK7pS7yXKulj0YmbBFDfHJzfw+gwNjiz
mLJWTM0tx+0uklDDGeoSmnWIWhK20uBIvmBJUoKqwbZIuGufGy8ZOc2DfI1cycpC
GnfKVaxOxnAihULqHXfK2YIXhvNYEY8aeXuSS+KvqW+ja9jYUbBur18LvUHBLeDE
Lx0naX5QYn5JwoPzzzulThEuDPy9z+x0K3eSV3WvhvLvXOvEK0sxMB+y3VIrQ/7P
dMZtYZ/XnFRcrJ3EZpcG0nEsCClOd7Hvuy5HemWElER443DPMDPxd+YzvkWmA05U
jvVxgLx/0mGHpTMIbPCsO3XeaySqfsTUkijM3gQpeJMUh4NR7dpsyYGL0HW4uP16
KHv4nTMgwhlJ07Cpz5WSQqFuwFRYeQlpaqtayJddKy2iBORQxZvnSlIrXy78F9i+
/F+G5MRgIfPTt82xc1mvvWh5mFInjrPHbmJEZQRz/4rVNVTk02iJkZ4RzZgCqufs
fwIBrYs9eVYyKcqmN/kdzylNJBp9n7Syu7PMNLt/8uBenKb3bHV317YuatNrhd09
Lbzos63/J21V5z5AZhFLmfzK11v7Q9J4ceD78zY0uTZptgD+SIp+CHOAHreojbY9
437fKLwGZMb5KAJLVbUEfjPMH8vP5Wbn7s7S+ZTYAlCbl17udZWVnhdjy/GX2c8e
NxbEGFq6uIwOOSZO+82LW2V4Hfx+w/nYcBr60YwlScnVHXhOr8SUN6+uw6xI+1jt
Aci3JnBfv3mnFNMZDp1CCr3myoDSO/F2rQ8k6avhTDI/0CjMJuRqyke63z4zk2ge
uw2mdAOrREjn5uwEKFDjPekj89MNAEKD4POyCEBQ0OGISUULonOb/ihakwFx20s6
bMzx+6jYqTrICf/LfEyNvt6xNgV+/CwAHJCJBAji+qTCh+ei/7nOp4gUKm4IuM4L
CQSGiB9LfnRJjEW2Fq6ZjGxZfYvNSB3AVKathrKgagKwXpvdIFXVlE1AQZwkbglA
bzWXppypcCJ/D3RvdOVgqKoNDaFoXG+q/jXZH+41I4VcDfk2Fd8aVqfUVqsqSWd0
brYKwRcU3vRWNDYXBxOVxh3tuvYsrh9aNT1P/+gY/FzevuDZaYHHTVT9gm1acWsQ
pHON+ZfmLVU0bSsDY/1qQHbKiVLyiCtvGkucoJMavIefoJ1siooiEV3Lhk7mk0vV
IjAlDT1tmhRHX8Ttl/YZzcbX49YnhIk7SPBigznd7P+0jiHcPyFUdmLvvfsBrIOl
4PmVVEZJcqoLrbLYHSxf/PgQjeqL5JjJeH3GNwc1tgC+UwOcS7g/MvTnvqTixb9f
8LnlADhsPdVUQOm+SYAtIoCvxgTGq7OWpDNkjXN1bmCCZjVKUzYkUAHS+cYWWOpK
UKd+YSTUWiZ1GTJOtlIeBYktTa6QQRGqMPF2WQzHVX5VTY8cK2mcHWJMbV2O3sb9
4dVDKT/QKb/fAL4U1uql/MoWGiurOaDRWZudbXb9iYI1nVtXGFmgNwqpT91YFRsL
OrSvyPKn2D0uUCU25d59w7pk1YazT0r55Bz+qhTLk3Dl5ihIBsb0MTUghvmqvrd0
Tu0dKp621Ju7+Ok1fgML4X4aU/D40uTXtUNpjU3l1O5K4s2NfWfzddXuyipyT9Ud
jExdImkJPSTeTiyeiFPyvloolb5AKrvcFv7TnngGey/CJjGJh+OdUqUpp7jkPUNj
5/5bT3Kp905yXtKCkrpDjzld/yOLU9oR6ac9FBBifoaW82qNJDRJ7nw3U1ImRZUe
8tJfZz9fqUk2KzbHOYB3ZbBy7qJeKFfvCTlfnD6A8F18cFmH48SPnBOIcMO1HXrk
IfUR3VoK+Y1IEIwTXTQJ/EL/8h3QGDkQeXsuBDk/HFv+IsKgZQxQ3tJioNrGgdhD
m55Jdgst1VFjAqjKTYg8PawjrHiObTaItY1lD58N4gtgUl7M1mIey+B3I7UjPf4d
cYIHWQ1/eTiNn/To8yUdkRNodsUepypwwAq1mpQ0lnf+0L8Qh1ZkDskNKk9CbHB3
cYB9ytnrZ/hRkiOanTiJnX/n1A+POl673l5hGrr1dYqLZjiBIoKviqmAf68Fq7ZJ
WxtCLD3Y3SwtllGG1DIXXOksYlVQzAIvDLSgNT4OyEm17YNtbYMBZ1yEOE5c68Fn
YuwXKsX8ihqCWOOgw+jO8fszfH6NR3q1ev543HLx+ejVztVbpX8YY5z/U5/hEx48
A/ej1kkge2hgusSY+LeLG0TCdIxfRx65u71WKlMo2SeyxZoNmhUM3EjMB9SQvS9d
XE9iyzb53Tl/nwEoT8XHxrcfBzd7txhNfl2ONcTyooU1srKpnezzL5ewjKCbOQRI
IWRi/B6RrPJ0TJ22aRuPjhlTHxyDz/hDpPtjpPgUTqQYQsoM10vaTQCcb35n9hfC
Na62PTwo33yzNSzzVI2J2z9OX/8d/kSo52wgtYq5AuVz6V3Vm3fcME8z7QeXtxYl
qHc30/J/xHrYXgtA1+acrtm0GirfBc2J/mXTGn830VeW18E/5XV13GcdtZirmWEk
oiDMAd8UhmC8qH4AjRoR6otmOkCurgt8s4Ahq1GMngjG6PG+CjCL+5xXrAo97Oj5
uFVYjWVM7/HmTumT20BQb15v76zLxKpf0Dv7sqNf9Ca0AfEexQiL4Y8VNrwR4MP3
I32hh2K7sO/bzyWDOkY77lvNIocu/HPYoQzGQx5byxfNEVETUhmvHg6oXjxN6ZyP
NsBmHkYv03BMzHT5JigOR2UQf4bpc6u1SmyOlE7UfGOMQd8n+BkSFCrzlE9BaH8z
cki7k5GVegZDtMj/yZX0plKHVlxxPdX7LT+X+F/+oc4Fw0IPch7Cumcn0UtYJ6jm
41GUjHS2b3GvlmI8D1zjUuXzaVYbE343SXwIxR+lVW9bY+A4BymYDTdV1D23y+KZ
V6QzIABg6UfnZMeV3aCEFBVNw/T3/bvkrETIJIZLeKR1aqS9WnQMJdZjxppjepcF
OJG49IhoTZDUT0S69B4bhKMTlMm4yqs7HptgKd7HOLAlTCKpg/4OlinstmSgJBPX
skIl3dJ7KNtNjN+k+9zl+awYc/52MnI0sZpXr3Lviw0JY7wlZxXXCUGBeSYXxqaL
QG1+xIMmv2lAcnx/Qxs7ro0M/sj6dB+5P3whOKaonRVmfDBaB5HbHI6qwUSJGAY6
RgfuFZ/bG6R6nthltTSUa6v8Z6MRFYZTQhiGtOPFOVuEog7iKCl6dPP9gZfc+Xpp
D8hHuZa3UFX+Axoa/lPb4HwjGKYO3o/tP20vXJLFu9uy6DVUbYJh9LQzqEnXzpqa
4fFCpPkuAvZEKPmOiLEGR8MJebmJm4QvlBQb+S9IMpsAr2I6cWm0dSsLWQH8rer1
AzgjV2R+fsO6vluwxOn+vL+CuEW3+BAzO+IrcNnib0TyueB9CCH+egzlpJvfbnxZ
m0fHvUiZCZC+GBlRuN4bp6Y7smMCitAsEYnA1rEz42rqs5+OvV7yUBNYEDRwyttI
QxCPiWP86xe+k09bIO72vjQwt+Ifms6/hoscRNnii87UV1Wnih+9nJCscRK1gA3b
eU8in/YFIvLVGHFrUzegSx+8WcA6nTKkNksHF59OIbrCyddfDGvgQqPIsEXGFxy4
pbTJJgHrCBbQyuoHh9c86dbZKgkNxum0JRuOLe2dRgFHoFwz4ZQcEnGxXI/7Ztix
NFC2cQRnoNEe1j0+0IMAeikm9s8fdVaWpPxFrfSAj9GV0goyaA7qR/el0HFkRElX
2v4Yj6NKhwiHPL6oHlMnjsTsOWvZPpbUsZ4ZNZ9RGqIzx+BeejSmlbj6jsvOnBCl
2i5bXp/cF+hs+m02kCXzaqwlUFJFn5S7ZRBTKCFJNGYJfwAd6v27Vo2WqjsjQFl3
P5OzooLv8yIkzWIr+e28LZFfp5WluAPaC7e0h9QhRy9gw4QVApTNnW1oS05MXFx/
6ehVlny7kt+auDG9P3N/fKGch3Zlo7Rr5tEx6+y3j6ai06xrwyEe761A4ajzHNsv
X7DFadsfXJ107t4AaSXBdQ87XE563V91J7jLt9HwiK6SpCEdLXeLEWZTlpDXzFfP
u5tmbjpdc08G29psxNIDkHAWe8Ft6ixlbeWfh3shqhqJhFaldERvKEeQmzFNfTnt
uGyn4GzLwB4sYVnNKIcjuFy6OEgiKOPMgYdynZe31W587GSXyf3BlJfO9QPfxNKE
sv+qbvZnyZ7u0cbqpKjD2bIE1+H4qCZlLKiRKjLgiSCO4PIdALQzultDQs/2/GBj
dxm1Bg4ln4Y8v0rAL985Kd6DqZgvOrzeMnQqRosKjVDZY65fHkwD+ubOBeRxlXTy
Sh+k9SmpFjStVTff3L0Qrps3TSShNrtZnMCcumJll+hC8UPMUihybpgd+XPRbT0g
VHzOSLQQkFvtOz/EXvjD4imOmaQKM1+kUCyJ99w0shJcjOOoGq6tmzDcXonY1t8e
J/xw93li6ZxfYId5xDvZ2HatqqHbEBtrRoP/vnhImF97G9dRWxzdq+r+8fCfe3wA
iHP6pZKa7691Va47cTdO/E9CUFF02H0nnu32qiaZx0r6xgnml+IQv5Bpdkx771qz
p/RDBZlJ4nZ9R2nfCAj5A8cB1nfyHLVxqF6zHtQyYCYMzaWmrhtvA+xYulVBjRNn
p2gcVZpzXZWbUJIWC512SqAE1VLzmEj/v36Mn+BXIwM+WkfjPyztNNXwBe6ez61p
vQ0J+P38GacEe/peLSSp3/g3x1O8xlHON7EtUGdWv8PdNloE+ehc5veMMxdZynPF
kdz+WJWJLCeSViF3tNizSdbUHV4HKLKWOIDQ5bkZSYbA3zeKvxIl86hLmVYMyHW2
4aLwffr7PAi1dZEFAMz41cECuzC6A9pTXYe6sVHYOkGCXS7bjrfjzM2o66DnTmUp
WSGUSSQNH46C9ViMlKQ/60xDAw0vT2KBpZZZSbzCMvMTLSDz7Uj7M+/1tm1dA16i
ihOJzUzsua8W0KcgGoys3sNhRVyXtwa2hPdpQ5v7ZYs5QL+Q4bpbDyytlN4IKvr6
4m+Ekundy679CIRQORudDspL3SDnOkiT3mLfWAiXXVtkmgk9Ur++P6xEr699FUtj
1BYIrxOSfuXpa+nXLMY/vEjxfzbLC10mnbXuGjVoahvlmRqaYB/FIFEgtdiIukdJ
U+ybL0mgA/+9gRLQqgBVrtiyImi25wamrlqhmTsawNev0hqRImoQY0H+K/ac4PUn
cHsDdQ0Wed0XC4hx+Ue5QHACiSESed1vh/Tph25qXFR5BXTHbv1ig1EWuJEI5Qjt
WxY5UGIA0rabgzjO0/k61aAL00969oVOZvqdNrFU+Q7R4SqDYB2m/ubqXveGtRKr
xAOspbsQnLrZnshjR2sGNkD74vCBVzfT+G5CReGOTly9h0lMDM9zYSxPMN1x9lAi
bwckTEZDZ/4Gb1hYvWC3hzY48fnKqCFEJ1kOY+2Qbwb965rhOY3svsYdXEzbHWOg
AVezKTZX0BiotPVHLXfWgBPCmLVkTmfX5TGWe3zlHWx8BhvgBGnfpWwub0ARW1XL
0jksiMaDaPeut2DPk1D+LjVmSLtpkVC3I05IU6DcdQp9HfeIkcwai866RePnYb1Q
AHxSh9BT7LMaxn2Cq81lM+euM/Wa4UDKKca2XkH4DScscjqN9nrCXpGg3RQevUEz
jj57UhdEj3L7FZ/N5tCB3YOgc0scQNNWou0YhYYFCBI/O8OzW8W16X7ZPFgg+vtZ
g1GWcdWl4t6TWeMIuvOBcR4OXkCnZYCy/5YZ/KHJKZKxfQ4RowhbQpR4ypqshSjK
XnastX1Y2s118A6R8nAkUQfJL0TJodqguQvp7jE6yCYd5f7Y2p37sp/1V66fiJpS
8ppFDUiCADBTy+pGFcPOSm0a7t7X/Tkzlmph/f/QPKUOZmJGeMU/eX0zJti+3rjh
VoZD6gqJMzmyQAVQ93I+V2JBH8kcQ0m9OmvDby9QOTGFSVINyFeDSi83KUZEh6TM
t/jXUcTzDDKH1UqyJuhjIwQVxn+dVlZLAXxDsQpSd8xWoB+h3qEuo3LHbyOKRuMk
XRU57KRWpDRJjWcZ8qasvQzErYnlFFrxmO6hT35xGAe53+RJWKtU99d62E5aNVgP
QPot2sQ2BCK3l1TzZqtC9JkBTkm8ROqfinNZ8DFemvQffAgXExoo65IGtXGVNbiq
g4Efdy+4xiuWgY1C+h43qBQ6KgqhEvJJsX3V9fsbmFFlnaUiEhL399BAHP1QCUHu
IlXrQYfTxZt8JoJ44GT4Y1QJoz+FPN6q/itMxFsFe95SJzP4lXeY9/f/guWqC44R
f90C3YnoWAQrdkX7WmpqNDqfhKPuauo4K9Wb945JvCZ610AaI8A82x9dMPuj/BsJ
98Es4VszcC1+UPC/1b6t6GkIUYN6l5/PTJM4MUGUkmb7tq71+CsXL9heZcvG+5mI
3vOqcUpXTQ7aayPY1cAedaxFnmpnadhGrFRmBpGUmrCVnyTFSFmEPUgsuuLdvLLe
89aVLDNFx6MKCeNrVc4dN97wKOl0mExZ6DtqMoazRdXItUSWNeOq8q+CX8gmTYst
vtW5NPL7RqvWdSmKEZpMwNj/gPIfwUmpkHYYN55YIphHn7DDdYDvvCNeesL1NdKz
CQscUoahw7XhI0zgeQ4Wb5tisASYBWlyROQqC2heIq3/eg2wO0tEBYToWiDo7YB0
Hl1csudlRgi83hejaG6OkLcqkJ2TO4+5lTgQ+4SXxGlQjQhw4u8NBsLCNwLpCbSD
S2fsO5dvM7sf/rUc8+BZu1fv4iPTHiLT4X0iKTAJsGAYS1BQ3T2D95jb+NOAp3vO
iRI56tTlfOEQfMTCu8a8520AD/3qTOf3RzMOHWAMfHAZ5U+Nb6LTbh+lUsHeh+IH
g4fumWm61b7fhkjPtu6P6XL135yMztsU9no4CWZDI/o8o+wQoKD7rS+LIAdwXZwD
ucRTwnUy6JZ5JzSP3SGV9AoakcHZCoH00gnQ9NleFX5Watqv9udBcIwsbBVAdIRX
IAOHgtNSGrpjCHRCRHCeupmazNUC4ILw0vZUCc72kVfplCi9m2x2tPNOpm8CzV3i
5/nJtkewreyieMW2HVWO7YOPvQoZcwoctm29b6rsoK7v6wQ05HdlS8kJEfNwY+Xb
NmVb0vHqgBqj7+rmh69XpZ+BKZxHt/q07BSMWMP85bkZ23CJhIGYTNyflwaauSnM
A5tiXmRUwqrWAIDYyiuF9xkwbbQnzbdZ0mGjp4CfSlF1khqsxEJUEbL7pOk4aR2h
A2NAEZd3V9eKMvbHT0y0zh7V5H6S/nysfXK7u0VR0dQlzlYHGUl2f5n5HTaV5F6k
nYSSnb4z8B/E+SWDIaZfnpezOQZ5ooh3lqaKxmjSPlCQ/lPWRlGr5YuDLX/mAGXW
1l24FGw+twsyR8il11KW9u8ouLLPG0gtR0rBlndOpGLxV0ubMk9MJbm/b5zO4n2c
WkrsGR49JjtpIBNkESDC2k8vP9BFQC4DKfcm9yxPalVtEG5i+b5mRjoRsV6Sl5aJ
suGBBVfXE3h1+QY6ZC/0WrhWjgyyN6ZQQzI5r7z5auYdboJM2oIns9Hi/H6a8q/j
ALqLkuZP8DZeKM9csX0Z7FYkdj/iDrgVE+Pk/Jqhu8a/UDxhWuA5oGKaIRnS++zo
JrB6wQeCwfudGSbjEBLB4Ui78vux/TvC3dnSJT/PraqDCy0BI9iriowPUtHSXe7W
pq/OiQuXeUIN+/Fy5jbkKy2waTIAZkqry6XzrARVeizD2x2PPCl1Gm0LhqbxA9Zw
Zdu1LJJFozGUH+rkbWIn5wca+g0R4NCfVhnjqyy5haVoN8+BtFI5sRQnAPYdOkNj
1TGgEv/VZVWzVgVKu2UQb3wu3/3S/LzJTu1mTkWTptHhFqacSxcow0knayn+vTRu
GBzjzejY//X8yBhKDhrsCn1B0tzBBkUTONOPStZzdZQQxMxgPn7ZaB7YNcFNxX1e
4rI4dimAVlWCvAxIgsaL0FRC8mvadGjwV9v2+Ie/TNMeA0afhxutZfMSxwOYH7NI
7okHP2380M9sqv5cnPQBDhBoqR43fWDEWKVnFa+swNDDE34oSRBl9fyqV1bFb85l
ktNoJAHILbbZGTJ8JEENW4fAWZkW9V8LevExIIqR8AG75EkYE9ht8HwX1Al9u00i
+tbcqNcOnbe5JnLr31fqw3WzqeAiVpCIcGKDKyzk59sS4vejLkkppOcKq/eGkX77
isbSGx0seMwGTZ1lF1r44xuasOgGulcVN9lt5ZLrulH7mQXl+YJ2PqgSZ8e9UY4g
j/B/FrYgsaTPtmjSsRVUZflSUmXufmeEGa2uCkH0CPOSR2ymQRFmDoJz80Yxkk5H
Q/ZCfL2t13DEJE8FakinN5XTfTlcGIxdLhnu++6iR90KoJkZ8+Fox02mEzFbIvuV
o88QvBcayZM63GsQYS9mMvdeLZz3TMR7ghZ7o3FP5BVfjki+y0OvOKN0Qz31ZHj4
Zysa1iuQdY2qSBSVIh8Z8c/DstbK4NJuyVxkqWfVfSAxfxRIa9NKj1kXzulvDanS
Ah/Ub+H46zX9qpMJfin1dQYt41YJOZ5M7rEyOH6XRodkDRIOwvgmX1E/XfZ9Xp/Q
cFLefJjyXYYuLureeNo67CJ9g6BV+ojsxAi9MM7GCl+hd+Wp/A8wdm5WpQmMmYGA
kPh7rKydOiwNytTSX5ezJkfoBNrLsnLojXrV1x7y6MvBbtpg+o8QoHwdALVTPt4q
Gu4QwkGmHg9HnUAQnKYdUwBnTRpZk7b0mhdiBQloI+V+PYa4ftbqKdfaLm5TXP27
cy6B9gXygqMRFuBzAr+lT36DknN0eW6mywp58I/lCpHInz3ZBQfLIjDbk/++rK8m
+FTbp4DqpgD1uOspoPmMeCf75fKfEe70soHmPTIFZ1GYG9mw2M55hewnIWPHVMeQ
M2fkEvhVlvE1X1sQwcnfk5d/OnY/o3YhVlJRA5ol2XHReIK0JXQbITzboIsdMMHC
sLBQE15Th2VZdGJKmL4I/RMe3yigJxxY/WNyaYz+ZeOE4Ap8rwkRck/cR87deX4y
CCUVAfWkiCJiYDMKkdZyfabVkCq2WaDOtqs5H18Bkh7yUPs17P3zonAJovGY09iS
0Q5dgGD82LLG4iZM5zSj11UBPtal+aLqR0hOupsAI0KfscizWN13AQpXhzoYhiZp
tAxD5X3TQtpZXkHnWvr2IKd5YEaGbkLZjIgRt1/KrgowNscC+zL5oObFbAZ1RdIN
MTJsoysNDuvzudn3SkDk+mV8ADIg6VXljyLZuLZx9aVMxUI+5hm/zcsUSXPa82yB
nba6rxFM8srHmdup89g5a9Ovnt1uT2SzhjssXcwErzXsWUq4Sk6He8tP+QWYg/39
+h0BtSz9Wyzyv2sGm4XL7uU9/uagCah5tTSEhmJgCF+EcTR4eXtgFIXYor+x983W
S6pg/vOtcim7o72CVa14L0pcMgBS7ciZPVVXI0bha7cBP3bE2TaMh5Uc6c/MoVFJ
XLEip2xhD9aImLD217iBGy8kJe6nZKNV6hZvo+z0xf+37VfgS0jvnvckR/xo1V9R
woUAEa81+Z3V6VwhPEA6VPBV4mycIujhuWKFhGlPJ9XJrscyZj6UFilzI2DzjDsa
x7udbx0quVm0a4R5iw4/xUjLyEa6rZzoQ7Sbp2jMWsvFeLmBzbrA1fGxoRrLIJJ7
wqFo2At36rPjwyaQn1bNA3nRsj2odXySySgBnDsu9av6sPcxbeWx1cggpIKIV138
AxUBuxzFZphXRPkJNsqHy/9eBnUw6olG6v/1bje0V5/J3SePHDJkIddEHvoDwafz
oKFB50N8yDQVOvEzarRok6Hv1xxkty461sao156bpt+OI1cQAm79kZGOIeLq9XbW
yM22NBtYMGJaBZ7Wkd7kJGeHq7kDpZvU93m4QXQdI8j015IDs0q0Qe+a6Y4Pf2vb
UqKVagTMqcofmcj88VI0+Vb7uvNMzr9cEF9rIEB2wBmw7xZMXfjJfan9yembFIzp
6HbVJWV4n9nAc64KcoZjYcxkHhy8f44Q0QlsdWJHTlHqAMWXUuFYMYzc4OZy6Ytx
sTSr79sPUvjweuC+9iQlqMbl1rkjrUjGOa4p+ZAa51kdo49g69G4Tv9UbbyFAhcQ
U1s3+V2RnxnFuoho2LY0VvTUVJ0SXQDhQ3FND3IbIF7lPuzN7Y+t0dXR68vsrVfY
8I1NFZ2X+ZLALjmRiPWl+Uv+mbZnUetYbURcqGfnH75/CF2HUhD/20CLZdhrq+fk
LGS9ZgBWe0DRW4XGsiiAAdWAoxbX+KSlX/Ka7tJo4GJ5sB0WZdWPXFeQ0QE+RRku
epdOWyY6Nag06UHdD1Hyuzlh1Bbh2kxb3SrUOczVISLx4K1iZH77DWNjlf4iFFhV
y+cAuValPs4lFhT/BDO81vUn1cwjFBEOdMXFM1prseS64BBiIR2pBnwy9uCQ9H1J
YqJbjlV/NZuWlYQ+1ehcxlojiM5YtRlpW/MRMcCVKqX/Lip94ZAp0Gs80IXJ0HY7
nhw1CF+8GbPGgeD53PdR+n/reoM70Tc+733BI2XDVqEho7bn6/A0o0v/whFcng3i
6C3X0Bx6WxkFteZKdFuEKF6TVSZ1uX8ktxvuDw+qnqw7xZDw3ue9saZVdsOjzFsm
PIJX4DjV/LwvfYuBz15sjZ/+Mb9zMWIHq+rBcvgICAAlua9lAvEq65bPw3GNP/9A
+Y7bKZcwcwKnNi+ZzYnmu/9GiQlv8GMba+vfOCqMcLDqmj5wIGSD1kYgXL6hoexD
qqfdU5m8NMlJTCr5IAy6ZIVWA2/oFbqJH25P4UR3+kk5koUSZ1tS7paRRFIM8yII
0NEoO53OH667d2kt50QTqjGoIdASyz/uYOJmVXeuCw7KtgvokmGvr4y3ZNsK/O1s
YLMIepehCQpWrqVgTpXrVOJ+zdrg3ey4u9pGdz9aJ4feHjIE4MQ2RP+HedE0e5e8
aSbVt/143WP8Dpkm8akompG6jOOykmZ+/Qije1optWDvStMXKc2tlYCWfBkYYAeo
pmFNXyHLlb4IL/d935KHJkRV3W5D1AwywMwsMThc5wnzzBoZgHfC6jMdd6DfbgWL
Rpy84sgX+/ASb3Kbkne20u8JV31aEHBVEVojagCbHsGIe8Dbf+xTX6NY5hxmHzKE
fvK5e2ukLQafF5WH4vic2ObWQTU1PW+Iz9exR/dwL1gBkGN86VcUHzFaxS6pULRs
gRNAi9JKtP1MyiGN9sQbx1hPh/7BjQj82Rypyw4rUfedQ6hDEWWEo2naL0AKJLQj
OLTFp9sf9b2pUIGPWoRxt155Ry1FSWeiQXPFuWHm+12A/4HLCdSrZEEK58mHdGqd
fmqU9c60e517dSksNYUQLueylgUO4ly3gqFNZIt7R1DG5l2hSJEgR/9RVH/xKRHm
POij64HS5P/WP0Y/OXNI0csSNevFzB2zuFTquHa8ad2r6GWugsZ0h3Z4rRswIRPE
rs4Gdr5aSo/k35zkle1Dj5nDrvuxNAb/PvT5hDXB43tUwxb+AGQ554Mw8zaULyn3
dxpL8jeHTIlrvILstvVRVnVOWPmSdhuyvpS1kmBJqmLxkxZJsWRFAGnwn8TjRIAL
I14ZOa/iBWAAFe+y/8xVWsRLJQcUZjjD46XXM8F2ey9cF1b2qnpbt2ExyMmHpMef
Wy8cGYO5uIPIP2Qt7UGARhaMgnu3pQgrURaTy0UA5pR1bXBfLsCA+ADPe9tz8yW5
l6LPmo9/D2cG/Yc2YcNXpLK7ze/eA6LzyUIBvivPh+D5FrmqQlL98RGZJirDwrAr
N6rADnsUSXwt4onT5gyahids3M5rUCyMwpQJ/Ol/pnKEc+chfjXwLlnj8np36NhG
ogDRERCam5GZ5TEurNg5SUtqPhgyyAcBUY1iNxJWRBP1xwytt8iiglhVOlcalsDY
zjwXuBhw5geejj8YFobcBIQorWipkbWZG85fmPqO85tAep3hHIxONl8/2oHX1G6Q
NKnjwWZFBFyq6H0UUH4q1pbNPYpD/LTaSFuEwa8XQaG7Biz9Jy2iqXIIVPbAGmCE
hK2Jqj3ZmifrdECvR2c8mBB9AYK8rDngocmZ1j38gRFirEjNgtzTZQnFabRA3YZK
vIzO0ngANmDCL6KnvxmdoLZHgASxvdnqG5sp5NDW0WZ8Ef1+NV6A600VHbttZeSb
ba8OhmOA1U7bX3gBgdQNDn3ZiCvTEcVXeWkXig5iOw3yeMBrK9TDE62Ouj3w2B2v
QTFj0LXvHBnO9GA6Zz411Qg+UxRBCorllw5eHlRHXAd153IaWhU2583f4WwAgvbM
PCZdNz2/4cPFn2aJK0Px3Gg9TS44IbLG4BjX64lEbEXWqPkiQbAJEoBfzUuAqNtG
i9cy5qXRmy07NH6//1t+OsrGXim0ZIFQUaIBb227U69zap1r1cfnj/WR8wVR+v8q
dkpnENXN8TkNI+7L79AGUqG4aiqGgrGNe4qQ5NlxATWnk62q7ktEHhJ9w7ZQemYz
OUawMx7ZhmVMXOnw/MH50MhRoGFOl7aewwNHGI58zFU7yyS1enm25W6TY6teNUWs
1pkfwnlYNWyTGuRjqlk4ei7K2wceIXo0gFFCpeqE3byDlsQFZVmU2aPKw7fm+UsD
1J6XoWcUxvSdJvPv3YkxgnQrAGLwgRq87Ym/T8N8UY7+iCbY/R4Gb9prEgi6jgwS
OX/+yLQJ/z+oSsfJdpUVChGvhToed7hhR7ViVkR1JY3hMfhMez1Zct9QEqoDLG3Q
K1EnIlr+P5HdrfrmShi0uTcQzG3xR+mskZvC9C1QXPP1leVPeC/nkhB73e05o4Lc
q2xKx0k+qhdm26sCAfeVisDz3aO5so+b4oKJBghDT2XCw3lzW4Wb7Xu6eU5ewWOC
IUirBgSWmTFW8FF4J3gAajfAMOPStK6bnVYTs4W6IC6bnxi3tZRdKzVxSlMGW+26
fHXQDr8jdBVlGl8bbgcNumcCT8ZEePPQhnSjNDx/mS45bJkEQCkAdG+FM2Jn80SH
rVqKNCI/0fSDd8KtZR9vw+E6omT516m4iAQLr93VT8/1JccdrUxltkp2runjr5bo
ijPAY+W5wM4mjhf0Vz2JjELmsPCI3/lrwmG2yDSQODMadUbxYD8Le8dxaDLxDbxR
LXn7DgkcKnPSvY5KX1QgDddMD8gSXHNpy33JM+eynbw2XCj/9ar8Xp6kWar2m0KG
g2e3pdW/BXOtPicVNoxd2vzPMGz7hMyK6PqBIObP4EEZZWg5Ixy8ZGxFepDqaxGV
VT1OSjIdJ+T5eCEzu22wwMm56zzX/kp7Z65eMen0gWwba1m6jrmduXRIulnYFYQs
YFUpvztFDIDKZQrExV1VbPiP+C4HHvVlYaLZScnmjmpIkNCms/Pkzpq0g0fhx3Yd
DznAxl4kOrfNxqJ7FhjZiFgt/oLxJsfHXDc0nTFAtC4ovya72tH22eKnjL6ubGzr
WXNCi622t6I0gQr4QhshlN6NVWrMAydDpol0UMBYIE0Sw+mI0K8ZY54M1dmvlYrR
rvqHbGtECscYtd3wHrNbw+MULMYyqIG4xbpgt0BBcbzgZIYIeb7Kv4FNxafMO0QX
TIZgnk3Gc+rUddC5gZ2EcMNd+2BVcd7L8iiXQAt9nEGBryJEx8IraDL147/9FOxI
8TEjYA/QkrzimIBGcukvZP22Ijbyvlh3dEnXclNorKUgOEt5KC7kZC5gAMRJnnW/
2ri+/roDdBWUahp3nKBgSXL12LhBVFNiXtrdB5UceFj7mQj6FwO3QMHH8nSNhyw9
K2Rg4h8FLHMdVt5Iz60ABDVWtGwsiGuJoOJIGAC8//qTGDYRUhhhP9GYz4JiOWjA
T2x+HQocnQaI5k+Aoe5lHPyGaGySpSmrE5L4Dg4OIgZJ8Gnz56maIGwsOTaANP1P
fHH0Bo9/OpCRoFOrdKSlqyfj58gxnq3S838QMc8gSnN1Ol/r8GjjjFjEO41W8pfM
Hsej8E8jTY/OMLYS3rpR0meSeUtXP+PmoQ9EnOJRd+b6vsFhJj4lFr6cVT3spxm7
tLAh/7B/l1wI9MscaDFw7afpNy1ltLeRwfmSOanqsz+sJhI0Zar4df3rRSIy96dV
GTIBJAde94FIemAi6v3POpLf+BwWUJr8q1Ora8P4mbeUidynY6ajvW523K3jtklu
/J0VQs4Dwp78vLx0A0q3Ocg7Klk+4KRA7tgTHFPdMFt7kLbUW7YOV3ce3QioNnMR
eKytW6jkG1YMGp0fcz+btoHU3cJMfmaLGRIk9ph44ChoZVU6BSZ/1Rn+mU3ObyQx
A/zeYgoTViJKaZzH30S1rRZUgRLS+Q6m0TCD+Uj4NpGsmwr0MD4695zUXiqhBfi/
Krc/kjuobm6l5LLyKGNvuezpaK4oOiz8H/SAai0Fz/ETjcyz0rQFPdd1GqaSYcDW
k3cIBfwLHEaVDmH6pRXiDWkxryDYeNHY90Oaqqg/SqpdJdveA8O0vhEPzEQ9zpJB
kfwOS7D2AA7v3DBSaL2oi49Ms40kuRpBVsijznCGDQMWAjOHsITUQSGYk0ossPIP
EXRCbNCKm+AXs1HnAwhR2UywncfqyfpeRj8tW+Q8wAomKGFZCpnrpKF9eu36n2eP
D0Tw1aDWrwYv/DJo6iiGpM6N2Xo6VrTry7LRfrx6ADe/WVMc60vdbCbwT7YbkWUf
hF1xkUYqG6rU4J9fo4yfhcBH/4BTY/d5TTp08mjfqOYLKdAkI8NeNY5hGLxSND+0
FYv2SSDtqOJKFRiqMX8agIv6C91mnVoFRzpvOqDwHk0Mr6RMQxOTzGYVkZUgMelS
+SKlkP9sZsVjXpU3TGXOJ/SjbhKKgLwgWVeYX2puqBWFTLZIQbig+V/yE5fVXDx1
Q+vMgdyu/bAJ172qM2X6vWMHs8o/7cJGOeXa5UwUk715LBS0fiieOcpBPMkYaeZN
t3K/dXP1wpRjw4N1MaqPL3CIkzrckYNtfJ0RDGS9oDU4xhxFNTRxqiJRF84pHbY4
AF6J487eUjviP2pS0th+SIFzlstCOekUCk0w8bop/wd7IQSqfaOkbc9+Kq+pLmvr
uXkOiptLp8Ob5SbkRxvwGcZXKfQutnn1ch7sYCEyWMOsYZhSizNzY3QKRcN8MLMW
lbbJyMIWovmixR4wUdJ4fEuZ2bKmMulUROKa+7fIcuD8jYRhoyHOwqv4ngt7MzPR
JfeMQtyABRntt614fx7OEmtD0TA106+vxmU+SnHocBfCwif33+pLY03R6iaZGG+P
Uy7ftxnSigbawQrtEOQEsoYCTNftzCTC9Ob4KMIsf3ZIHj7z4nmibmTdi9x4oRbf
LCKWkX+fboYqeNEYeJJFskXWFc24yFQ26EOFa23db/LZjrJzU3BSZdxMn6z70+Il
oXcSnUN9ASYKzvABO0635Vv8TnRXx2CrdJR2pvlBj8V0OPIWYg2IvJNAq+WVJfjk
LHJX5VkxutjTESVPQk8KGzU0bClpsIiu+dGPPhfnbGMMw9ELVlcFPdUJJNFWzHLG
Uf6LEuhegpBMLu0fwP+oe+q16AgxMJKf3CzwBHTvkF1M0cLJvE9hQuzpyXAHrHw2
4xtBGuRQfh+xUrPEgkvwfGC8tTCLtQj9npd+5JVqFW3PJNWjnDHXbBk3hnoYNL0R
WYKP5FaIahZmuniuKN6gtPN/lufv2ULecC/W7I5HPt06o4y9+p8ILZU+C1GLvZvq
ETSRM227wqQ8euEIuvomt8xsUV7HEYHc0d/LsXfpicaA4jqxNNFOadisDU9FV7ud
oJAO2KhIeB4sPFtBb51ma4smaZRk/wAXutAWnB7C3inBZcbrx36iFytrNdqMIZ1M
zGE9tSF7ByzCc4iUTCxo27NPP8Zp/1MR3dlSplKn+W/docIW1lP1LW0gCMNZQNPN
JgIFefRG+/3Rc1OuepVojguBNJ+VChUMR8qYGhdWh8PBKe9/jPZvmQ/G1zuOJaNb
8OX27aVfothhUy06av9hVgGlSvz7ofFi4ohtZNHa3BaQBvOwZuZVxfUkMAJD2CJ8
evSP2R5yEdVcmV2UamzFxkmWVHw+yLdUKJ2mEiVrxU9Imps0ccfs5rXOUSlkrH9s
MBx7CxKG2QSvoobt8n/BFgQqaRst+kxnWo7t+RLNGJgP21Tj8XeClB6q4jMV2MzW
bcIy3guQyNjDKVsZX2KocX4ALBmK/KMZnUQs/vDJTVr8F1/AzjDRo7QyvbJZWj0t
xwgn6GkgcOqrgcZMxg+JfjJEGmX24X2Rq0l1Fvu2l0Iy7Bz3fj6nexGEz2SvBmas
A4/54T6BQMZ+wE6MZPvOP9Ccevq4B/YO2fDorIxvtBL892PSe8CCF9iSuheoyDpz
AV2n59xWs+DOpa1CtkNdk/uK5oW0a4lMqbhbmg6cXUnkcEu7AdfluYe1vtxblx9y
OS/KHGiGSddFPZuxBgEGIuCXPH5nKC2qA8epc3dOvRxtTfDgSx1qxIH+BvZ/Qaum
2Q/cIwjWPqUwehHBfCaZhEB3DuGmEANDPToB6QweACehLEjsnrZZKvQCEM71Ow5S
YdWhBWpyhyMr64PEH6jXmbiJG7xX1KZr2d56hqvdetQG6o4kMOKby5K5LpEe+V4X
cq9fD9ApMtWe3VNofWjpDCKkNQwCgQ/jXcyBIeFOJa3Q7krRYgOa3jOti1sTNuaN
NLptXePebUSJbDNCv3M6YeSvAvr78SDfQDtytbMvwNJzGxC5UN1XhlEeUwAdDZSG
HmLnFWNK6KD8DdtucmQpZhp/Cox9NbFTnJeKf8J+8w+EsYcEJ0UBqTs+FcAdzjiM
oaQPqXe2USQepAbzfF5SuZHVfRIflFZka2DLF5zP6iQ52ZMe3vYHOstD0GY5KIa/
rdmU/olNOHcDV+0AbXS9PdLJIruBxMCzkV4rx2z9FfOqawZiH0zDQ8jl+tABCLtT
L00QAikG2uSP5ZtxEvZJbo20yXoFcCSKF1TA1X0igfYVskqX1M9+Wi+BS5r3atAo
C+ePAROKzcrz4sQ04DgYkIWy/PBDOQ0FYjOrQN1Lz/+SyBkdkZeIbrPzo+FTzYTt
s3m4xTpAq7DFD8re99AdriIs/wGfkKx+XcMfUz+SoYZh6TOe0WVpoJoL7NPr0e91
jSZG9+gGX5Crdtcsd4mXj0m2t6tL0RKz4aHYJUWVeNbBVxklv/RyKIkjc3KfIMy+
4LgNrDVpJ1yY5/E9/TB4czyi6aTsEWn4FyWlkU0Y+XxlZfVZAiX+I7DbJlwCBY26
7S4kSJz+O531lO6Ayr86g1EzrthKQZ2Co2wzIApSBOEIlgWhXsxyRWfxVW9H7LnQ
BBrOdnQY1l47D3VB9GDmxA+fxlJaGr/7dTj9XBDPeGr8QxPzg2UfvPkGy0KzL/M0
7A8s8ptQufdHPESETeE3mfr9F2eguiQCvvVZ19M5rpqRn6MCndEv5Rg1n/wyzptt
hgcEj8hEN8wcE68FLv/UKFOZBG/qwrr69bZf9YY7OS2+rlkVakDv7/0YqSshzgIY
NL+Aft2oxG0OBB+jNz+BSBY4O1X+ffngaUi65HwzyyUtzyqvkfq/fjbgnzLrw13o
njOcyEECIgpSlnLFFifPpAEiUDFw0OhGhMs5WbRQ2H0FY6cL5vyriBmS9sX5XJE1
1qqOP+ZErUVy+uKwVeZrHNWEQTRzA+xh4v71S0xmqbWb9SYUO/YUPM30btNIPUtm
qtlw5wPe2IthXvXiLmA8pB1qvGxsEu4gHLW3B47DoQlhIyhQhd36XROkA13SKVUL
v7j6FNOkUHc6r+0f3uhcWg2VWFTUJWbNlqXNmU3wubK4qGPxmmFbaG929lS0fGMU
mHoGrLXZmsl5/ZYwW/3qs20zDDdWouBvQOIQcyXlmQC8eFTNT3FN0KvAyOCHwPZ1
9Hm3sWsRPa/ie7sPHqZ8bfa8kGb+OsCh3PlkkHzEr21MLtG9vBVW1Fz5fV8lsovt
V8Re6s+OMpr6V2qTTpGRU7dGEse4AlBdv/NJKNJE0hRDYX6Ck2lOu9KW+ihe5WiL
Ai6wgnq74zaH9h2+1j+Dz4YMZgb53Bu574AqIRqYGzMgdL70htlkPGEDHfm0pHwS
pNszuFuK3DepmGVmWcF6FMbtkGg78S/fjNr+dZsyWIe2FwhhBFffvLBwjfhjw8v7
n26fa0me/mE+IDrI3gh9s2pIvjLQVXQwnJFVzh0968giXGmy4ukDHVH/DZJciJbu
uU1meSFjTsbS2Ua2ClKxZ2+a54PvWjrJQ2i1pSW5/ZtHCRt8J4sHmI6e2/rzLOhN
1u3vISGMZ/616F19dWkeQtYST6mj8DST2t8W98w45K02nnUhZ2LqTNmbnZyOmyb2
ULqM9sFBfJqM4gvC31DtOYjRqlBs/wb4wmX90v5oTRuouFdbVHDuvI4vtDltxsRr
JNoju6QPwLRvi2oClQ9DTqhnTtw9kkzNI+703xnLxfmyBuHh2umFA+HO62SM9NKh
QN9qK0gvpQEEJ0VTp2zJT7iPmUEfNJltbivziJ6+ruq6xVCOtzstKp9To+uw3TUp
FnziTxhio/GTz5DEwjPZKLAAPn46LouuKug1DUF808mL7C/FY7H5XzjP0aKQKbDg
oa9pfZb/7GcDXiX2nXYNTagFb3oWmJBVuqkbYIeP2uGORCMBKosf6NX/IytLDaDC
lAOvKvMb4tWhLSwMWyCLTS5OKExfojVTFtqq1s4quTZTDHc1UQWjzxYpr1qE9ZI3
7CC3Rk/vdJqmpsCC86KGUfiCsSV6nzH+zYZrj6EKVPmK9dy6Ix+7hOxVYzLnlTqD
ulV2nG0OuUV3QboNNSppDFoiNrp03q7qLfYFQQ42EZvWXpHBTURaM4WzC38vBGAl
JhpRx0nMWU5dmsGfW6H3mZgaXQ3v1V2X2rwlVWbslPnIx+aQY4PzYJA/maumHest
zrEHlL789wPPN10wkUQVshb8UioqLEYQ6xkF+DTdJMBn2QEXr1onPlMzPtQC19F3
DdDIvdyZOqACF6cQsUyjKtqh/gVHpgwUt/X+WwFBG+VCYxOI112WpV17IVl2n0Uf
B+F3jN7p6LNFBUqNTvSMe6ZpRiPDpFe/4F3Zq303W+jbSnSXKFZDMbsev+kLXtt+
E/2SZjAPXsfR/q0Jg7KG1hxykYME5EyJEMM/O6QG9RawX5/jYowDQW7908tPBOhH
gcwIS1qtWGWqS4uPK3fk4RhX6n2M44ztzfoke+GczDwB6hjtmhK4DjfeUaLjTeLP
UHiMdQ8cn6sOneV3YFycux6D6J0q1bSsBBDTgy0XZ4YFT35bao2+Rq/XZDOvWgmz
6mXckA8DUTE6757FWZoZ2j5Kasjh4pHbC+x4+5OIZ8DedSzEu/jXcl4of2udDvRl
d7AljVZORUtCrlon8PQ6XqwzIq5239mMF9LgTLcBQpUex1EnpsgwNSj1a1jS+gzj
G+k1LuIg0Jwfb3gYZ4jVqGD3Hqyt5DNAaXM1A1AFgjNUfYgbjTy9u7v+jvV90VPn
5/RHQ9C6KTQoWeL2f52WhSW7JOrgcqXlaaWeFLc88EgCJzPHV9RmeDDvyAY+MGUX
B8PLxxdMLu/Yz+7H2uvsUomlHCrvUd7P+d0R4K7r8Dz9T50uMSYCOro83PvubySs
aO4HwlYOcCMAmtiXURbDXiKrG1s0WbMReD13CwhmeypAujQ7rMW/0son5yPUMV2Y
aqiZfDYDDjlKkr79UMfvtI1PBelXlUktnghLRMulNZkdzeh2eJw1g0ovAp+Z9zGp
DOnE3JGn/S/GiR/tOxddVCBRinL8SfDtYOIxdveBmSWQCvhdTRQU+rsc/nceImfP
yWb6DpaNwRqaodschYQu4Z23MTKN6JX61Ct4DU1eiBRIwwqYzceOjXRY9HlCieSo
NrbcWfwgIIGyOxSuL4Vdm35Fozy3iqZzD5DxkwlpVNE6t3vZsMvctq3447fg+hIR
7aXFKcDlyKtmZsGF+su+H3nCg1tM0fTTG5svqIucREHoPyfQ+RfAE9FYa/I2CAtJ
E9JbabFoYb/AF9HECkzakb/7l+G6FNvEqCPpJmJW04Yo1YSfP3J9OyWImveQ9Wui
NwM9WNl3Tr4iIAafyJtU+45cdO1G5fCnbuVoZiXKq5zeIW7uEWjRIhkE5NYMMg28
f+zxNZi+vMv4ClPVpc/OqMroNuTA+b812KElOpePyV4rQ/qe52uPJ/O2vQRD7L84
J2u5JKQFGFtHtUviXSASg9Ace93CYd1fb9qTj+l0gVyrAsnd3J1s4oEyrKVrCYKC
evJscPe0i6IKeUPD47DnhpvvZrLsWlaqVgT1+1pu60dCnRVhgWHfY84/auqy5O7g
s+41HnT5CxjoFLLUmE4Nqdu600r9qxttlqGclXobatPWdTmSc2PntKLxyw3CFDGw
i9y5Hb5KOTYIud1k09b/fZnYQEmXcz46j/sFNeBSJwnaI9kmIF7m2c1awtOmai58
ZVyI5pylEsgmPnd/S4CzobEjyZ4CTemf3cd9jEw1GShOOEHgdWJ50H9XyQ3O2bvo
t0jmkyyrnDsJqLyDH6e/g/9WALu8Xl+vIPBcwu+4T8PKbE5S3LzsECZ2oKwXghV7
akNk2awN49/EIAWmcTWz7V03tHl9mxvMtkaHidY3p+mOnJQt6msml8It6JSnPi1S
0LQ5L5FMwSZ9/ksiKZUV18Dpm5f6PZiUogwX1kdU+U07qt6sVBzY6JbiOACFuyrt
TNisvpNosdOC85yDKUSQU6bZV+Uw6PHU8novROw54ePgV0FreoBjCUK9L8Ug2Mjq
ghtZtE457psQ303RsAyp+15L6dTJw7WkfjncrtQNEgtXgGPnTJUTc7/sLT7FcYmC
UPkisV1lqnhqzt4a2zb7g6hKT7sqvdcvGVfmgbwwf3yF76H2AF9JjLce5JJAin2n
3ro9+JiNAqMZHjtOVoFPr45TvBuSyNjzctTp75KkXfGmiSF4dAl2aaFclSNpc1y6
uxhrHyu1ztxjD4ShFFNHDRDoUUY+AwefGD5JF2huNlIfCfnhIdfduv5/wB+k+Xty
DaEe4Z85AwRGGQduRNK79D9oEUCe2E5gTBrelxD7HUVfN4VP+RscpYuI2sniBrx3
Mq6ZEhpbd1N96NzidGexx4J8tZyn80QanCtxQ6hVGE5jBc2wM1AbzsQXTrER+BA0
pkn70waeMCZlEzzPHILATsqiKomA5xz/tZYr5EdREqMqM7d537beTRQy+wWqSvzm
zueGBg9m2I6TrjXk6bcoI6AuyxDpGBKcWf0JhB2e7+J7eG53maP21HeGvjlYl+R1
yrFvcVHzljioRhUWFA0N5BaJbsLob5D+kFFLFqD/zA0sA5UDYYpM3cthHnEg7VuG
uqwfmU4Hj/UGCsJa1e/DiP5oouUz5X9fvvztfV/f13wDOwwrFMDhM3KPrUDbYTuq
MIyCE87/XPMwmd1RWRbk1R44aRrvUM9yASl2NMOSshY0LZaiufEuSIV/sY+rwX2P
SeNS6RZeBifVn24sLL3o/5MirSl8WAntGjQvUNGER4IKdcjvgS2Q7kbuemy6Jek/
DNj1Y9oF5Tap0FRgM4huNZFaltliJaPodXwHN+lnRnD4MDiNiah70wp6fjPSm0y4
ZBY3RdxwoFL3Nwnf/dDxMcT8NbNYJJ1cfa/zj+wA8VXGM+E/tjZLone/6DJIV6D/
kWFyeEepMTbTC9G5vJEd+nATmIav6pJ0eOOzQAli8vPwdtKh9kt0/miKsF1drdhb
1ZOxMNn0dQrLpo6khe+IKRVHaLQMsvQZvIMq8AI40nLUSsko2Qt3wQD6DBQs3bzP
oeO/hezfgZy4uT4opG1fv1v5C+cbFjpmJh54AjQ17dj+iq0jTg84N96y3UBZub8Q
PdZZiDjriInFbcfhjp8PoBDi/cCE98jkvuKW2l35nahxwU9lq3mSCRMn9LbDeiQi
BKkXqs+FgpQhtSbORi8NSz2VGdUISHiULo65IMQSy78sqLgaUonCU6iWEB+rdRbH
XqAT5roy5AfGzPQUei0AaOgYzCz4SmSTj2cf3X31GmUPEiVMycbHzkuL2ha2SUcd
HV8TFxL7x7dn1NRY6HVO92lPAykkzrKiEYObjP83QvoQ1gLEtdBTLvhmPNhmHZXk
3g6vGwHT9fwdTeMVG7Kx/t+OSjqNz5GVMe0iW60gdWaMBC1DXBMpc11lJMfl+s8N
yxnbIzZ0W172vDv2Egh7oonK/sBQYBPuUusd7jWj/0SXGQllf5s3zD7QO3wYdxhQ
xqrsFXThFrcI/LGzLpeJgjIgeEcKh+amL3PZjRVRJDJMgi4VACw893kKc9yqscLy
2Kiz0iUA/Fhy6qnujVYuebAGubrp7mlZXTTzBz6N+LysbJMrzypiAjlo14DDNyda
Rot2/HfxhIGCmdwXTn+Q1DY1oQodplZj8Yv8t2JktJEO/OPX+yPz/kyEoESwf3Pa
kVWn66o5Vp90jUwJSjpCGTfv6MWqLrhih5AsKi213P/eGYHNnf8cUctChHMc9YeR
cIaPEFNIRj3KyAJHyKnF0OGXgO3sPjZrvKEBUMeyWqE52aTtrOm9DgSK8/zyJXXN
AjvvmxGrF5KzgqjgbhPU0TmN1Y/NLeG7bEpZ5h2QYlYgNlg1WV7LP2X5zPh7thkk
7dzFZS8iNPjNmGa+FhnikOqfelvLN38VtTm2INLTSItoIdmjHCBI036V54BIkZv1
IVU3SQ7lZrw/M90+qjqjKblYmvGEWeoub8R2R9M+5+iD2aEpFCYHsIcBIi1JNNG+
WgYYnue6ozsZFELmClp82VI1Rvn7orLFSMEZrNJOWOCWgbawBQw90s6WjIdaInMd
/IBXd4aVpSIixC8fcg1DvmM40J6AlX5PT+KZFeJDfkxG1/ZRrCKMdoshmuTybhvv
DkFzYUPy6g0+BGRqf2sKfGgwA3sDBkI+qVcS8PLAUW2JYNIWO4ZHSxlYpO9b/GLm
Wde0w+/XjA0ByCaxjXLcWczUwWR5AaXPp1mOM5RTzrPaloguqkME2XG1YsgpKIku
V5fM1OgCAFXL3uRoOtUHYEZMKbR+yJ2romPvg3ZJNACcaOCTcLokSsoN4acvjaAa
CbPsBmX1O3OJJVWsPuxdTytbL1pg9t/si3DGFqU3/ZlkrrPjvzOI5eAUrngNI86L
abZoqyc3tJ7dWA/a9SIPj1XLmfDl3ZzmcpbmPSToIDmy3ZylPl1J+vYqLv3jJh7/
wq3g8vSVS4wPLdOsjMQrWEoV9OkcF+S9vNFfFXgBSCA8odxzuH5CMKJyMixqIqi0
bgTRlkVzSA9AvIJueis4wOnDWPqzURkChUrU4JxD4vI8lxUq6I4OuY0Yh+RnjqRO
Xv21gdYr69zD9vuIjVfzaVzOBnNyZ7gTYdgpfzkkYXbfOPvNaKMO+zFVx6qpLMgt
4cthSmoC62uOwaqLUMluOYBmqgXWNLWYbGpGnbAtozc3mJqoH45TFL6JojjuOk+b
/3XX5Z9juh7JsGObC7X7SV7FO+muE0tnaICHO1NUSLFQoNtRsqvNZTloSiWLX7mt
8ueOnPg9egoP0OMOoCBl6TKUvk3SZRPSzNpMiGs2OhB6Ec6uR8HbKnrALTHsIaxA
O1PveiAI2VMpFl/26HYsKN+R3q4gks9LZE8IJlUMPSahxomOcEfUw6QJRP2NHYqo
/82bnfCbAGotTFBLUL65lHCFlBP3vwYBvjj2UnnE3XoGetB5N1yx6tKi2WpZMHdR
xFpHUespIMuzPlR03TcNAeNfn3d742FlS9nF7Zf8T8SMApgUkGmEsmysotk7/5Fo
Lq30FzB/+WdBCkX3qJ2wdxza0tvAX7ECB8uSi4DmduixHLRH1d4UQCuzym4AyC4Z
J7XgcSB5PF4hLdAqOBSZgk7aN3BjQ8BW2ktivHmlnVJKqiTj3yZu8/nzF3f/vJwA
TvqkmDcgbOr7Taw0A8itHFHkNKuSkslsNQC0qppqv0Jwt7O5ET3JXc1yKKx1DbWS
qSm/t3eI1Ro3XxxBTYidU+mzcBfoYvANTdIO9MVxTZ2u6oFU6weOvzonGpK1k/wp
KTGJF1M+tf5KsQfJehzRfy9Gaw2sWIoDx3GwZfzVuITupCnwoUB+hstO5xKVfP7j
KCH2u0bQm4oDYilmXVzujvq/UvKrkBUQyBRKcnRQ5bJoqeufRssdv2KeI9aFN07o
oAmkCupbt/1wzwQpFIxWqr8BMA6GIcOhZl9GdPU8hVohzQb8SX9pe9uH4JZ7LK75
1MsD63kQ1r4L/5CBOgjl45o3Am/tCXL1NvfUYyy4CZQ/ZlnxBgSw5wCwQNWLjcIJ
VbRoRnxgIdUntbC6bvqvpRkjuCwLaggIh8WcdbB/j5wHkIG6smiWmsbOcEkKKCxp
bWBdcZp28HGRCEDRKzzxe8ld0KYDTeBaJB0WZUldpLXYTv5M+iF4DvAXeHnzDfvZ
fGoAqEARMylUJdZaObuYZtlL9QT8furUaY6EasO+X09FNBTgm2nS5K2d8kB6Y5ge
ZCwavx9rLeU6e7QKW1hxa139PJXFCBjDx1Y8wKP4GWrvUkgi6lpIklX+Lrf1ZVwh
Csay8qkKkc8YRQt5ROtoz26wYxYxNwc9VvY8uGdbrHeYB1Y39ume++AHiPcICyE1
vDBbFnPRa8KIrH9jUNZKtN9uPmtrcAlGlTB4OneDOHhMgOYLjkaPK0SpeBP+MG1i
sWx0YECEC/cz1mTlxG/IV70ifjRWTMF04jCSqnBnVFY7awgM2td/9mJPxyEsp9dP
vY2DjemeTBEp6O8RL/QnfZJWITU6GsGBif1Z5k3OePDTn6qQNuw5jVFzhoI82kmO
coEVuS5wjox9qM207FPNi0TijMn9NKMvP7qCvR4zrWiqLMJVS7/isdqsORHOY3tZ
iyPD7owoTPMIjvK4CoAocAC+MG0CsE2zwmEi4kElHBqVKprn2ZxtsDSJXa381lFT
LBLWxp9wteHsRiI/z/H5efNnxyfu+JSpZKlxtextz1/0xYlZChF2SBnLNfhkwxrj
1Y/kfm0/xL3h8Ot0Abc1QGXoW4PeSFnsTSQewFHG2HKK6hOiZRuW6QZ2OOfGUI8T
PZdxtPpv9p6XbKFHS0jOUFj27EgCp7f0o7dFhS2Cv8YaFi1x3o4ESMt6GCn0Bz1/
p0EQ3uDHySZcOHnsIk+PT1K3f2l79WAswltVYIT8LTnK1uSS/GZexpWjssDCHYyP
ncxlLXsJvG5YyhNhjRLYf7wbpntol1TmUxaFJAX52QRwL5d5tTqIkN2IJ0vknDV3
5CaTBfhvbfY/DCDwmO+9dkgpZDtwzvhKeFu9hopkTG/of8ryDfGdor6rvXjd6y/O
zec837w1/YV4HyMWhPNYmERnH2GHO8iDkz0Egbw2aT/TpEI9dBdyADeut8f/hn5o
b0TI3RR9OR7+qOLIY9biSBw8c3pJgSa6hNaimUDps2l2YbMcUme8TCZ4qYqGOO71
JHN4O73HbRZHpqRMyaBLycMqmNzJFuK92piTEG1FYyRJERvkq69HNGtMslMuCemZ
Rs9KtXJ/0wZVBXsepMvI+cMTNcffhfZWJWWpNlWeSs8M7HlTamGCPKSHP51nRV/D
lgPPSjGJNm1e2zmvNUQObIfTFroo/cdWcPpHqFSTgzcnkCLgErI05GkiwCMnaix9
5Rx1n+m5rCtO38Zo/VaIeKacJ1Oan5AvAvN68vJjCknsVlJEe5WIyt3yq7rJcV6f
wCSerCVEYtMI2e/B4rxOxge2AqHTQRhbVX10VsAaS9gdcfl6hFRNlcJPBGVvhhwM
YTize5ygByMD/TUqGyD6aH+NoGZ6fpYteZa2kmHz/uE9vmu7dL63UpSr6qZVxcua
Gadw+B4Q2/mI2KQg+LXEfBWtULjxBPzAiJDjIHEKv/LG+cHrMBmlUH7gTR515Rtd
zIGsr2WAAJe4jdM9qnVX8H7SDGRVktWVZZCrQI7zT6Cl6V+9bK6Hjjo2ISkICsaY
b+zJSeMHYpdpPHZLdYlxnXpPzHwP17Vf7GtBK5NI8cFJbMdWvPekHUGQPpQH8sSa
l+5L0ngcjeMuvRmLLzoYPmWe+MXpW/XiG7IGulpv8jJVSGe88wmRT5FPHZ/DYG/Z
mO7UhH9CMII/bqbx+tFrZxXKHNmB4bIv1ZaBLwgH/r6wyW9z7DIlbr5nAcv+i0/k
EMCQ8NHeopcvqYgN2PMZq5h8HWfINt3rhT2oTA5X10AQ1Ugo1dft8QfLQBOWPoTt
WL7vfOajkkcdRypjRVyeyUFrH0zpDPqdcW7Q/5w1iqaVJKoxQQZqTza1k1/c0j2B
cSS3X56DCukK3uwZ9tBt6XuLm1xe4dArGkK4mYtQ9MyNIux1OuDkwuXDhE9PXQ25
byJvXHOihTkioONudEhoKITpCD3C6OvV4Lz5n9PLmxJd65Slrs/Ffa5XG2Rx2c61
juVkFe5Gcxc3Z67ZWLp7WMU9DXoGftF77iwr9090JbGHBsevFcz+WHQ5sIQXcG4n
Oj9vsIedVRLSbTOaptN/6WB8mBxyHf/XF4U0hPDBCkJ3nKKYJjSztFms93CDQDpF
EB3fg/Xc25zbqHi/x1XKNKiAsjVHftuOjW7YS1cxWkWdphwdH+MRauZLU0VZ0tJv
6l6HJvCnwTgBWDPt1EYUle54iQCTqBfwpuLZ5e0ImG+OUyisGzbkUxpmTahSI8aT
2KI3XHiLz4hp+4hRoPtqEBderrC82YJcbvUKe8KIwdLtfQ/V2Ko7ZrypSV6RI3P7
NBU4yG4ThjkeANU4el2NvDlGACfLWdi2J1u5qA6hmNcv01N4asb93xlmHnKWErsX
SxQ/h3NgU7amojZmANtToW5mC7g7eEEqJXkVrxRytakdScp1N6KCrflOUUQOmIT/
A70KmNJn2KZXZNE3IPFuo/RoEdJDt61NB0F4wN5bjZnxMgqAvLGuD8cIIlMnyK//
ktkQVHUjSviZh2ePvq98PuWiqsVHcBbc8t5B3gI+wUYTkJvRgM+r0VodCMMIoxnw
r7Xw+SsXV/SskvaB0VMyFU9LTGV9dejraK+3yhQneSK9B1wNMBlNXPNtRMLnjgM1
n/B7gD1pEZfDSxAtrgARvWkItAijh9Y+XBJeWZr7WYcZV8TVbkb9Vk089TloN/57
29QNb8aGBe77+ufXDRyEE7VbgCl7iHfmvJsu19KtWUnrwQ8HAOn3+xzd0EJsmMAH
yWkPhyqOHkrtEzO4h91CL0vUu5IsaLPMes6AyJejUO+Zbke+4dl76UqwffzL+wL6
lobFYi5ssNVPpi5Nzw6tvjNicu03SyJCnkusVfyh17/rExCKfbsk+lwtt12huApw
y5Mt0CPb6AGopvg2WB5gw5roVUDE526Ptu5VnEUnDzkkISCXwaPNjNAw6dYv7fjA
aRGN0v2q2MM+XyncQjtMi8CcVCUskIrE+9YrBwoRZClwLawPKFhUnUf6AMa4MFB2
nduKDf4g6gE9FnBrUXTPYhQcuM0OqikIHhAMSeSi0JT7ZBv/BgkV8p9j4Ke0JJ0A
9E39sKXIknXHEOy3YpqA8rCVyT09vneFX1uE8eu0iT1nBcJCFHeC6jHdhhpLz4Df
8kl4llUruOTqGOvr6pJo9IlZzyRW6D0eP5bZXenmvP7nKzDchp7SdlhcH6w71Y0c
JQIgeYZ5HthjqP0CfwnT6uq58blxBJnWTkwlOJ9R3hYWdFQL3g0je3CDnA7ON66C
lNhpXNUhPI+RJHtjozntOSVCZjK2uzVXcQxlvq2R5RCKVjB7AQ2vpoxGcNIFnVpt
YGwQBMQGSXjbPG35HkMF2uDWGyVJqd9b/BkuiN7k6E4+qW81PRPVlf4NL0oaMFow
jceyPbOpX8BTR737nZzoEP52Xu/meYJrt3BbjGZfMKoY3Zo8+bMQ+KW404FfFNz7
VPVyR3P1smelQk/vcvnhhsqpmga8GRtYRQ7wZzm/hIIgP4dAqoDplMuMWqj+wJKc
h3/P3LIZn/EiOTr8j+XIOnbBzBVnw3Va0BTYuWEpl2UhzmFMUQX3IAHuXkVa/2Sy
zr2DKA/0Vy3tou0WD5tfPcomm3pxG0U3m+x+Tw8tcH6uSkWNciygXPDUdIyvlC30
jh7idKuTvgyDBfGxqBfcFf4ORmctdPLERevTtqcVMY+XW4tCInMHv/yBJ9MqQgKE
jqPQHUzRXs4RXyUld7mKfrZW8prijjoxlQ0IMp5EmveAU4VsCrChegZEetVgDTtY
L9Cd+qzjFadQ98F7fWwxo4F5NfRWS/PFxtsKWhajKJWhP8K167zOuGgx5tYIVEbt
Bwqfu/ArAnCcOobvJgYO2HOi7NbiZwco2TMuNJD5tdIX3u1W8wLkADjdnvI/uiUR
3W5jKUQ1DbBqDXHhcBEE+Q3gyeDiRHAB8rIfpx+oKZjbbNAvgfHRsIt6YZuWjthw
FB0ZqX0TBIjNEXZA2UWVdOJjCeA4NrS/MXTfhAsSMqP1Eew0hnfdgQ+OXi3jTomq
/PAzJypuKNezmulIY+uNW5xqgh2OunzzpbTQyBBRYLEiY7OEEvz1gO82pJoJqZmL
/VmVNRvM6HZacpMsDdXlW7SmWvtLAQDzPEaUYPBKReTXCFz+BWXIAbbZ0Ew5vJ/c
JNOQXf2np6NLFVPMgzkpqzjzcXO9IZHihWLyXQzi/RlA8YxsDC6EYuD06LV8VXJn
FYuiav2YJy9NfcuXDS7NAdEqAqBdIBYgJgP4MpByPPMc3hM1cnZ/1Z3TsCl2D6Ms
dF9OJAr2KNPHhsrr4Y5vrCLb1JxxON2sMtCHPmFpJQD8vIC7TjyMUfvAfUGCX+bt
CO+qTxbbMjQYnlk5QmT3VTExXhPZAMmegRpMzeTGLs9+ZRBsBIZbCPUhOiBRQLsI
Upqgm6l5iBeyLrM8yh7CZ7OZetiIjhG4j/8fe1E7EusRgYqfQp3nzkUHnXAnr7n7
cEQc0NQE0o+e+rAdNys7firotpwetg4fBNW0vghxRnHVYEYhk+JORZD3lNlifdi1
k5ePK0VjUWfZtQn38gYLcy7NuYwWkd0GVGgO3Mt8US7jMHPTfaSGUn1ie5GCRW+E
AjKLSdfFCpvDj0OMrX+XeExEkzRfnCv85VIaz/rUVuobYVaHdCk2Ou6LVWPl6Buh
vwCyrDDoI3sU49Epxyl7wvUWUKhUwWYx5t2ALUmUPnpnZt1XM/ruktVmwthR3PdM
yWJLN/O6cO2APxf79BldyfuOLG6E5mfzZPE+MHUGwQupNH2nZzHKk1qZxFEYqZko
SJecf1EpACRrCsyxquJDFXx88X/VQ/3g2tcUGEqetRpETjVXUsiLFgXJF5YsidEc
KGMGvu/ZjzVWWiFbfyLDqczEcGa2CD+sXc5pi07ghiohIE9RtHnEYtNyVU7Hr74E
pQ5TGzByHIMMV38XI7NAEbQjxZuW7YMv5MwFgorLUnLdr7XJTv7YdM9gTzHGdqll
wBtyX8nUZFjYasbrKrFsxBi3SOC5PYmhuO7vWgHHp4Wb0bhOolWgbYnOk/Wno467
GbWR0zmjz9tiXl0AAiAOMSOMnPoDL2uj7Y5keSCMCoqKmMvhi8z5veSf/7eb82q6
ohFmk8RePUzHU266ahmdfebGbFqa6B/haVrfiOI3J+TMdIvjI8XPx68J4Jke+ThH
gPBxT4V4fb59BViXRdeNIb6fcPc5/EO654chxTWFMwCtaW5ALLAFOBdTaIDUEic9
YxcKAgYaQJ7xIoB3cWRvMeLTkiLaeMCwG9NHqzayue3erwyTNyZBCwm0/wwXOa6v
Z7VAjYlCbJjByI6pVerJSaEW7ICKNCt9eXdQkJvDyaqLXVC3snmUXMCizknZhefy
yLs5ziJlvTcjBwIun1hhc/VouPyvmhv5Pkg0u5iUCn+AFwCVJYHCpVvu0dIvbJgT
s3w5PA5O72RnBl0ju1re1hOjozL+RzCgkApsxs/PES6UFni1XE59JhTVEonVMnnH
6Jn5C+bkAPlktBKImCZbpisRVqwoAF1BBWcxuX+6ZTvQmhn/DR/KxnF+QiFC1hXn
p25rLQFOKuNlTHxl9hnng1b4zjPJRllICcthNzyOUAlD2Oemjmj+7SlPhGaaYml0
+Jxy14lvDLv1t8fIfLIVlwBJppxuS311cgguhZm+qV9k5j4XobloSRxOehOTPaM2
+wes/oe8ryu45I0P7XY7i2iJwSvJ/g3f8KI7zSIgiFA3/0JRMMkyMlS2uvslqtnn
xS/rgLNVLVS958+4O2olYvfvdE3Cul7vd2chCYE+LSZ1pxQRQmNHSqjEALPqztGt
Fu+pPLi5EI6PuQJtknxBoYdgwA9VyleQWi46lAuyHXfNTa1ljoPSHDbK5x1FP+jp
yEFsV0cY00hrmTfUBKksDIitsNeZROa7NtiIb444YpPHTKNgcnj+UacwbnVlY5xX
GbpXg+z3LtF/WrC92vAESwsjiUAHM8NBcpYBQeJLmh4q3ViXyI4dS+M4aLtGGZZk
ZC/pYrjtcKB5LJQ80/GDLKmYoezpCb6TqliqqL38duZ1ShzCl/4ky1Vbq3V1ADFq
dgNAk8QrAURM3vg2RK8gH0v43SFsAdojF41SGiU4xhl/25ca+JlXTI9FUvWcNskO
0CE6usyZaFewmkwgKG+176OYZY1DPyKiEg1vy7MLxL9+Apf7L4n819N9K5DWYI7z
80IEBhoHsptfw8wX8/xkQ4ItxkJrN0tyIgfhs+ukUczuHb+5gJj3p16YC5dN9b1J
+174NLfA5iAnOv4Hs057lADBdbb8Ttj+2Li1+UCbwGUnr9JI/+qnWX4oxc02nXo/
Z1sMW2RFsDuazGAUtEoMM8CKtdHv3hQA6i235+hFujI2K1JIzNZSTz95RuKKFIhd
lIV4dfpskvl+galpRQ/yLMq2MTpZpdAtgQEJk+5GivjrPAzixY2s/puE/+jvYpAQ
H1KN2UTbIEUoaKmGEPyKpSVLYCxXpGNb3KA6Pb43CZKk/QLKsox9iykymPKe+nDh
mLhkynyzQMeDSyn3wbiKtQpkeR0vccHnp9AiVUthJ9TNy2y+adwu6Y+RoVVJTkLp
FyRzOAFNAc1MB/aFkppLfzvy1WH2JEJZsrdiqfTeXoc5f7yTsGq1FPD+TCqbDL5E
Sur7tdd9kpqpdOD8/AU/0V1FP4WamiJMeacJloz0+R/p7sTCMKNpmofnnx3bfmLO
KgJYawAQG1NVqT6ROdhYJqb6Rhvn72lDThYS0GtvJZbGj8KbVC9lNrk5YcWwdblb
iW2FYYMWY3sfOE8FU7PH3KahC5rfhmhcXmZeP1Bf1VLjwZOXeMtTC7yHbVtWMhfB
T7IQnRyukkWoxUvfiT53oKJfu5Zp/ssUC9FxkRdYSUufr8GH4LqTThXDPaJXFEtK
QcC4ySigZncEmrByMS14X7prAMSmrj7ZxTSzgodpmrLdtlkK67otY4KGP2jUX1Li
caxSjB96wviAznXBGfxmgNqnqz9cp4m8STbNmKCSNi1xIiPNZVpc4LpDA5f6UQmn
hix23V8CcumSB2nPiX4eQUlCRDprL6iXHLCM3IkQbPXFs+aKerKCKcVlKXuwlBd/
eUA2b+wNvjf4j55NBHipSRKRLfCjJUNwO5EeT6Sep6SHZuj8ABdOdXueNCOiyb3b
AljK00M3yleLDlcgXMV3RiBihuSqEHV557DPsEV0pyKYKLZJXZCuzX3voGnLcqnT
iuzvcHtnLAzRCPhoMliqbVEyqrGP+bXWD5Lc6vbusk3+nDMAR+h36dfATn8085oj
vuquLSYhLUo/kyZrbNnD6HZH9UfBKd4fzcsOrYFdqhBF1gS3m5e9gWAsmUp8+dg4
XiiCb9erLPsdKhgw0xVYWKJwzp7rpJI2M08SwSfXojFRYApnXKoY24SL26+qcsGA
6bggmm7ND6eE2hKzQ9RAXbgUidqEZ3hislw8S2CWtU47jU9BUTp6PIxy4DESySDn
yE6tWjh67Yj5eiQETyn0kIA8EWTggLVUJYqJccTxlp/arayFNFBV3EwzIZU71gJa
Zs+Jevsk5zkVZpxKpcu411iX7rVVrHOwaORLS/Hny6qvYEougH2T/60Y2dq35WdU
ib55JqPXc5FwKYoo0PDEgrAgdWp5Ms2VI8oS1FT7YNyzpXymW+I2xZko4Oytyhgj
1b49kidUlDy4VsV4An8+2VgEBO8nnsuF0fVyjbP1x0sYMworBIf2JLb2ixvHe4dN
7ntDxq8RkTaqOf367DL2jvRR44WYrf7xAIS0IY9MxfaE150YdaoM667Ak+zzK9cp
SQY53+v2xmw4n96izBUV418ZDk1Rcp6cgpC6rrpSPaKl3QiKZaW3s2hVRAFNsHiO
D6JsgdmtHiCqk6U217/eJeSlWTRy/fo+rN0K+7U+csu+751I7s4cSajsC9Bky363
erylCm8uT0L/Wxs2iUBT/sH+zmarKoRQ4UYwAbm/KcoPij5Bsu281axFIlta19SC
oOGI6Zw1aXlDTHqRkajlxvKceQZtyF9vWVygyFlypCzgvv3kDUwaQ5HAoJ0+vQHU
pFG1WXvabLBiAwtZNl2Hy4c7Rhh3g1cZOmGm8JvPXkVRk74W0Zo8V75Q1FLvwKoQ
Q7N9Y8YVYkNKhhH61ijV4os4ExfELT4ju2nWYRhLgbOZ4glk/GOG1B6Ll/ruSLLz
EnvRl8X5a669LZYiJrMBnHgS/kYJIunPVTwDAYGvG5fiuPTAJ5mhVihC6LRc3v8t
nVhEZ5qHh9D8M/7xBgNYrKXNGC8qyoFKlfHjlNs/JbJWaJi7l3X69fHeH6/S1vHy
mT66Bq9ruFTL/+Ad09KuRMwEDvxehduiQdwKhgeEZUsxi87RsBNEnWkHBdZGg8Zr
xxxlLwBr9MArMXB3X4drJ5qErkqSKMuTr+epJRA0GtyiFceCkZndr2JKkpfucf/Y
Bl3q8qipCsovDUGrtcdI8rbP2YOrYbNFfz7cIaVqk5C8PMF+qOrROLxZKA8FJbwk
+QJgIHxK9L4oW/pNVtOFYxwqVmIe5rZnA9h/P7/6pEd7N02bYsCzMGpe2vlL6buo
vspDaCIH3jawCLEJttAAnI+5Y/Ql63dh3oeBe4uxwUOZyTA+OIFcvzO6L1YJMyxS
2WU3MjQ2Sg88/yvBjUDb2YKkP29PGMnOrz6dyjOAqTPceraihIcZuoBRzP8XmZBL
Tic1VEpbQ2U2ehUPV+vgQY7a54gBU2UE30ng4gaYVg8J3VRYM0xyyjHjP0r/dbC9
NtZNJiNfbgZPUZDieJDR94sPRScr7uOl85w2FvqAi4vwHl/DSfPvXxBPmvxlMXOG
gxgP3Wb5w+iES0hkx37t4ujfq+jKTh7OToD/oQSoemiJCIWfZy/k1o+4YfRZhWXA
FEv76ihOG/OeVNWZ9QRXUrntulmoeEsQlxAK6EFvAqWvuB0BytKsDFp1AEP2khG/
Q7XlTKjfhUu3z1gd15lMyDheA2ugNtbhJeLNJR3g8ERwJ/DLOcs61QqT0GNQbRWv
xc7KQ+XMQHOw5FCLOXffdBkTmbnqYy6wmmSEOT5E4NNvbpF92Yjqg5bEL/6RgcOw
SVyN+E4aRuPMJnK12yWwbMsCjwS999tFmJiKSSEsK6rQRIUiuhi0/PboZPsKf3Bt
rNPrUMBQADmRWE08E4Fbeq6ZQQ25XsrU6up/A7PBEIRaF7CtT4ldW2CCcuDrURUu
5TeeDcgk+EVOXZoJNzwhCUhM5Ch22Bc0Z6yr/umXRkb0ssNDb5UKqfDlhDuX0UUQ
4DRNYHK4JYEm2qcOElUPDt/1xN4t1O5u07pbtydcOyIBVO6+vtgqigi1jVXBv5ZX
+Pj7jRGDt3h+LiSeF3NJ1KE+c2TN+Wa/ae94R7owlYqx3U9IZ+FY0agd6ey5yodR
p86GE0vqw/uGvG5C0QLdg6IX0hM6VJVyUIJ+YzLm5wylL6bqxii9EOPlJV2Z/V1U
7zvR+t1xOOpm/D8c5fGvFPHgO8cb//WkoZ8s5mF6DVFps8fTGuCEbzQhhiThbKJQ
rrg0qOTJQxc+nZlv44SFPOB7dxpeL8ab1iWp0KSewFO3QpcdUn6EOPPjgd9V8hhS
O3verc5Aa0wT5hfKIRg/DbbTSv4lDWg1fCiM5/Ot0BtzlqFmZmkGzZ/F3o/Yf53/
aiFrfrLMuXntntYOOXuvE/EBes8BDfTSwGKKTfNSSc34NMWMYh7RnSWlo4ERmZrf
i7yV0htF2qlnH36BscGWIpPtiCh4RwP9f7/xWsoQDQvFzw5BjgdtWq7uXlgWhHNS
l8yRqyBbzT9ZoxoYM1unRryvydSFZTNuGJFa1+X+RSnkzDt+0DEOXJv/frSo0XeF
Orp4AoqZ9PZNvhwMJrwZHp9SocatEReb2V8wv8zIsC9emduVKgxAfVIT8vova8BC
+3aCnJnHOrZq0hoYmqdo3rXcZG8izNpkuiqxDoD0og1my0gM6qK3+IMQ5j9awXoL
T9clb8Yf9Ita5bkQxzs65iuCX7Eudz9vR+k3pGjPeY/Jv9TWsk5ZMIoCllG8kDuF
kHYfkcmBpacxgIMFznvTnWNbUeVRU+youzqHAmY0kgH6oogmQCxMQpwW31P37w9r
2MuATNB1XNttzxz7LjYvQWGrkHXqFqMxsctOVOBn9Hi8FdqyzRB7Unqp69+cIcLi
KE+jOhGKXgEIbjGXGt2ugzAeDpNU0916fbWn6hbaZ+h8KBqCPcgWPj5wjiiM94Ve
RZdWutAgd3tmU/drHXRjHAOOHxFAZR6PV7WVS16V2S4Hjg6358d700G5S1nCO3k6
pvan+QUlNIO96j7WK1g2Djt5wGYcXb82t4u1NH1KiZCFZyFlCjUMstLelZUpaTr8
JMggj3eV4PKCcLIhlfyidqBxv0Ctv2G98jGups0fN8ganWUZ+a/3/4/UYBbXL0jx
SvDkFWXtaaYoTibD+ZqL6AWsWyTlIzFcXHhk8AMBFyWH80CVrrOaBfZY3EhQOLAo
UFvzsQcY/Y579BOgqnLeco9wtRUN8P7WG43+/mZ8PrY5o4tQ1pqRMNskiJHPwmBQ
KZgQOPLTqfs+rcsGSL89vkMGYRStsSxPZAfPoFsFDOVWnN9MPmRWyvdRRft2kMDo
dYUwMXTuBFgApG2hsbSJRaOBTL5IIvu8dwRxJqa83/SwrGE5ov+uKmvk6bsSjZl7
TT30tPlESGHlJ/VPObEPv7J6lnByFGC4y8eYCaqx6EcRSfauIYFhUrqhQU2ZnIDn
CqsuHRyVCuBfUBiKBmOHwXLId83ziv2YBs1K5WbA/5RhIhZfjDsG79puVJh+1oHM
D1/TEmep9wwD8d5oOuOCzY+t4A9xkCXAGQDgJLozyUXUVjRlXKnecDQZu9+k1Xw9
pIZEHqd+AkpT6hq4kKDrSrHSO0h3ESPd4vV0ytUH/G9Pu6M0tL0jac4H4gCbtkbI
3pzrBsT0hwWHjzdebHsdfn6wGNs1D2rHSlbuVmDJi+7HkUuK4ufryO6uV/M/IMEu
2pMOa5q+Y5q8y1E6G0MG9aG6Z318iMRGoxlXRM9RrPBv9Adt4YH5ZRWMT2QYT7fV
KOBUGkYw67htERuACYZQoYCcK/20GVSzF8bESPsIMQudm94J9HA1kQbsy2pLWm8h
kSZRh0oVt0ZUv/wdUWUy050nWA0musMszhd0iN9JEx8Fx30eenKe7hTYUHrCYMjY
VC3fLAuTlT4nZ+EYyr4m5r+ewXp9Rpjp7pEwaBV8J05d1JLRoFaF87UQNfSJ6Wnz
Xn9xdrL79/nPeDdZAMfUkTne8UHBaZQyj6TgX/o817+0qeoJf/wwEzRY8GS2bOJb
jWwK3j74dJtonimNMFTzITLAuvjMk2qZSoaUqbqOu83nZoHTb8wnuSmONRzpZYLA
A093P6073/fEkBudryKKPtbgJGzHhw/lDMLaYHiFH8YFPvvT+t1GLtZYVMdbtszb
/UooPKCRgp3q+OJnFlrgOP1pYp5TLBLCa0XvFPC2QfulILJW+nN5hG/IDn0+aRH/
TvTkBa8zhysQaZyaBpcL6BfS7NduH+cKVcYbvT14/zqYVSE/RmyhnMFlwK62psvG
ITy3D+vvH8V/0kggLBNV1jjOVJQi4pckOC1D95lXG7nt1P+51I4TcC2dtaZtjCQB
680vpsKuWEiy7/jOjP5JbB/HxC/inpZ7Vefy0Ik7PA5IQ3j238eOS0SEGJGkNBuM
pe0WaT0hE3N0Yjd/gFaFv1q50ii665VikTvfAs+Nutx4Q1G3lYhugIH4xL7n/zys
Lm10cdVXfUqhACSv/ulXB+cKf4eQdqP78B6I+sLpXM7mjos/YhbjaNypB5G80QxD
l+ii+EITqdRr0emLwN3trneVwWqgsc51v0jWih0hzW1WTfidhKYx7FqnK9XnO6LD
NICZrF+DsP+Gm8z2VzWVt6g9jEaihdZmDTFAncvR20JvUYVqUQGSWEserlWBvC+c
jgYfz3PZxijiPlAI0QphlubV02HYL6q3jsOHg9dUpSlsu+iWHlbzBZ1lCFNluNwn
CLcPKLnTj47gN8kg0a8y5ykBdgli+5Hsb273bBW5+hn6li846Px2Rx6AAtH1GT7H
r28jsfCDR6mJ2qjaLXESckD7voAzWlj2AiS27+vGaHDnA0GQ97DKHYOFoYhbgZu8
KHviWI0n0QPk91blf8Au+SBXQ2QiAFf068UUuwmOVDbxTCJE4ZdtJn5nlAtb9rYG
tHPwBds2Mji08MTKVCTOrR8QGW2qGnbeXnLV2kb3ysMMUdegmria9NNOqTldORzU
+eqk8MAdMrQU80U8NQUQCn/wX3Ei0DNfTQGvM7FzopkBtRt2Da6AmyE0s2tXA6Co
7MinK3sPjFgB21N+o7p/6I2ZW+ZqwkffryiODggcBSPBd3HCGZ9jxq0K5xRqqPd7
rpCn0bmdfDvNjwNhoohgS5suU2iQksZ6ZoV/x9B7mqyNm8ke0RqfWuGqDbC0qvGi
cQ6RmnxIZOJPJFw0l+ZqufTC31MFcKtNO4JAMDmzX/WcF802ZS8NF2Zev/VunxgJ
jPTilSKioQr0V1wj3f+3+gBhJBKCPnBZ0h171JykuFaY62hEem0p6ZIRhc5jg7B9
rGH7kk68XWbzItd0/aEdjw0xVnibUL1el/MSls3LsYjhZyWhB0FARvDvYhxfMMVu
9I6L7BzpKgzawWQIePqVwihi0wKrTHWVtFktAL+Jo236mI7G+FOV8rJU49KVxk3j
sA8z6E9IbkogtR4SltLaDaI0pPC5HmW+TQ8Vcsfo+6CUC+QNUzcQfDqs4+Is3DwV
urxqUjqrjySDqU5P3DpODXbbZoVxE/dIkB0bv6mAb89JZt6aRB2YcqVvUslF6qDQ
VMVS9A80tdjl6hA0b/MM1vSrtsElgWd3Dw2qgOqen+b5WJlxumyl5NYrdbNk+lav
chjaKBj29cLL/VmtB7QG7B91e3vKmaEDpj6ixpoBP7UVjBB06rvHeMzjIH8ovd5a
/WyOhuuqXrcvF5trUv8XUZarS4HYvipWZdSm5oebmBOC6Uyf5TOHc0UteiciP43I
Rx2tZteXT4zHT0UoMxJ4mNVOqnJAFuPALlLLRKiDcRWTLLKCpu3nxP9rrCzaDioU
lqVibIlVU2b7SFq9WW1Rc8z8zqknON0gcEACcgBtQfgCiY6qRChrc5n01v/jYxfp
bUnSgzDch4RQOinoJBzBTivIBlHf+hc78pCLHAUXUs3WYIDzoDQQV5f2kCohJj/i
lBDFWPgNHv1QPS1XjDK8hJ7rmhfGPv+6MnWajZ+CjDJbb9gHX5VxURIGkcOEzKtn
UTDEDAWF7Ft3b8xa8kBQqK4lTKL/3s7F+oejnmcOvXUWX+h15d/luW99yr152/zM
zg4bt5PETIG+GJpMW0b8WzINXdZf4X16LPxTcafvier/fb1UpPIoavi87IzHp54M
jMHxYLiVfxpmEvVNFygnE04ZlGq3DgYTTNfR/OGjTE9LTRdMWpSxC2WtJmDxb8/Z
TpScNhnkdYOA/CYiKxzQBBdzbnO/K5hrCl4qKTQbXHKc19GHeaaVGF+AU4BhXiRN
tgs5qHQ9tjA63pBB6ZLPBnMBmu0wBtPHfWqQNdGibr1tWxEoRyWyzHljiKJQygJh
h2Y0O4jGQyAxUnuuEHNGGyBHPzli1TZ+/81ZzbdbUklEKKTLjtCqlFzRomjczM/i
J+OEIIuDLItSwECKvwfmNS4RzUzaqPveEE3f7kc3OIzdqTYUpRtwhdS3Xqb4aipX
sP8KsRUDsLpPtUNBppC0tL0iJfzP0MYaLFCyPnzrmUQaCIWl8hTuuC8aUuOa2E2O
mmR5KH73jKMibgh+nAm9Ih3g0mmBNAgO/BKVd71vQsKTumQNJIxMCVBISK9Jgl2T
yxlfVZ8fio8ENsvBImxILlnCYf9URIUEyXY5wHeA2Xn7UlpIwVaFj5ofQAndwXZA
fxAy2TnyJcThmxjRNHkyngJeycCwcM7U2PX8JPXeEFY+FBh2oDOqVTM28cIHoioI
wIB2kP5+C1GicenhV8cSgmUg/CA1SpmjJeSmktY/F0v7GX3MbSF8BoBpeMxkQHKI
EgSdG7ttyMgnJ+hPbtsQ9jB2eUa3HrTUDla0CnF3dTyfRGwcpEMwCaZJ4fhHMMEY
xiBp+aQ2Gvboa3gE5ecFSJ7FuRI2rzdU19TndoVqrawc2Etm5JN0g65JqanQ2bUC
7Ssy2QIrnkVZz/VJrE7j0oBQMdEjgZygdyUFIfBynVqERfNxBbgZljR0nNS6UNV3
S/BKtMxVgF7p+Jm8ENOEdB6c4aLdy+qNf+RJMrjYUDpHxTuPQ59kHzObx3b0BxYM
3T3ix/vShuWlSRagjZt1/JyWZ71RxoJARDUvrwuM4IqYAoia6Li7qKaSsRIM4KPs
EOj/E4xxFDugUZYdEoYhT9BP7pd0s9POoVI7ZQ1iLxi7A+Hjq2mo3in3lVzDOZ3i
HW/RAr0zWE3I+KG5S7gSTcKcSCZUa0uLgeT+K7o0D2Rm27VZ5ob+CtHUHofVMWnS
W5vNd2kDcSLGdPNPfHPgdXATeFyqpgUEsgU06mavirTV8zIKdmufseN+EZ5QpBES
zj3bw6Xd9C7g9dbJ5Mk92ucfuplibAYN/BOllJLRf4ymZE7r4549XRx2f7Mjq7pd
P53vYkHundW94xZ7KJxnZO5/DQJ/rDi4HyXmbmP6PNpOiQYmjhhxscuezxti1pXx
S78yzmtdgZ5Q50tcsszENBmOTrbEpLDM0Uc7r0bpWCUMSjZX45fUTODe/6X3ctSw
HsDyiJGJlhvj6bmmxExuMuImNU+2tD7SfEovu2TbmU0aqgBvOGp7QJUBn7GLmIu3
aZwKl1RbUvE8MWyW/RckBxvyyiBViul9cy8XleebyDAyr+kfQizfs37W/1GLASih
24ob6XuSaBqMy70EkdEhUSvpSHARWSETks9Z2qC3q/2v0dxNbKqU/ZId16eeOniq
mDIYR3jCoVQB4Qse7N/w7x2TCAoMVCODEFBVc0d4KHE/VfSZl6Mv8dR1jk1RNQgG
ORqVyt8poa7WQ0N7CxtB6hl+Y5T4KqcyFIlMYmiWAjHEVmA9iUU8iFbwM9gCfYWo
W4M47DlsuvtePmZjTIMHOzUD2iaVjPcMI2yj6b707diH5IOpitjSAgw9PiqSgWzJ
PilfzPLA7BBlZjOVLV47u+dYPYHw/AhD+gBEZCDIXHFDsD5YOTxvG050RqKYFX1W
q2pAn17bVcVWzDETV5ZzKa54ZnbO1BgmqJ3R/WYTJ9+hs6QkaF+Fgw8b2JdDYKCw
DN2eXKguQkkZy802WIYerMLa/Iz0c436tyDGupWXe2Ei7qsy3gmCkcyhxYlDBD2D
WsVtnVC6yCeEX1efSJqAd5dpyZ+Lb8EHG0kV4DiHvy4/hd/K0g25ihEHPHIJwDDu
ghQc0ZfLiFZZXMrkaNxlXtcYT3wc6l249z2xz/joTjVlczmQZ3MOcbEQorfBHVBT
pOK1nCIaoUFt4z45Gp5eY3e1Tna+opvAjIcw+aeiHwl6FqImF1X6gpuQ1FSAsfe9
ofjd5iiU6LfWCVzDgqNPGMHoTZgQhPRJC9BqCNoCbKHK37Oyyqqg/gnF2JDlOeBy
rvTmspMcjkqaT1zlMt0kW1//i0raDv4cl6wKTVaiAgaLxMCYP7VgA9tjI09z/Iv9
A9HBMZ6ItOA5vFfhuC+/vof3Hf4fz8M6dkyJS2hDVdo7TJMplcJxJRV+2pzInhBp
VizXGUXmly+hIWVSKfG6lOL2X//D4vuGgpvT2JSomkqJSFHGHtWxr4uA3nAYJHPl
8kEreXBYyldQ/AbcuR2rV8DFCFjJCsgWgmDjGXCTKBLUPclJSZuFB6K1jDvAxOLF
abHzVaMyzKc2xo1CSzc3i+82qE+cIvjzICe9UayIPoxFAlWZOhzk9MriFMW11O0F
S5jsTc/PCakuGlYNju3uqP7os5Cxnz7ykXuTRIT4Nc1AeNs2Rfjtg0eeekEZLIk6
U3hXU5b2h7QwTjHceMrHfh6ghRoHFZ5teDGS4lLLX+Nv6+tf3EX5DVTW3tBBCPqV
W9WQC8lBu+Vf/Cwp9fNdbJ7yOx0ibYpgABzPdnMMfPBLbhRdVF4x8K2+JKEOl3UT
5QocstANy/k4hgMJ6L98oW2uXkb8bc8VTfWQT+iItf6+oabnC83mSgk5rVx/WNKN
O/RVwh594BkDMx8pF45AWsFayf1mB4Km9KLmSiJL4Zix6V374b6fOeGVBXxqKMtH
5bByKBDlDvve0UQZEBlgq4HoUO+qy7M+0dwjYhl/VUxb55W2r0YnTJR+j6vga4wN
hZBcPmKBcooCUQgVqawh6jRybmSRdke/2USNk/91mKoHpRu2L9Awg7VStE+iHB7b
peHyOnRxjBICBW9cWRZ543bCJqQmWriL66g9LiccZQjq1TUYPh/iBD7WBOWtL2Vi
lwMEmfY0Nxf5rZ5h84aZLVYS9mEDpF1iSJMZ2xVfSuyEfM2Ed+Oyeki/PrcWGi2a
Ux6P9oavNDyagUJWABWynSASD/IDpntfaZcha22RWSEq03nHNA2Xa9LDx2BMO3tu
deh5aGLNYQJ4i38kMMgVfrzAGyHhGEELbJfoJ+BUUWFH/4lI8CKV8qwcGQ8jgAiy
nZf5YX+gfLh43shiLEak4YLWhCHHCvYv5uaIYl3If3bCUCQNJ1+zMmCt3nPSCSzO
32ym/a1Ox1J4AvAzODn40Ku2M4oY4HI1wEFIIZJcgpaenz6XqNvTl+LkOOu8Dmr/
KD3LLFJ1cbcYPB7c5oiIICSh5a8xsa2CtlvG4C8tpc7PyxC32QimiPBfJdQh1cqm
2VQdWGEpEKLxuJgONbhwJmD32+2ftNpI4/FJpXN1pmcN5BpcZDbUhuRk6aN5pKUI
Epp+6WFsLHg/TSkyQ3h8B1v7jZfjf5IhWjaaHfT6WdjMvdjPPeyFAiWjBooHv6bg
GzZEfG4SEEHpIktWV0nEZxa9YsVUKfAzvtq00wM1hVqGxZ10UUTGCSHS2IWyFfVY
b7HUTVXkYHO/OCnwsNAdv46Z2wylH/s7sBvUz3d6UZ55o9RqenD78lI9FjLjmQOY
msQPRqm5abAQl4QQX6/y2fQcc0pAlIZRTqpbtz6Pe3XiidWGYUrctZqThI8+Xblg
rX7w8OFfNWdh+SObAxRvpftF6TJOzl4dmJLOPqNj9mw4ZzL4IuaEG1hWaaODcEdH
ylWmNtT9eoZUwlrNHsyii3M3paeUwIrVeFzC/cFTjevuV324UWmDFHIPrJvl/mVS
3Yr8XqXKJ+fMUihkP8gBvKwqkV8SrQgzKTdT4IqVTj1Z9PR8l4ELl41dmX9Ug8dd
52QxGgRRDD2JHzYmlN3gt+mB/FfOAC00cGDNGahHNr40KXjLhm8Gt5rYkrdAGlxj
QWGJ/FETWxF35O753cN9jMhqV32s0Rs0fPU3TE1y7SYDmCTpUNLQ4QaFBvU/BiuN
KJ/faLV1yo7qoXRyHxMKnQHx/cV5/ZIiHFSCFdCbkmTTwh7CR/JBrn8BYjp3catC
w25LbGWRYMDMgSvDKhi6J6lGRXzQaO6+awUmaKbPGXpu5N2MceTfC4rB5YaAqja1
vhedG9sTmbYoJzEXQ9Cfstc9NaZLekKgLTld2y0dLDbizqbnBSJQ4nxxVIW3zWMS
tMxbetOaPCxAUwRzc38pZt2lyenypyPdl+8Qx54a2BhopnM/ZCbQxyehpzVJTgU8
kCPT1SkUYsoSqp+B32JhFOYgDaxtUhFwprRJr52nUOXTZWf2Pl4+lwTY2Pc5nmLQ
AgbzD7lxpv13BZTJYvyNAXXBuFKIUZBFBCVTXfISmbBelFxVMS8LLl7QWMaVcyFV
iEZv9W3u1dR5ZYsY/cBObaZYa0rUabfuyapNVbeBGUay3O5UJWzTUTV2NX2uvfRw
TLW5JFTzk/w8j1Rx8jGPWsLligyi0TFxOORvHbdhAFMmWgCOAv5c+sYzHQngUIcq
HCfL8+oCOIVh63jnj7zf/rM0pLxxBUbOzYxON2vct8kLK3RjiYr5syC0vLmlAdy9
GN6cIXSYH7n1H067hSVtWgTmtzcEovRE1/W+M0Zg32rACBVqStQalfTmtAxqAHgH
LgZrAgvYUSTmhXU9As6T0GmFy8c8VB/KopvrXps9xwE2Fd7CzzPMz2QMjWlkfytT
HGl28ITSwwsQPNgKBrnvcGjZfdz6rbd2SqQwE5dk41+SNlD0L1yeWi3T8+jh8DLO
6YTxE419ENKD9w15ICQqlHtDl32Q2WDU5124E9SH3KQyvYxEEOCp9TukC1nlQGzj
ug8kNgpzEU1/xwT4SNIqQl0H7AWFNfG3skYkwYOYvmS6/4O2CI2RKjeXOPqCgw73
GfIzg2t797A8lpAztNI8tukbRc1iGbr9oPzHEPJ58a+lk3LkeIYSFGbdwWEPAiFE
rO+a61Dpv/3doP/fGnrMCnvgMUeE+nV3ScAKBLwk3B9A/6lDESqqUHr5Zv6qzH92
pyeCVW6ljhGn3m/Ahy7rxOFajNasxOxVE72zKwv+Pb0RyoTsd3k1ZpRhAIBaE8ID
97tKFHXoU1X54qfrhXv16q0PCFz4cngc/lmn/lo0ZbYIrWBKYWRs+wERhL4VJuxt
yetNRAz/i4sI+Z9r9/F1gJgxTz32M5h2rs95m0WgjlVrxaEHeLV9LYEwg/7L80J7
/Zphigod/I0pfc17uD5IqgaQROHEdONTS8D+J/F2/FpbOCfLwe7c7rXg7QsqAS/X
lAQoxjL8tFGBH7gK0VwfTSi3rJrD4pAvRuLtC4eJ+QQHCBE2A3oVvDKB5JdPOBOj
VDWc9n6iNJJdwraHwxN6WVEbRj975QidCd+Ab1Lw4KZ9qV9VoadvRuF7xKikURkY
U2n5Qd3qNX+CNJxn3BwfahK/d86HiLEUctxj2w/tlG01pAHhrgZEF8WHYSkNXXCS
uCdHKMTzdbxBFKp9svkTFDsAZCVz3xO9HLfR+cchWZ96PXnaAO3cYqhKx6+sUXlR
hTlAyOwQPHQftxoTEpr8XB9Zmyh8/HpC8SwTPUWFearHAyoogsxocRmHL1lpiXNy
yfUiYaoIi6oAl4dlwF0ZY4sESYQ4bOXQp77B17Au6xEINko0hVzSPgtJmxGggGrF
ss112uEBRKDstaKTxouU9Kh/T6aeyjNP734EHqiLorIzl/yJstIedbzXaltAdQSD
bbyb+8+trb9yeyaLAViXXzrRrv9qpSgpOottl86YIfABZNMzp5ZXNses+Pm64twU
X+p8jRVvbneBHmOR+xmJnUg5HvQRxkguE3vhPYKUbTRuNUhsbiZtTRMhItDRKdKA
TfE+FPD/9PDpNh0DGor7jSqybAOiM8SdupwqIwCiZxdLFDmpnbMZMPCPDV0wYqsb
nxl1G3kRYwQXHUznxahjJf+mhG8U3v3wcHsNF4riz/j7Ap1lRHu602x/arAzehQA
qsPOLx6/3bdCQ+9mhfFYSDtOREHzN0ZoYoy9LQoEGRIMGeQVPdoyvguHb0yiTUDK
I9/rAFw52MqhJxA0KlNubbkHZCvGa6AZtYtTo5BjznGjlkJEyY3t3IGMFOxMSVii
cWD0V0biQhCUdAhdV2nyS+MiAOzDIWP+9wO10d/U5Qec3mZJ9WbZFy5FlnZBEpJa
wHdnlQIFjbPLEuyMWH6f2FzSdEB8WhwCH72F58Wh1he7MuPTngF1Xg80WfhumUpX
n82AXcx8Rs68s5dpUg84yIEie8c686wVI8wYQ1cTUyPHM2MoeXmMeyI4lwNBOrD8
ZoQU2YyFDgqZnJck7XgaJrzIV/D3aOm/YWZVyWOKD3IQ3e7LF2REPNH5AANBaZSE
0JWXZpK0cDQ6Nu0nYUyALrNfzVWGkf5LhSWC0I6Ichx7H2TGASlkgBWhqbRsP+6D
icmrRK/BDYAHUW0FLEdr/+GFJH/R38dOjlJjvbgcz0gUatcH0gL8itcDuJt2wEIf
SgR5XODkZfLVHVpyj7RqAsrqZ4ihgRr8On/haZolbwifVEl8sSc8L8a149lK/i/b
lb252gvbBJwqz5k/qGlbo3xy3oIKUGCG42/JyGaO0PexGIXV315vEjzjU6lXv163
995zfvR4eS4m9nx6guCNCY5A0zDDbyRFSwN2DnF0y5NLrwG7y8xw5zpfmMIoTIPV
KDLmVuJ+fBfL4bXYPQ9qCI/rU0QJ50hOWWq1KuZqUUz/tqhweIw6IQY2fzcZ1aoq
XO2h/pT8G0nxW9yK/od0dQjgDxag3nKq2Dq2GYReVFI8VWdsPZndUrMU2wNo05di
0fH85xewN4vQBYdNWX/dzC9foUQZzo2gaF6kUMUfnpaJIIkyg7TNAsHjFlQ9sPJh
cOeGitKXdFcMKUcOuuHFuJ8DtYWjAF4geoscEoV+m9AgqFZ7lXkR8LJeqK5FAc25
1iZKIYtueAlZuYR8ykAFMLx0saM0IUBQHeDfVDp1q2OfmOLTdRR09z2lyzPOCbNx
ihjuPGPH56YKJoI0tAKQkBhNMpKCPRbLlJHHVyp/nEZm+TKb5ti05yhP2mCqU7DQ
RSov/qT6CQk81HtK2lk9EI75HTBX5wv9MmAVRtd3vs3un14sjhIvAyS0tsys7uDn
n5gGB1fcCxcTLffkOp5XJUiQO/f/AKb/ksGrBFkJLyzX8sSgAZLvloTz1ITOQxkW
lSHpw3mGTtrTN9YGnECZpGIcLNFJ0aLVBXo4UTI22TvRXPH6KXvTEP/w4kYUBvhi
vVeHzywakXUkJKzwYTRTQ6K3zJ7NPbE/986uwUhvjdN2iHJbKIpSadXJ/+IjhIhl
/RMSWL3ZAM7dQgH+haQjQ7/CE7Wono869/D0R7s1HMUeJ1vCcmqcCGUrUnTBdcnO
KX9YAvmMkCpvncS6okiLSZGkBIAPRo2q9/qyFqh7NvSsL+YAOU46nU7Mh0lCYGul
jQOYk0IyENZPuY+YIJdWNEEOXSrAZ+fRlYCOTHZoFKTEPjD8BMzxkGqQcH32HlJW
XlKMoqKRI66QJUo9MOPFHHu7bN4Vapk7ujQ6n8xG5PenkUqlIheK28pBECAIUmXy
VSLN4bYxiIWIx2YUCIPCs2wFCxCfd9Om/+9hvvzDwn+I+NASEgSN4QoWLji37UT4
hJ/1Ln4Y+eGRMNPDp0MFj7CIpKOPlxFlWlvuvwEj+5S5qwBD6GyCg02dPPVa4tXJ
2OA4/oH3hTss1s+wIMZ73d8V3HTN9NOt3A6Fm8HqWAGlllxoorHaHX3m4hPApL8G
OuBaHtgfZ3PAAG+fauZ/BlrvMIgtZ+8iKX81t0FJnGLJbATSQuTIZGhx9hgp+4FH
eXMvgeQ9GaJhF0SIDztBwQVDcGMkJZy9Ec7GFCV0n/+5NEfyVHhkduMeA7dZtM8G
O3VVQlawRC00P8cJKbsE0XXk8TwikR34xTIckvVeqC3jKYLrAtTCGGcwR3fA2VgL
ugfbXv/RhLL2L2kljfc8rs/BtolmPRkBJw7sf9TKOcn5SFK/fXz0yZzQj3SxGAtm
3D/+e6lYMbRN7AA/FHrxHnB7FzJvicb6ydxvDRkUFldMaabl1GwTH3kGJUNHBqv6
6emNhX2B7HpLC9xLS284RlpmuEQHk4jjO3N02TR/b4G1p5aSBQe43mKigVwfJhuB
i5Arb5NJ8zIMAoT/XxRtSo16yYe6+AHGwfDEAyDlM/wUNDJLrs09KYx7qQBLy4o/
631FRqKImxcgwZQYEHRJeubfxAxZgKHjhnyXEj9f9Scr1mo14Aavujbl6dPDyfKF
+ltcEE2Y+HRPpFvaaN4nYNNdHPin86rlGtGO9b+MwWmCSfVKQo9Q0S/lBModZtYh
XhJrDkiXOJqeKd/Aj3JGVGQagJKDitdmlS1IboWh/tIeQlR39fusRlQz8uOhTDhJ
oOTTBphPBkP9coV6QXyyjgFwFQVUvdMNZ8NP7+FdtxoYxPHM/XwIyvi+4g32lHzz
ObncqZNMBncMGLg2Ubeb8txFq/vs0AGFjllmGkaBDh2SCWDxtvi8r87ZT584Pky9
uoN4C4fCPtQbDtpEsDzvb2A/BeliWaiRKl5ncEgGp0mamVxtS1h41HVdKbAdCyYB
L+TFM7SXnNZ8I9vodqYpMlaN57TUV3wT5Hr9C2wFho9zhNlbRfbCyzadvwnC+8fc
UTFSQjo67cN+o2KRIf/zdWkD6j6MW+uiebjHe9wmd/1R6NZtc35efV3rYNM2CGCk
1UJPRooYMITEL/Gw2Qv0GghcFx3wv7Npl+II1F4gKosxO6LNCGFmrQB3ORwM7ddu
qsY1EWmRmu4dvccXCeR3duaPLTU8u7vV72H9DviuSoblC5RtnhGpO6qE7DQbmzUZ
GpO0Dcp+12zwELbuvUAzoBzxn4hAiZ8qwH0ieym/xdvJZsthGGhGCdm+nYqyfkF3
rmyVtbgMNm0z7Fd8yTtUenXMaSiDA7OgGdVR/0mJdUyFUfJBFiP3U5xtcI21z4xs
/BBP+Rx7PSwvg/LhlterlYHN4Mbev0RBT5qFxpJkotM7qd/ufBmw2aS3SxWKh9nX
Wndp91ftTuu704U+Z99eidr0d2u8ZXZwLh8v0xX9GaE1SplrPiPV/LQZ43Cy69Jg
v8jjDfnAtDa3MlOywtAXuP7hA8/nZYdMTfjSiuYZV6pDOsauExqEkTzeZhCE/arV
HF+qJEhAjEJnLdnaksPfhdobg5Xy+9aORC8YXObU7STO5/m3xTeHfcc605tUcwKq
RGDNBwa4E4OGfAlwNTw8537856tuEBgsJd+9OmLk5o0sFH0gG1/mTfR4RU3ZHQxe
R/yYsdky4RFzB5kCkvPcYQo4Jls1Q5v//1e4+j6sHiBFEI3ixN6YNTLaR8bYEz0N
9ejblrWjkafMD2S8Hj0HafBN1a7eneR7uwewNGG9JMouK0rWmjOejcOC5koc9yLq
eVloehqNhof4snhBN69YDS4osDwvLgFs2PQ85ufJ6aAKJnZDzfm33LlCv7VU9t1V
TjjMoSI4Z4fMfo0U7iopQ9a6ifFwnYE6GkqY2ZoUABtsAUM53OVbN4hPJVBLVRPa
YSWhjH+86Ywqvf2QsDaeCfdrkpr7gi4mq8QbS25LnaJyOjZn4d1K5DknLBQc9CVF
XH2S1ooJUCAWhp0gDga5xvqGCQdfLTwKxqB7dj7/p99NkzAqKzikzr7xAjayY/pW
1MSCizRkDQZeyUqXKgc//HJrvF19ClnwxVjf4jB/je/vly02Mhl87RjHl8zSCvop
wt8KOfr5ptIwlUqr4L6ZKTm3HxiMg8ejzObxtgy7QRa6RT8OEZUj29Z0GmkAHrbf
SwCkgvOWjGZRUhgZi9MJ5GIx0ged2PDVeZ1pU2ZXX4bhohiN7IZJCBfDaYUXbqvY
vTjpMmCYojtdoP7F/kmfkTNscFCy2S4hVhE3qO4yWPocwf7ugqi3GzpqZJwc2ptV
mg1MOAPvZ7vMkwR3lYLZTB35XS1zP2UUYYaJkVLT+HmF1sU/Y4ll03ZYaCQLgceO
qZo7sKtmHyi++q/atY7W7zrs8nUYNrMwBJWY+J1LBP2g/bE6Wt++GLVFkXRZRxzi
KMorQnGIi7brArECTnwIuDVeAqWVrcqdoq2n5uqTs5oovDjW8G2Va2EZK+HVQa/Q
LNrZhEBVxrUq5mwxHpEc6sHNnjZjPRym7KMvuHqmUlLpaTpd/dvK5FEHSaktxCC9
NLQLhQLhDzzb1x6Ago7AJV4dpVBFAoyd7I9sbIiU3/anZtUmK5WfHEwF22JIykwD
YzMli1nfhmbBqp2YCIjeCDzXWck0bfyZ1mw9zqLFTugJTi1tsH848M+yyQSWaMNp
2Q0WU07Sa4i3rqQXxASHuzkFYKhSc2sujb/D/KVGaEVwvnFL8CgCOiCphIw8sWJ/
3M4dXIhQsRifmh5FVXt5bJSCKkMi6S9FC8IvWA7HXxC61RVV0VujGw/YsdCxEc5q
3bicIjkGGVD5XpuXISkR2JX1lT9xggDkFjR8TFp+++O5+4v6jXGpB2s8f5YggCqT
X9d3vjgjUskq8IoOV5tc/JkVNogEw0yV6HF+24ZmPenBtMrST26clxdTZbV6kCxd
0zr0yh+9/AA16BqUyUFgjLdeHKSbCi95h31AFh9k9kqJGZyFyKuovkRrMiW/F4jJ
R3MGM+phfsTt/0lWu3HWxn+YC4tR5dq2W8fBDOjmE7F/DEgIBEkw9SI91IaH4gmy
YwJRIekSWVjfCqCTNnkP/QHOcjNULI3876ACivxjE8i79qHfVZWqlN1+D6zF0d5D
IP5JGnJwJmIdrVfKmpu5pdXKsFSs8O2LDdgp2TEt4wnraClqH0Z3eVubD7dpyP99
cWNyduftCOdJ5zW55Kdeiawlsw5BlTOPAe9fz4Re2U8yisJL1iIS17/MwV/552Ua
i/1REwaYIEJelzRMe0gBZIltfm0scW/HzmiAYY7o60N2UpjUWLN85nI9kpdNWJqq
f3Xq+5SMHmkK4Oln2hV8sYZN1/0v2DoAgRWbX+ZnW5K/XY1CezxKYwMmNA/6x6Qi
+Kscv2xL0r97/BmXyTmoH+MJcOn9PB0FOozDusdXm1Cx7mMV+FpU8MpzBsMEi8Zv
t5qHYj4RkgrUuU/DTCieztfFRE8gpK8wmFYvbHS+FRlkxQ6WYq/Kt0C7u/syJzrT
jCtVRjKFFvei0fgmnHSqiw5pOcQ10/dWtamdnrNUEXZsqTerqm0HBM5ebJdfmYl3
7YVYIdhPobjao7xdMsM45ElIrnFQnWDBmoi2rsNjdsqGkL9KO2jf5mMdEctU8MPC
QsKnkev9AVJV3l0afvxalLww4rHR5cqramuMcuc0PJCiJKCdBFYWUPR7ZXRHNfE3
PbDKegoc8BcarzfS4XEApCWYVO1JjUOMGEcjmRAXlyDVfGecanhVfEcvDOul41ZY
kV0fDJoBZDlqLze1EzuXfWyWDFpw6ioMR2kfb4DoVetaukSEzO/ssl6HhKdTIkSU
68LYh+7ewd27LxT1lpmtTzoh+TTMOW0ooG+TwUPaDzuXQZZHrORnpojsXPSm5/rl
HUADpOQ+edPZwIfG6lugqYoYlg55l6AkBGlEgxV/D781VcKTHrLfNDR3OaXdWkyl
wXKjUsPEDU0xii3C3g7BDUB6mlH4TlXM2MF6ojEEZm4L4TuksAMUTcKYgpBH4e73
OOaVrgExY+ZAOhsmIFsVe8PXayAxdBVNTuUI+JlL/r/xsVVpqN9TQrXGhhmtQApP
cLDuI4pQSYnOxb5o1uOOvnJawDJCorQK7JCrGcGgteSjaPQDQsRLP40wTUVKWo95
7Oe6lwhxGOrG9herJa3QF7rH3r0yYCOrP7WZNsHkv47bGIDhH75gsXUuyuDirmKB
TcBo+MqPoqbKvFXsmT22Qx/2/xuGKwxjrw6XniQhb1zc1ZcvlkoQdULS6b6Aeh3u
F/CdP2WvVzU6mooxD968WRtY0AJFnt4JG99ga87eE8YfC/5hGaTPm499my3rftYu
gTziwyItSqFKGVFoUtqpnDqepyyncMERD4rJj++oN/PsYAsAam1/GQyykNBe3Zkn
zhlqbLo9/+H5YFt9ktHfw6s8u/ycw2M73qJy1IUz+kdXcOaVMorJu38oQar8GAnE
gyq//OcS75CxX+xHONh0ld6i2tPaX+y5UU3UespxiNBho9O4/QMBEp0hDPzZLM/h
hWzaK5MBx0PdAtDp5Zl4J31zK21vdU66E0CCs9I9s8ap84PO1oO2DosxXiiDrwcp
OJsdKrl0dZlYcJia9B57kwd3DwuvfKA9+utLAm9u0DqHzSYBIJD9I/6mbcx9UyI9
DkULTf4452SDZFErdeF5WOp1mE6W7A/XCN2P3LCs414PRBJHPz2TTPoXqJYdOPYL
57iY8yhVFU8xXFYyvvFTuDNCoU0n0o89XlVXI/+IACpCuEWgWz3aUjsu8dUkAsL+
BeDvZMHBCwOjAyXDdUcsLr1vNRQsY9U+5O7ga6D3V1i4RygGx5BtdbxenoTDuVJX
qPUK3SeIzuVfjADSdQfXK+3zVyrBPwK+KBJPqARDYIqi7RwsGWSf1cvKzVtNaefl
rBdzdXzyREuiH3xDPB/o1gphtr+/YBsfDi5iEuukVAtWAkj8XB6Zv2TWHaRQ4zth
zav97U7YtbiZZmlCNbaohMyja5Zc1QPyXj9/b6TnlRJQGpqMUlKQgKKkK/Tz8HNq
FMcZqufUcfnLCPlxVxsVSxKcrlUFRz54VXBlaKUyxJh+1zvLzc4itYoBnHIQT8iD
joNEu8z04mS0Yn3DdReK0qNwVZmZeUB1U3O8GENvDo472pYhHeFoMCgLEXmKdZNe
kmKmZ+vNZFRcNiCS0/Q02Nh3bAONhro7/AWoLMiT3CL288h0kWbPA68/qQWiCHcG
ZU/lwzBmMC1oiadQNsiScDGYLXMiMiTG9AdLNmglftyCsu8BJlIbi3O+NHRYQFMe
A5V+QGVoCeR4VluEyYxHscIecRxg+LRKsFasCtFaT3/z3OqQs4guDuax3VhWb0l3
M2f/mgYQEA7O24R84HZ4a+jv3OAKD+teK+05L844NVggu2UbN5cEtuCSxQmQ7kPb
uSoZrwe+KEKvHHkwPdZU2CTG4kZeFcREx18oWDPbPzDofIO8O1W0kthGE8S42gty
KjdztP6CUAeJfac6oxT8Uq9rmzlXYY+V6bHMiBpnjNefvE7JOW1lm2jIs3g3aYNT
P8tgP8lLeg0KxKeRL9WcdLYAmu6v/sVxmIeQUfMfj/2W7oLUs7hF0f1aSiChtqqL
s1p1kCuV1H8ZxSPcNxrluzi77/YT9YuC2KF1PJ3vNmcxPt03pILMhnIqV3Fw4Djh
YA7yGcqiqnzGpuOrZA8kFHZL+BwQWtoWZvANJZLOFzH3sAdMajABJj8xgiPr6bPG
pmsc5UFJA0kq2ZvvGXf/h7tD2TeNv95rHVCpGRqqdbdK/93LYPp9BUp58t+F3euK
tF6tEV1Kz4B196GNPOZ2xzbe9m1N6+Bc0I1q42qJWCvsiKT3Nf3tlZWJRE9F/DIB
KrlDVXY9YHJWgzyvUZ0PdggX6+rwxH/W2orFaQC5G5RHktlRXZovPvJ3E5sxdicD
JjszRU611SKOu/uBf43ta+qrVSimjHooN4VZz3r0eIB76fNLpCoXzhW74S2ny8DF
vGVVO4vgmGgnjrOH3HKpuhuz4PIX14j+hRLhT0gsZ5142SlkfYLnTgoh+wWBc0fC
C3xmbTXj8fFNo1u8S5WtGE09zPCVxs4VlNYcFpd9PA1ngIsRKJ6gfw5ymrohoBDD
o8A2H5rrKwta7a1UZbkFMaL2+/1VmtXHGOk7cGKHb4Nkgkj+QLE/MP6tStyhWoLu
HFZpHJTAbazDQFMYOI88AsTXPI50Fs0w1DYN7prqVX0UwCt+g+jnp2Xdp54xtyYL
bH2RTPHeZpEGPtlI2UAuvrfQN3L2hdRYYS1hYXCdzhdzTCtJvJ56hSOr0xN2b2YA
5o24NaY9x6vJlhTu5rrZfwfZyRqezA3uUiIihs8fN4dU3GvckIWCT8OL7fvBdJPn
Hf+KkZw2XoCHIUvreavU8Ur9tnkdDjFqfxvf60zf+PFrmFfHBuDTcqOfL2zPyfA/
5blB8f9SpJWbHZRlwCCwUvDByJsu6ecbG1Rq3jNWJaJitdShnuOEba4FNDX/Iph9
65auZ7UNAK3mLeZ/wE14ykNmqVF8BxMGVFvrCYrK7UX1KEWdtemsvb1Af/SjIrqZ
Bhrs8NpTnp2lvoFO6rDwKyFHQK2HPRmzokJbTuHoWKJPzl5RY5mZm2yxRiyGDgI+
vGLlvyfEbrXcHmAFjw2wS+7SONCr9YWqo+S+nBpqu+ElRcI4sU4B1IrAmwH9YuaH
fHZFDUJhR8aCj+byTZhG4PTykqqWxpnB3htfBXfxtKa4ZqRzzARro7IBMgUKFN1d
rv6Hthiw2zmK5XRXZEFF5n6+iOtMwAf3oSl4ec54Pf1CMfnxyiE5PrjCFEywzVkb
FvtwgklcHsIrwrUIr7EAP7UMhAb/oFswsDd43NzDIEI4Pipgogp5REwtzWzggWzR
gAiabhr9m+UFdeF6zRi+eKTFe+TCUfFcRVZMshlZODWtK+hKpoky1S3SmjR4/4rj
1c2QPgUN65IfnhGlUrDu7cXOsy/TjJBvuItTwQ3RdJT5pGfIQtTGlQF2T6vMSauY
DLrpc8081xZN0bTNZDmeIkP2Ryf1e8/5zS1f1BK9ZqEDlCGqdHpfR+2MHkjd8RwQ
DcLAEmf6lxycAGWD7VJg1YzhV4Pu+H9nxjVyxmJs48xjbOUIXbg0zKZyBrpyj2/f
+aTnauu+CzMeVomfTovCUjHJ8VQbdUIz8RumB2sBrB9OZyH4RAorlWEZlOi/C+1C
LU+LNCmAYOi9E/DMVhpK9nh12pEPx4r6UhZjMapdLtPZgsX7uQNiTO74Zt+vzkdG
ME2Q0hKVtVWMgNKNlnr8RdvJlphGbQw2Yl0ZJk2bU9iyhjxrGS3bwbwEjQsmzvjv
7R/t2r/t6qCJWTZ3lPD5RlTwTlgdLr9L5RhKXY9TePbBG8s4Y5IbnCsX6FYpEXDE
JAtIUkjeySW+Rg/Dn7cf2l7itqkpAvNzDXJ+CgLix7BOR+3D17/Q89eL2O5ai3ss
1y6aElkt/XOsDkyYDVTsltDWTcoWpaY/cN14h+ZzdUN4t/yZcEOrG9WpGlaWNQ5L
Um7v2efRo0K6jvwgN7rFwgkBnDXpHKmDnBG7VE5fnTfuHEB5re2JqHFk/ufyArFb
vfSDN8ZfskKGwE0cvivtTXWf2k2RPlKYOsxFOatNgxTmlHCx3l8dERabHfbFbyqf
2V7sRQUchvYZjSLSPRIyZpZvuM/J527l3ghhi3yRPAJY9E6P8lLzxZHM3VrMv5Jy
qndw9G4IZyc+aRS6uqoV8sl/ocHGmQkcDbs4e7RGE2oMzI/j+51cmaHBepnxW1bW
8vSMKWUpOix1EqIxwjCDm12kZIaV2ovOhLeIjFTDT0nvlNpXTDcu5u36MYlnqede
5KznH2LUUljbeV2+G4ZmtAR4ZKxxFpzfTDmnk+GZJxN+kNYsa+UHZKtSP0jMamdW
2l1pw7yd3SofEw980yBMgFajZWWyBnCId9m6Cl+dCMh61g8bPCf9Qy21+NT7QRvV
WSS0Q8lX2/5g+u+NbNCjQAV3ARcaCVrjNnzgzlcnRMMwJe0K2KwpINpzlcyZ3yI6
nGkviMRIb/cQvwjO18CoKGnEklvGEAJ/8Eo///cT8a7ZnWqtVxOzoW1hHUJ7vUEt
m9GM7Z92JzrSgFuPtTwtrtpyyWVw4X3toQOMiZjRWaAcGX1y+w6vv8vKKmiJ+UIH
A0agc61QF5LQ+XlhaAbc7l5r0niNPdhf2KhL/YpGmuSw0or/KunlsV9xSqKWsoMp
5NUSmw+2gFA1lFlnnUY93jTpSS4A8MxIz+nfFcgNPLGyM4FUcHP4wvaW1RIpnlT5
Gdwrwq7RMcOnsY5nj9jFdKYDNfmRK+mg3fGpSf93QlF+426V8uiV77S6hK6oZzGo
95UAUeqAGYSnjPYniQWj8Ij2998rKKvO4bQqILN4KoUyWDKrITE/r42gaXdwV2VE
Dsyw5UJAPuOR+ukjH+kyb+IkIhz+0ZSMz6IFL12XBnrLBDD5DN0ff6WcLBBkRPLX
kICvDcMKuquWYY05v7Xaj9cZi274yyyZJSkin77UH0/wMKVinN4B9OaHOIbCIr3b
d+5jWdjub7O7GWtN3rNp5N+CuriwNT1zUbhFYsmZZRKqD/MWphib2ml3IyeY5Q3d
j9/xxG/PBTuW/kGSn56E67zGMGJ4dUetYwgXM96Q4MensSK/PZ3J1Rulm7mVaPzt
qqhdZRAlg/PtBHatqEY+SrhQ2eF2YKbUQiw+GMgpFgaojyZHHb6KuPYkMgmKewQs
7z8r1J28BHAFHfoHCE8Z/HsWsGJf206SomSY2J4ZllJmsmDwxbbsYgk5Rji4PeVi
MW8M58nMi526+V3wEICeKQn5KSp4+uVFvLx06/CfyOHJkXKTrOxVyktxA6OvwRZn
Z3kNodftI9R7wPW4HfWrPb/IZ9juUOa4LpvPEs5NdeyK9nISOnAn5vbJNx1/cWeF
d52LK2RdVNe7NFhNVJ7AIF/gUCZNXOutzFwAyz5I3ING+QF/+6DkQcWryac1wlct
ladVWadLlOewMdT2Q2dxC9iAU1s4A0DZsGxsZXNzL4BLKE/Gm9hJOev2DSqNTwBW
MBbptQYOJXrXMCXPU9sM0bgYT/gI3z8yQPKH8a2PcZxKBeMCvyXJBSh1aNOrQiGr
AJDpKpNZsj9Mz59GwCj89YOY0C9sZQMnW7BSAqPWj4rxYKSeyyhH9xvc8ll4Mx8A
CZByk9L52aWAzJLDAmZcdPJXyfhKPVz9FMT2x86iqcZOGxSNXQaiRzOYme8yKjFl
LuwRHeoszrBi2AzQ9odaZFLF54wshYU/+mCT9WaXvnWHZ1FCMxbfH1ZWJOeDKEzj
HSqolEQqwhNbKsZtz/aAMkLNsHFmuhPIilKRTvkDGl4Xv4QhxO4u8NTU989JowFr
DBRhjOPE7OsL+BPPHDkKCgIa0Ivul0im3li68jjzkzlILM5VizxT2xE9qN0AeLXp
I3H8VgRwgKGEsWBBtjyjS9XU5Rrkt6b9ylTyWe+UAd/N4yDWeHXWhd3yR/gs5z3I
wqaGXrzYOpWNQFcTudYRE3qibC24J77PahJ1/N3y41VGooyBaKVyjyjR3pDl2mmn
rA8QpGJrZ6rT1tA78ef/vSbILiYV66T8qcZBA6j7E0+Ir5iCXFk/sS23ceXnCtcz
uqlk/IEk0ncQqZIgg44+dyKZqQjXWpvuwYg2lZhbqA8LAblSTqUOP8C6uuU0BduP
cnTgzqY1ol6kj6B+JmFdVMCeoczoS8BY6HAaJaIG9PvWme/rv4iDB9P62N9wDx/e
u/HleG/NXph8lS4CpzX3GV9VmM3bwaT487sD4mCZhU2kVdCe017Ne4fdK5kgoXSS
6ToimNvl8m25VVWpTY1ndXuT/HkzG88yMLKQcUogI7cxgOf9g0C7QOebwAff71TW
Xdjk/AYKU3TeIOg6BEWvhYLLZAjGXVss+da8PdWr/7D/1TnVLL8OOwQ+vb9jQczw
spxt2nFP6lXc45l1TEgsJdOUdjYlsj7Ap0b++//ly0ve4+AFt1BNoUJ6gCCevKph
ndzFkM2K/Oe1l6nrCYdqQhoH5dcMWdw1PttCXDev8RMp9ogST9Ghkz4iaubuFFMo
x7Y1zTfdUbm6dh1XwRio9aIBL7+dZpCHB/cx5/pgBgVY2IuWX1Moe6d4eYVcEutV
afugeBCaazMhu8uNhdScgfCtS/ZGdMAZK+ZMTCwlUrwDIS8GE2JyJTY0tRKhHU2L
ca3/X3dYMTlNaPFIy7JLEVJywlS30yqXDjR5PfbSf2jFn8DtaWUvEXx36PVt4VHX
UVrMmNPukHXhqO9okV0KzVOx03dur+uSZGTRh3VEqdRTvhTMycG2eYtZ+NTUtzmb
O9Dkz7wJ9EhR2vrCVHGUG/Vi7d34rOt0Em8UhNGrl/tSk7X+/xX2Vfb1bbp9ZLWI
vpv5Ige9kKJvVidTJFxsYxk3294ozs9mzcdyrrtSVPhixSCoYUaVyS+UrSY6s7iB
rrqYSuX6PjG78zf18n3ECig5+u4JNrub1n2tFbIDezS4kzfq6yT4GqY84NH+GPQy
FZLec371oFcBTvvwlElxLIIIN+oIjLL8ZpRTx0vS9speJ0iBKlSNkT0x21eRbMKd
NOh8ChgjMnIudbtrbBYxkbGtqHpwpM+MhkJA3KK1jrYQBJLc3fKPATdhEP3TeKxE
gTaS9R8yCiFL+e7uP4a56ask72t0UBWXIfB/KZOX95o3UwLoIWKbcZXACK04lqQ+
ywN5cqt/pqcv/T0vWCA+50wQ+RlsvCaN8TYKG7nSS18NhSBj2RzIENP8TQ+mEqaX
0XHIpMFAPKs8h7bVxOQgs4Cde41tXs+aQNQyY4smVMp1LOkX/9Cyx0vDvpL6rVbs
vD+H2dR9t6TYqaozdvcKcQrjBuI7qTHQsQyS55h++JODZitl4PA/2E2g5fPGTW3Q
lujBArO5VBAOGW87XAoQ1lcAqYbVp/OrEs5ttIos9LGVfJPmMSBrH669mSAuBBt1
SaOrOgUg61n7BI5LokQRrHzbSnQ6Oa4KGACAwn/o0wCAD+qSGdVBzz6i8lWjEIAf
WIdGAN0Lisiy3o3/8dJ104jiHzWkwW/w77Yh6o/h7QFb0tMFd9JyeX2F8VM4iC5h
yG8xxBe3/eqn8EPBlRLmPklkWErRsm2WkFF9icouLMIMDyIHaTlRq3cDmsbQF8d6
I1NwqyA9iEt2gJ5qXBSY8cDmVc0x3aXH27RtFguaqEyc7niP4MvKPpo5qNQFW0ZM
tSDgqEBGYi+fFhOit8Q8b5wXFBxHUkGXmmS/6s3iG7EquvKvXxgVfCvZ++NZv+q8
dwETQllNpFUHVlag8a4LdWCojoIUkij94ycxD17g8VHM5RuH3U8cb193HhktuzNT
ZhjCc1C8/XfLmGr6mUF1q1ak+3sN3f0QHG5vvqGiQav/1apywrlaE8pl+lQFEJS8
NlidYX9ESdkF9Ivity4hkcD41VGq0vyTUhv35gIF1UblCUr4EacvCgOBTibfDd7T
pivOWAxlrVcvhq3CJPqF3i0I1u4le4BKYS+XkVlLnfWWaYaWu+tcjJavIaf2sGmu
2W/JTS1nsIDN2k9GS3ywuvOlKRLwbK+6SEZ7L1y3x7+SRj4MJaw2FGlrYXJxKTHp
bUNpUp8V5/XSmyvXJ5kdE0O7CRDhGLLwIMTtE8TIqpMU7xWGWi8qkNnYoGKijmwY
yW/Z0jxBo8iPCZG0gX4bjhmWkm2S46nQGgsDnlm7ml6zIWmdzbXNUcsFWTpqCpKK
hWDMu5JRYDR6ItwXFDCVk28jXqGc+BONzK/hPRlhnAbBo4sMjUx/22yyUedr33wj
X/3mox90EltesgdwKPjV1MtDhO2C9adXsbfKDtPBOdQvqWCqSPxuvws/NWDrz+ei
zZdw6BWq1CfFdlhZZBHcGRyBN3Tlrxnmd7WmL3g6KY+jOInaieT8+DbxiU6ewiv+
b3WJd3niV8Glc1AgWbuTgPpGRcpObbNXQcUJ+xhzJEMOH6mXzMAoXygfTNq3vEbb
fJPxGmdbvshAJODZ6NybxY4Eq2Z+YY1/IjtlbquU/Hd5OJT7+vLrg+sV0G3B1iej
FjasIoL+SsNQEJQPq38woFaB9Vtz2DqSsyVw5rM0CLsE1akRde8z5KvNy43c2mdD
Y/TvrL95f2U7wHbfeIAPwCBdOxpO4GZx9VMqrkdfgO8kpGIu4UfxgSQ+ZIk2fw4q
ATta1un1YSQJs6bn3ZKm7fWmVWkowPnuwUQZ8lt6TR8JzY1FvdvDAJcabawjGGVF
Jcgmv7AqozqYLVhFf5STPagpeN71VrrPbcFGTWkZwDtiyhVeKyomCvAJatugVC7/
I5z5Q2FYDqXM/mdDOKwCwKzfaBdxnPFklQHZMzAsZb73wPCIiINBmrE12NQ7axkn
nuglFzbchGv2iJ6p/+s1t2hfwJU8pEVw19Itni44tdUXEO1+Mc64qofPKHDUFJzs
JO2eg5QVeA8dPQFJzPgNUVkqnE+UIAxRiByzAfiijdYeGJW78Dj/jQVtL2kcW/6C
1MzcY1nZ9iSpBH6X+H/FH1gm/L+n5tN2d1sU5CbH9l6+zns2h1XXgNly4hGq6E5V
VObEU50Gy74JRB9u3vWpdrUT7LlZCAXq1HNed8awVYGUb2aJ3VDbeXzzC23F+brU
/HKbmFdLaGLiCHDhurGZkbvzUqyanPvY04w9Uh6K+TiSH7r630iZhEe0N011o+9l
Wcm8j+o9vjYEqHtM+7C6pdjL2xk+ssNvUSbzS23tgV3TAYCkFEZm/gMya8E4gwyw
+ZyiwucYuRi/3gv4pUcolyPKEVCna+Dl/6ymgJH0Buu6tkGJXkKgQnVQLftR6Q0A
uYnaL5O97qEhN9vr6Z/ZuHq4zNl0wazDMcE43GhomlgOCSzVeZqpzCl4g6b5h2kh
Af6Y3UXdWLZG+ZowlNX7CmfMI3++sNGgmyDJnTdgrB4OzUPxX2p7ZfQMEfWgnNcz
7hbtuAPk+n1f9ECWDeUr1hU8dXwF5fSS9JUPLmPPkFQXynDE2Stb3OWNcFgVEiCy
Fy2fz1IfjI1r+S1M/Caryq/GM2a2hIYQyTUrrUEXtiQVCrlVItTL0Ied74Pvfk5O
iEXcMTLC7AAsL87ZeMdCIR0WyPU8S9ORepFR3JbB98u4TvZKmsWWjZhb8/zqMr1/
wbgiG5nGxCUc9VI6fiYhBnfWcYUYhrSzUJHeZXolTcpDodzMiUhpK7TSw24iSMnT
UmWIKFhxtUJTg8wuJ9PjiC988wNmrOkDxQau9gGlNu5V10jH+Z0Lxygw4fFGum3i
qKxrjXe+qDpAnGP/Q7nnSY7QphS1MfqABgenUwXvKquKGxuzDiOlk7VZ0WNx09iZ
CfB2vWKRnKO1v3JbWuuUNrFeVm2/PyAuhCgIfHsCjUJZ/90+wvn+k8uu1LFfVnsf
yLagDLgW6nCjqtPTbjdREN2adFWUXjVxaHmp80UiCJa/Pj2JHww6YgJ7FJeWxW2d
edAWgAILlVnTCACtYFXR2A93RB14X2LsEa/T2Re8EAz68Q0ae1BAKhbw/VeARZyK
UevPo8Z4kunZYvpBNzwcsxgbupbRhNp1avhzBa+8hq9XeIqJ5Q0oUv/rnNPeUZiI
cZC9/143KsQ7ttzr6/Fsvjk6LnCudB5xNhnHhK0Ace5KWd83QBs0UFRi2Z/M2iXK
mSCbmcSHEevWU9jS5AuFCwEeCdKeZMjjm1Ovk8E6MwxJ68hb1iCS8Ta2q+uJtdr3
3ARW4VYHpPyxrnhT4LpIfgpFdOWAUbi+1/YF+AjT01gusgem3HxxE8B5ukgNqEQ6
zC/9xhOKvQNqv1rI7b6wg74H7Gz8DrFMCFnV13czRHFI9byryvaO99bL0bITWvwl
CPKhM9BXmYPaG8wQFiYR8CYdWuDcESOMpTz8nY4QVbRA4xzKnlC6vh1Pjy/NN8hc
WTsBE2LQeeTTvW2zmu59+BA3G8mahkceGvthOv3XStNM73g8sxzUYX87F/kLAupb
FnD365SIrzY+Ln+k7+ENfWqltJABcQrxqbHWUV6gTyPsJlTB6+WUuruTNeQtjMKw
Rt7QyG1sLZUqvFB/QTCSK6Evqr1hukSFjqXcqZr01rPIxxPLKHPS9hHEAOFMwM9k
EJGXc+EkljUXRV++/tTB/6mxdxQj9ER0n+xzlNWJr4qIujpKFzQempnD1zWme23/
0E7aV0PJxoA5g/V8J7ywBM4b27F2uYqmNAwycwLqRh4gdfcoMqvztu0jVHRsfUeQ
zCAhM54O8uB238wXm+UpqfSarpJ21fb7ld66C+7XhqwwY+UEytAFjbhsmig3vk6N
84aRGwKxZ03hkUMshdP8xIDaizET6KbYfPZ8bO9FAgCKSp0pGY0aB61Kd8XdsrzX
VbR1BDtEOh1qkJIC5q/FmUN9GuqX2Jux06x8FreUTBJsy47V9PQWB+LV8WMno0bo
8KR1+Y9YEce4TLi4MB7ojT7WKQFPc5Nj0En21W9yYi6JvJPcalT59l1rtuMNZF9g
tUUmVLJWRJOU/Yyi5KAUdzM6C+ZqxH5LviZGTyfv92mW4xjGfEbSfdLMnEzOLX6c
ib9ayWLtj4/vtKzuNVQW4jIxTAkVF/X+0mRWDavDHdp+or6bFVk8EA/bDVD9hbSR
EiS2j76XOkK3mpXD+qSQJWRb6XSrbRc6m8rhTHNKBIaicwPvdp6OvSWY7NTY7Ujk
Q9HrA7+Tu/C4hdu/UTxDkmchJKUzZ0RVLTrvm6RMMtCp4vUDeMjXK98FaNZL7w/r
pHEMzvUFej371WsASK9F9Rnz4CLRpyDSQzzsjwWrL/xcGbPBRa0qCOFbteyZqOAL
GCTOCT41lqUibh8tZdF7i47xosvfP2AwDqOVX6arxKPOMzqHPzhzXgybJdHBS1lJ
Gr4PBzyd/c85IuoJJ2v+RQ+hybGinT6sQGL597Kb+cpJwwM6SGNDfRdHhsra0z8F
6TQGm8XbqbLHYS7FlwrJsFYcVJFGM2D1VvN49HtaRaMXvw6EfQthNEpRkPYZVtGO
38OXCQ7NAm2eNGwFIF59UZ65on8fDXD2mSpwUO2xKjP61n4MKHxqmcJ3sPACUFNg
FOKxhY5wfj1jJ26VMDnvXov4IGzk2SWjlER3qCOOOQK5Mly0wxA5KtzA7+CpsoYi
cH8x78KJEQnHQ/43VTSx51krHVkPkaZNagdOQv8AVYOdwbZe60E+xppdr9klrat+
w8RAZdHKjMn3N+p5QA+DnxPNEXCEnNc9BfjuDk+zSv5tRP2wSPb2/MtUNCVW9l0U
ys59w2qk2EWWLfYzfl67KlBy2La+Ez1VBSqpENJA9XZ6Y3VyTQXs5zKAFclJidhB
ngNtArV8m9K8ddaaT/e3GVcczCeEGTc/LpPVI2r2eRPPMAmEuSKi9ZnR1x1QYiOq
3cTJWlettDZipCfWN4oNkCOghoM0GdCM813A/tLK9JFuSH3vuBBJs5YmMody6ks4
zOKRwvqSdg5FIYM3pwdexbLORWtnNqYMCGqPq3PLsh4joWHx1JCB1g/hIaRESfRJ
N4qpu+J8Oj30AY5zqZcaKpCb22cWy4dWu7x+4wzM+diO4HxZUd7gUTbaaodfn0ai
e7hulrs0HoiHtM3VxYtEHoJ6BGnJvikbgWrMPDWxdVzNCLdxpRrb+XaNKIcYHnlJ
qBoDqRE6UIDxHIh3QId4xKqPV6YGP3NOBnwDxLZ12S5PblBTsP+HV6j38Czr0SZr
r33i7aD/+ykILyttGn98c3Cx2QLz3j/W+aqOxKc/PxjfEOb1LkonO7waSPtnO5Jh
POts+znJxHCdAupHHpDqlfL7oBqF27o1hYRnWx/ltVGGZ/IIFxltNupuyCwREm5m
0JmEqRFgBhv0OiOBweqwpt7H5utv1c25e9fVaH8kZjgDd/LgmQtxLnuk0MRmaIgD
VZ8z/buaHeKfiLjngmipG2yLUYocfOaN3d5CMMvCL3lttUm9FhjxQE7LrSirETFB
mTtvAxjYDpsNBOBMbdP/+lR+G3/NW8M59rhxiY95NfNeM/90PTEZt1sb8FdlbKV9
zFixpUpv0JQMzGnJqXKbfzE9fji5hJt+LwYVlKehtZAN+U9mVYPd70J+nNFyl5oi
IBd3lIzqaiNdRwpgFLYr89UFPhpclMUs13Y3IwUpwrKcl1auX6UKlwzeXe7e+dDb
ZuVVB2YODWrIXC1T5Mve2/jhbjzeknp2Trvd+JQjBOxPYA9PGBQcQUaQF+iof9td
IwXDKbs1w2bwrePQnT0as6HvT0v266dYtblkTX4Wsb/StgswxdV9ZciqYmnRMAx0
gIKDrSUe3jj/yTltPotSRAYFJo8icnlSWC7x3DEL0+cQxh/s9re8MbQJfydxBtfw
FQHpxsAuHHGQ98O4TLffpNTipOcz2lQZCg4e1kj3ExWvNP6jz71lI0Avzshscdqv
CkTmXLACD/W69csd9ccQyE6Q8waTACxqmQws7gIwakKoXwGg+n3/XCKoWZH8NpyR
uzkC4qnH/058pGvqf1Bz4qHGa2wyjPYJu4uW/DJ4JjH5nreBTstClEATqqvgoAiP
tp7DmQ/DHsrKyaROISjh2RUzLbxsG4NEQRvnHk+vzOQASxxqM1dUkfip3FEci1NF
LnuyJx57PYLFOtXakfu6/j/nKZakbXmV+vcbvMmq6QqQXLWL3D8p58AoQJQguADt
JuM1GgALNxMCWHhNA3nUAg0x3wpd0YX2CWqEyv3B2OJ3lb72P8pLYod5w+qHmow8
sjIY1u9AxGZBed/kFR7/hBrQLT2dMiIwSQ0KYjr5YYhjKw2fSfQDSurh+SvewRkG
dihgr2C+FU/+uqZH942xAoA7f/6iQMFKJAGlyINcS4VhrTsmP4Y1blgqjRUParGM
vrLZ68O0J//vVBYbwiuqYBeNY+lRqsj+8Sc1LNU4kB2a9KkrVyIYGzoIyghvKtBr
w1tx6DQUDhW30pqC7jhpqWl+a4yaJDa9UzXXqEvdO5HP/TmDHkillvmGgZpavZJM
yKxAeSFtVOMqRsmyt/ZB9oHzfujC5S3yF+3xFJT0GwaAH/wmIs4N+FwSVJUssZJo
rpWrJWm/atFTIGWJq0d6YEqL1gXiXqQYbK7ErNQ0xxLwrc8qZZ9C/yWW45QWHjlP
5CTXVZnV/U2g06A0eFUalXEzlCrXyuoW/BwuVOyS8+gkNTRR/rZmBDoKZ0Loufvs
6zEVmTbzmvT5KHtc+ZWi0mKSaj/EueH4EUgKgZtomSI5DJ/pABk0mKhNm1WPkL1I
W/28vbH0HXSxrvApIQ/Juh1AuXDy9qGol5578QZn1LjoiTyN38Lo3/CHuVVjHSFt
/TyenSt7ovcN2+SEY/m8k35Bo1sMOuEM4wU78jTT7JaDRgoq21onkQs+84W5o2gV
7PFJsYpgi5AxtTQDK1cVpxP0ioeqdr3bUAsYNwRzzYtMLufhpxOLlZlqVNdRPwNh
lS2+nXGsGhPaCMgNG2zSA+Hs9uJ0WqW8YkJrZEulUrdgmcIQALn65SMvITbfdZBn
P3DGE3IUSlCps2+PF3jYBfRGDiHwlvKcCo2XrVb4Skw+ysWAuSgFyia94j4e/u6A
T56kf9kOP81y4JYXj2OGMST01+UOgJe+4Fi5Dz2662XP6p83Kz5sFNILnrGt+ek/
MEWR6RYW4fap9sl1LVe2hvPzcLVV8Tz27IYNj37YNmErbCEXX0sZ7/qGG+mYfi9k
jVj9wTV6w9jKAvwOlikZfR4de0uFPVB73s53fyVnXtZ2CXmyPm7xwDIdinWVNUPh
s16DU7J+PgFSpcdye7JM5dlNun7jtNE0V49f/2VOBTAJQLaPc39xX6XPpezxtSip
MSGtGTDnmpzYWBtz2zUJUao9DrQjzOKzNC2LVHtFZoRn+3OJZCe8pXfW5dDv2TDR
hddqmDjezW8OXQjCDLNv7VLOCmDG0Kx9X+AniJugX66XDOPobSrMPvkHkgyepucX
YN5hvWvXnFpg/6O+XvCf94ry472l9RLrdQFDH2qxsoMPI7aTSZi7mkukkJu12uAC
GQ44rXXIm/vyW0NgfRYxJkFA2FnDOsPPaYbnYrymuXbiq0WrFZNE4/fBqFFRiSZ0
zezrY40L0bN15Mx6aWtUfYrA9ZIScjOie/EYoEpk89/oYuIHfQsHhLpmxM1gmyVF
Yf8AmO478+CQJmbXBO1g/YN+tyEqpsxo1hNyA25HqtTi80juRk1PKq+MFShN7Whz
l88PW+hYmUwlZneAo0KkU8t6096XJRGHGyvZiB2wG9SGxv/iFKM95HpgvbAxlsye
JC0bk75TTn2BfQPmZcWyVp2RBRvbpNjtL3jqP5p5GbxpvmFRyzPNDgyFFX6CaZ7p
hgZG1a+5QSJlReQ8tsV+MO4uPVJRqjBPHM9QZ3kEeTtLULe7l8sJ2LnZH/nF0laK
t7eZx5jOodfmE9f3FcpoHTfy8HCWcu3QTTQRtvajFcHfEFyXhG2pIp1XWkdC35us
ghZW065zBdIFfjVyWPeLE6Pc6ZN4qM6HePs/rn88zqqnxi4OlyQAyQOXJq2Hkbs8
gOqQYK7Uxwr1nNTHJafLy8RKn01pN2uz6iDHzH1MWivs7SxfW26f+xwzSlBc3NE0
FysP1CWZ+RFAovp0zGHTmEbvh48haojn6njV97ZvvGC5pClcgMioDkoEaI7C0Zse
nmGOYV6BrfWkU+KzF4QogsjFAs+VytJaRt0b3m+cQ0N5XabhR6KNJkVpsETNQ/1t
RDwwBHSPF1ni75FKZvCKs2wbukIJ3qoo0I/LMKgtL6PlVgqcZ+wfpX/etZpjJTuX
9zlr0R7Ee+IIYY02H5Fhm/NiWS0MNjzgtkPj7ijnjHmwvLcPWghvni7mElmDBwwO
8RxT7D/yTz2cpmnSFMCXMVJ7nwQVf0Dx80NifttWBLhVfaG2BPePKnTxeXbqdwyi
neow4txG2u7GHpFX0ULcmDUPsxf28hifCSxKxtKlBknQl/6bns4J5jghYMVn8+2G
3Q2+9htSrrdfrGhHWyFdwh3I9S7wfOXUmUSxzIl9DKI7MBxDAigwWXCCiq+fv4Jy
2M3HV5+4ZPqWztPn1hhfJXelHWVoLVO1hKXv7VQNVZ8DCKuax1mxeXSVo2eE/KM1
fVew0hoRdUBmdtIElsr+ANvseLoVrvbs7MBnNIAIeU0o14otHiklmhZv8olaRpni
GQYxZsRzSbvAVIS4hBg+xQBq9OjU46tP0/jLa3mbIKRhOqGAxLz9R+yxwg3ihPZd
EQyitYik+WbG458sEEpWR6N15r+XL2P4v1qd4do0PzWZ7TvVdFXchCUuK+AaFLfF
jrSPGiRY20yJdt2cumk2E3Do/Gvwt3iTAXwzbUEXLFX+7UV1L3LIv1Vn3oJ8nHH8
p59CQgRG87ib+TFbTNsT6Hd1hUdeWpsaGsChq6D0mObq/p+B3Rs9zFqgypOB353U
TbcKMoe7f4jFY8LvP2Wv/o/X0FMo4ahIqiI6JW92SdcgKO+DeEPK+KzRaIqga5d9
x0Jdg/za76gQw0WVw3ihpIY1j9MxqChJPAtPXSTBiqmf7Ts0FTPgey2RydwFCe+I
mTk2FjB42bLYewV2oxlQMDvLChZmGaGv0lI+pYeqXRjNCI5jdabXcvwJyxt8M2sx
PM9Uc6N348eCMCdTLcw9t+KI64tLKPffZbYCWx/VIU0rnPzTwZ3u8YpRFE5n0Xid
UBH2KuEtLE62tmvKJvgi9EwhQ9Y+vEA7PHMd5w54z8ef1irT+sR0/YDy8gdTLgYe
vtE0KldHe0/wkwWGE5DKbtfqJFJzlz/Q6hljC1esCaE996HW3qtIJbuiJShl6n9+
fKKYN78plcununisWCGEvuSqjmsl9sVWS6pshNYAIOR+IKayhVPFuuXrNW90t9Pf
YL0Sldwth1ncmMyT+0BGCG6eTXtVu1k2G0ltJL4LrMjDs8dFbobP2NwNwbTFaKTD
HZKEiT8CUUV47VpC4cyVijyY3PJE6V0RfDIATLc49LXs1Iw7r3XrM4SA5T2lLw7v
da8ZNpuBhTiDKa/2VYyLDRg4NxM3cWSCZWqNDykKH0uevC2kCkIYk3DzKEFxfkwx
dBIi6sTB56P+5m5CKn1D/chQIRRTxddDVByB/8iqQt9sBnyEoNbWbsllzyjEGOP3
6JR5ChNuugp7KsAeAtVbyf4n5trNFomD5mnKnPp8y6SDe+pNjrfZizsvFdn+o6cI
3BmgpQFM0+C78hT2onezd8ZM8u3WInKxiX28AG3VIgyAm2bRekhpOtTxU+bhlmLK
jLSBQT60eEdQd4z0D3BwXTJvvGErmegx79tVwXKGB8WRfMK2JsxDeyuyra/D2s4Z
uSujke+YEN/0ZCvFCzwHlcB611v3b415ryoClf/mOcfJlX4mDc7xZ5RcNdbL/R6v
GIRHDAy0n7XHFwHRwFhbi8KO+u7rLWd7R6ewtHHt7V/VvvJ+hyYgpSbMxCTvWWKe
G/JTZPGB5vcgtODS2dBRAmfL/VqLpBzcw8dBh5EQbg2mbOl7D4k2radcD3H5KFr1
MeIqItcsnN/F3VlmRPTo5y/bOKC1KEDUotgooB1eo7pEXT/nt8oGf8/PWtyg+1bm
V+vVnnGbTWs/TJG2itUgldCl419o2H6y2j5w/UjNTDg/HboxeeXIC3WFfRfRBRkI
BOMV04//0ZBBPYjSc4Qq4SgQ3EoKe7Z4H9G9Pog19wrDqA5fV+5ZdgH7+eJMBCCr
C/zIHBzS9kB3Aksw58uiRqtV6H78mAclBpmqtrQSBfpYAl29SFxNpCq03iRGvs8K
QKHfzMaMXi/gNfU5FXH/tgi09cjhlFYR6wYEbeSQ9mP4LkXOlbPB/XtQtxupbylh
m0BZZ0yjjpl029rvNNscbo6k+A8r96NlIRx3XYWyTfgoIijAAaZxSteMUtNHeOzQ
j1BEF1GlGNlN1RXZ8PNYrno4uFytghEffluhcmsPpKDnJ6QNgkX5O4Etmz1KKTVr
Ksg44jORC8rs2Aco+r0TM/FtgmRigZN8EUHIH10McQkR9qg6ZJz9ddMn78XLu1Ob
75Ve8ks6/6SonOOCsklfRjSKSsZmKQfKS3wZv1avY2mln+NUwNVtiCCH0MdJbK+O
cQbk2kdBPz+Zqw6wpQwuz9nI6//Wg994b+RChGEkl9tP3TufWZtFN5775HMsJwSp
lBE6y5pOBJdPTp0HngKjcfRtb/5qwChgQ6PJxCojyPPgFNWtKsNftBXrF2BwKJO3
92+8p4bvAX88XfMmmNiMhMYGdoU6f5IUfMAHwA9PHWWDv3kACfoKmwoZ0oBTszyE
uZyyNsHUVrY12n/jiq0rChrWfvxrCOM3USjM8uzKfR74EJ0bpsgwuusSiImwxwcJ
eNPNGgXTXPF9/CJZ6GL+eeUeDfp2mEN5J0uECswXn541cwzCULvlTGa1liJro6MG
agb1UiUTbhYxzuMEFPdoFgE0c8iGAwxY5KT7ztg4OF3+oBUp/dTSXSZn/iVebY2i
Uej6PFUhhJ0fowXHO3NcrUb2O62Wc7U/VWkxCWnN7uWi7XSmpLA0Y+TjZAbdb9uO
rmuKGE523PTwIeI93ycleL+qV/Jgw1JMeABpfwVdrBVh9jDF/bvTlAVmN1Gz3riJ
9gOrr3ECjwJL/0XWd/okJ7WM+lecAD62f7M/sjKXBaYNG/a+GbAvjkkQCVvmgzqk
JjNvfag8WF7ASDASKqsQ9kwrcqWDty2rZVi9qT9PavygY+p+gvauIZJJJAd3R9/A
Bhx25yfsYCbTnCWoHb01vUT/y5DY8oLwprMQkEQtUM2fJNOXDY3W6RII0RnuMPvD
nSLrbXKUQVPM4Fhc6XICpNyRs9QGuT9LPjAWN0dVV/TFpGFmkUmKE63KEP8kU20/
iFTZOnQmMcoGxhpcU0VrYE9aAFHZHeAA3k+BRZP8hbLU/qi/9ea/LKvpnGGkf/8s
9mecEeTDZ6LXxRKEKt2rCIx0v235Pl0Nf1/feD4TqyuQX5o9uLrLSKULRRx6GDT+
sv+p2AtuauXUwALMSPNLRSOUeEP5qd1Cx4osyUPOzX9OqxyEJBfrMVCDZYiIsCFq
ne4xNzuBKP/f2zEhofBo8VVnpzNiVw/jMfGFEbptRUUYTujD7czkzewSnDpmrvxr
nT3BhNHbyCJgmd/77BK+AGdqLCGjt9PNB2ZQfYYrNMOXtQRMkhw5iHSk7YOKlfRz
XHipCvghh0NRVizH01ye3+T6iufOiA6Dcxqr2+GNZiZ0khJ7jv+A3YLTdu1Ciopt
nTCTz5BMo41W5tcKLA5sSJSuaV9pJLLHhuKONrp2gG2kIdym//mrx8M5jwyfy+C8
KqnWmGeMBV6juMP3PHAQZpWbzPiv5zGi//vwVcIozjpFae9n9arrZEwOslj74WbX
dMx9mSF5hGln9CYz8HDNYHo/xsgmFbGvt/iNB3NWeuMjsO9zQa7amSIhZUkI+nFa
i8idl7LE6j9wLKRXvgyK3BfbbuA5xBOOWFGM4M6CTMNCSlYu/qn2Q4k/rgm2DIWw
iGCf6zTYqgLeweU9dWa+Xv8+z/uHpyjf5K0yqD3v34g3mZeTjzY/AfzQZQ8o3rs9
HWyFoj+MVB9SOh4TMzrfDvVCFJY/W4t7Muus2m+gl++SviSBJo1InZXtZ9jrw8jK
QGjXQqRl9HuAYDMTMgtbppvBAcT3xZBA9DSAiM1awA/ALaZ2z0xoSZb6/VzI1qpH
st9GxIKadF/dtdk0FT/YYwUUlhNRrdeE5sx1+cIkPwIH6xHPUsCGq43IkMU6m89O
OM+pxlaFlbPB4H6hAiBFSU4+tza2tvk/QITZzU2Uty0PXHOkzbQgeTM7fd2eTTAn
eeDG0fL1woJvm3m77tYCee+AnVOBRroXQGqeaqTVzBXMM5CNG1ethpOiHZCd1+R0
HLXZ1zsEImXrBvV0d9jNStmbUriwoLEcNdvFD88r/twQ9v3kR1oJPpfdw/weTPoV
XbGb4D+azshAK09Kkqj9OIod9Tj6837oAscAbn0k3PTx0xtIs57W6rnHllA362Zc
spemr+lXyqKJb52l1nh1vhB9HQ+fIhoVbUaLn1haaADMP03XmfDzNJH0B+slE8xG
t34Hb6siTrSV5lYb09Une8bpF2lPiT+FB78VFpGpVSChDrI/9Ql0aOr2hUS3b7zI
P4TzFNnFWksZopyA006hHVfJfS/qqsEVooVMen+aMmWLKJ/vYRV8usSWSxxcQTIR
Vv1uIUmPXar0zlecmepTNO4C/KxD9BdVJwovQwF4BcsAO4QlmmZkioCVzkEedA9o
rpHeU5OLjA/9edI6qLCMHUJ0nmCSq5wNL3Nk8+oZO5MFYN+JaIrqvB3usb/46Ob5
JxdraKjTR3GRGauT7va7bXPYpDTZFWnmo+b+nB23KYgUS0a5nKRKzLLfPesPd+4G
Gm9YI5lBpiHkDkwCPj6Bh61Hr/Y3J1209UJVByZO/1880CFJsgYqiCjTFyowIO0k
ZguCbdDgxEn65oEavzNiG2XuG6JGKtgeI3NIn/f8lecLQrfBIdM4nPg03fM4T5ab
t6p05x6cJwRNyqsjx97duVTqjLyMy5xDiGyJa4sXlKHotrL41PjP3BnKR1lT5bq+
AcwHjjvc8F5u4ehSuDD1LoHc34brSY8+KgRqxSIwfchNsF6G/IZv+fXcFvnBfMGR
EcTr6Jk7Y79uF42n8EeVbd2GwarwdumjdG9zYDvbi/q8JNcxn9RKIvw62SN5Oehk
m4JexlDk9sAdoHC7NfWrRE5kJToG8oaDqqq3uTL4kOpE+yZDNGREWKHHUcv7phIt
+uhjqbKcTZvH0D3xG+l68qh8+C+Xw8hLsK7fsLXRt0j/sQQrrATNwxI07xpzOkv6
nptV1yAmRtk/k1pKqk+Pq108VpYFnz84zGOTD0viouWak5XHssA8+l2SFs5fxJy6
KNrrgd3wXTVewKeP0aUIheIbSjFStthWVIsjWZzbqKFn3QIUIwedEFkA4U3GmfOb
5EizTWVXdOFNzNc7OiRc9yct2vDoMcXK3Nn1aaJa42ST5Xw/Wd/G97NxJwhDleWx
ydw9AKyX7CkktR4GyZ5oekzfdIQhRE/Y7w0MMyKjgpMVzTWY7fHswwc7OEVucG/T
xs0C98PseAWyR4V4D8pjWlBoWQ0v/5fM4VZHnRHbFkgDjYG+cU0p26wxwZXRoQyc
uLyFscWjnG/nb58Af/xWVzUJ80BklhG2xP0yCD5Y+YRvg+gMvyqpwkeRb2ZNXBL3
2s5Ra+gze3SY2p8hibsIA4YgcbCSk9zv00gg4powjIg0hUIkRK2CXeHgOvtOeK3J
CnWdawQLqxDInu1+hU45/vJBC0CDd7MS6it/MJFypdRgtlkSAVg5MQPkQ9kXbtTh
eclJOc3zpGgkhYrBXD8L52YvfMxemqduvYsojE7V7uN5WXnoe71L+8zzFxikMNej
W3/bINHWSfQRPuagBvyoXTloQB3dRBymPvf1pf/zydbJN3Q3lc/zNNypxOkg0lrR
x870x2arDAZSMJUPP9R3BXhjqtxrrrHi/+nnPR2lcXxuYixsVokFpumji7eEJMru
+rSYyL2VTH0zmgxtcP7GNr5kgnq/GAdipBwVRlOTbDWaHgnUqUs71ndNbR6tNBcI
sOS5hH02UvtJIbpqonEN0mXfSR0Sl4603iznmeVWRlcU5BP8reMb9baoAU5olLb2
RZH4ZmxzsiZHz6EhQUimdEV19En6be0oVoyskUuv7nvC/wiemsOdweZOh7IsPyWl
iWJJMaXbLb+FkWng1bwGineswLLHAD3Uc/57uvi/2vR4SCKZSafB5VErk4GVyAa1
S8xmXgZR9ymIBZrg73P5Ehgqkw4OcWNj90J0MfvXKLTJgU0J47M/vntEpPyeaJNn
8z3mFnp5YrEWB9WkdpjdHKSerTC5mrWVNOeMtFEmOo0XNDzCY7pOG/K6iEh/tMp6
VGwICFOGq7yVzlxa1wNuRSLW9wmyLYy0lKkyiLBYbGMBaoGjv0x034XCYaJiAl2E
jfAvreHz7fIjxvnaMwzB6W3h/3sEj3AGalju6xl6c8SRAOu13IPShnp675K+JiSx
ENFgllkCYzwxVee3PGPJp5Riv9UJW4L42P1JO89DnXyQhBgNY6CPy7x2BFBNtVVZ
WixIC8XMyIcCNxk0NhALsTAYAztkSemrLUytIJejl2uvGmdFTCmLVm4TbNBoas1Y
LYntX+GPEs06ZiMtwMe0hnXNuPIY40RvijxwdadT63d9MRiCY7WmdjTsNf6GKvdX
qfM/6l52CS3Ntb/iHiHs97mBKaLIMMh/XUWHlRqX9N/8deChBzrfsv0SUJajD5Qe
QYkbjnw81PKx+d4O391mZvdvhLsexbEMW75Ysg/3HW9sys/gqtRQfIH4C9Vtu9XZ
Tg1682t7sC9OFkCHoBq5k46h6rbFMYZADqRkie01xVqcEw+dIj7HNzFnNx8WUzh5
8WRKkEVxF5AWJaGMyHt48Uyip+lmyw2qlSoMfuaqs6ycuPc3d/Tx0CTlFdqHL6Bl
zc/DQfOaHnWz/H1gzPR1pPAS1wgoQ0wI9/6+OOkTkW24FqkS0Z7+dB17cVlkQklY
dSEI8PtMgF01J19+ovbsgV1kyMCsR+MFS6P+VPmHZ66Vk3wsI0m0Q76rPOQB2MG5
p6aqND/Xptzq7xrNl3ld6XagvYcO9R3NbV1a9k91sAnpI13C2zz9uB7SM5ZgDM9x
xXQ2RvO44qctxs2A/n1IJNDk9jSrCxcP+dqSk2mTXqbHFhYCQwDsMIx05KvaCBGX
xmEbjRxCDl6Y9xJUx+06INwQCTU8fwkJ+L9KBviT4hg/RBflF3u1a7HKZdY1w369
2n8rVVwJOdgN26w2/VhLl2bjgBXJAmWH2YtGU+KjZ6GBa9KoKHsdZ3xcUxigCor9
PI9Jnv+ZoPWbemSaVw//tKaP9xUBavIuPWKI4jjDt3K1PILR4uojNifdYWkBGU+q
vDF1d6+zpSpqsAdjmp9WWrKCuaYrkBqO69EyWoyDkkvgjeM/PJHLtsYLFsH7FczF
4+qY9kR/6iEhIc6sORSU5wu5d5aP9m06NzxbuDwTTJKlXagGZlKs4wh7B+EwPF93
wuDZ1XVZtMe9ZWjEex3TxYzLw/Yy9WU375LrpIHAandlUKovw/oeC+TpvBnKBvRr
ge235rqRVCqrD4VH5lwppfKeBanjbCJPz9SmlOxO91M5tsAMuHkGZzJNqXV8tw3h
+Dapk/AgDSXoz8JxWDRh4BTnMeo0qwbj9mW9Z98JrSXXmpRPb8u9N+yg0QRWnDCR
cT784oq/DlYsAGKWirNfG6Yiv1zNy+4060QPJkPQrsY/sg0jV1QFh1H5sPeoEh6s
+yjBuzC49Bn+LtieAljwBO/jOJ6/f8QWXAEunGWtCJYfZuPWwzCzKxbm6CiPFkJn
3fW1SLFhrvv9A+N43Zx+wDDKPwKU8H1WYZeI5+qYp810ijMfBFNE7xfO+nYdzJuk
A9e4WV1hzwm7NwZSOAd1YRJRy9P/uB7lKXAsLkcw5hU8mWzhpQ2y6zeA1RLHwPEK
ZEH8Zxezp7JqoXy1S9VBBkrY9impElVdYC9QxoA9FHMqvXWmHYHV1h+dD01txiIp
n2PoJdm5SaCv8P15V3lFk7lXes4DUwW3DZ2A4QLIOWVdGZz/isHJlixb286UlgWT
1l3ZiftbM5Eu9sGiKD7hd7r4UV8wG7KFTmk8JM7ULFlv1HrHtQ44ufCVciEnt5iO
odoBke0N9kYWjHwRsBnSAKO4Q6LSyIpKlJZvoBHm+LOvVf2LVBW6xiCIKBTT+lBM
Fyfi4HquFxNkGXRDOIKH7S07/M9zDk+ALojW1gG4wWV56fKnDUiPRcyCwvQUBYD0
+K36Fs53+6Z2ZbxTRtmbjs92vjMN54U52tqt7yXg1tCYUtk84a+VLQJsoRUTVVg6
sEGjK75GP8cGoo6bjxBWNbYW/ACd7VwzWahzI9t26BVP8g0FDL+d1WP+y30eDeor
GKMNFYQWFF75BQKl2mBZ6dbEtE0X0eb97zVyGVFETEz2bMXllexa9DxlH0WjkTy4
AB3kPRPzCdYxtBjTBcNx7Z6V1MEUI3e9hMd2zkYOfl1BlPUdcR4im6o36EFuVLlv
8/9T2D9MLSZv8qtyHRL+mL03iwbSC7eHvP/Fhed9cOO1m6u/rqsFBlbu5QhXZWm8
nP++t9oNqwCGiP7VE+z9ByFOZj9B0whb7uiwZuQ9YcfbsHvG1JZEm18TCOKTnmtl
ovTOseWxs7f4TDFnLiIIEdjLfD99K80JM/Wn00g8BtALjtLZSU7qpAp07b8PQUx0
ilRFhiEDRsSr2RZF6/91tZ85W4eHbb5oD+q7E+3gpBbPySgCKppIkV5ErbR/JbWq
kl+bQ16s9fLVPMmjJx7IgHJCrV1IqXwBW1340xEp9qAp5z/7CZUvOHfe7yfThDtZ
Vs4O4RvgOdtpu+ybm4t3Xqs6/Ux9pMUswdNjcXWQrQYx6vVrHSj381j22tU0SmWz
ty1z+PLF3HvH9cgrHrriZSOGPjGFRZcr9AULjvebcNGf9SEq9E6me7pETePmPEkM
jLh1Woo4JyXd18v4BlTOydiKlg5XwYHKQQDHrZseIExgWsSjakZFxhQHz+EGJ6je
qWxHXuorbdn8wRNCuPyoOtyPEy58tvtc7I2ODOigXuoKd2i1q4L1DdEnHbjJErrP
Dly7SKwpYumP5U3fQmIgpnngKW47OkR5G4texAgQtTtQFC0uu+PnoQxfqWeGnRlV
K3EKYJphqf5+QHWu6Hr0N/t+LmNl3+lsdxTK1l7RsYZVTFcOBDqqozgTn82vIFiS
ry09HSPhIPdixBQ6OhBdklN/vDJ2dWNJCtsJvPuf+L9KeKNP0sRvtm+VeZ4Gh5j2
j3VM4m7zTgvC5AlMIN/myjN9Gk8qi3PJLGY0R8KHtkVU4xF5BQzRTifNMKn2oTuY
w0xmXm7tQJ2pyJO4cu+kIrAghGelOcuDHUoCToj6m8K3D/EOjov9JCAqhYV6bT4a
TQvZHZtGRyq0/mt5HXZdw9/qNG/A3i1krbXeXLzdETrRN8p2r8CvrBU898MW0ZUY
PqgNAkFPvO0pn8XYchVtv4LDb4lE23YPULOR+A9necS/fRlc01z58UXnveKGVAFh
bSchZ05uEFX++PrIadyykDBKO7KNYzTyQY3htTxHELkR3QIbrF76CUCJrMe3cdln
lt6F2b4jz4c2fqvg4Iq03sldIir5n+sOhgHaug4l5z938fdjSZzQ2O1W5QhQIj1N
y1bL/jweDcWBLo7Xg6r5zggPioxekIB5rQegXNszxZnk4wh4xkKF0FbXXjVtIbEU
XNQFwfV6JYlQCg6cy7XoJVOQ7RgpaJ2MjgBXREMWjlB2jWJEeAKu2vYRJShEj0eT
bJNtnigpCAsUZsxVPKSyZP5jDSObdA/WV6MATwgly5XqQT0RZOgQ7Pb0a2yzkwb8
cv7vTGbZY1APt9PjgqpQe+d4bMQAy5KHkdXbdrIHJG4Bln5Khe30u4XqnpjBZSnV
5tT04SZWgXKu0kguxcl5XHPinI+h0k2/TAh+jtncNw5Xyil8XtnEFkbG06Jbo4e+
v0pTNo7weP1ijTz1NxLJk58c//iqR1sSd9oAvxe4A1oPF9CaTp6EDFecaPkSV5X3
6okD/1E8EoV/6DXwancgnx629sD0wVbIursmeQZlWmyiKXLnjR8hSoTUU1QwOQat
0C01HIqbLNJ+z2ByonktHK9iJVJMHqsxDNs2j6QVnT/AlT3eHlmVelQNY3DKtXIo
K7qxW5vKQekN97Yi+9KGuyHhw9MrE0rsQ3aaGISlEBjjTdYmOjUkpIxhgcwLlcEi
qFa4NWKK5T0oam4DgEgZy7P3HDyLfzJLtns0RO8rUrlecnv/SDeVLn7UxKBMNxAZ
zQjifJjp2d+tMC+BZ1iqeUGwJjqLggH31NjKso/QxdxszVqAvQUkQx1PNUBAF8fv
uSuCyciLDfMa6cALvMxJ60O91SCSdl/G2jcBZ4yVVrGI+QxtIU6HXCro66eLcA+W
CYn7FaVmpTzwjdzfo1nwOp6U5AyUxuSGqvB8TDZISntwhelBqoX1VSvoVxclZOLi
j2gKd1WQYjOcmvFZb/tHTLUAQCn9yL1sUSlUNoJOSq6GwVmTt9/yLHXemSfrwZsI
1Iq/NTcpJhirjw4ZzbRjfNMx5c40pMiVHLnFM1yJc2lovcMpDrZPrMivtrec+1CT
YV/l6mYKBPLKHwnmquq0LJxzvwFqqoVi/6nbNknyTQnJHQFtO/5yrb3bHjh+e8HV
njl4AIDw13bp02qeEdvvjj9OJcbkQTHmIWodzgQqn2T9rnevJtNI0roXSMe91tZd
K/GS1sZC1TKoUOgaEtTm22IHbtc1N3kjHFPRp5cA7/l2z7OfrIhlH0nAN3nAwgCi
ee6xMZ2KjCoDSMKqY5LOOu8ZA1txwNsKJDyaY48SQ5PWyAM1033daRTLMYiJOeub
lRabaSewRcgTI4nVkR5E3vxK+RBN9MTbJCDb/+ECXqjFHoq2btaJ2UCOlZ8uoKKo
dPmN1urDN172eLvrD6PuhQ3EgBtdlQ0fAGs+I5hh8nNJNdWGM+W9cRJElT7et+ZG
sOTzfIambsQoqc9ispmVfXhRKvvrP1PK5ymEvvIuddiAjV7ZxsC0MIRo+SioXExr
vvR7FFvwkBlMYHXr98LH27UpWgqUDr8mOPiSPZ9Le9kw7fXbIiIRr49adn/zGede
cB964+rP2SSmw5Dhfeq8VkYb9xCxyagNeBvgMSnNpDF2CNBvkh/s8s/pRWbbBLqR
KiQnqCVTOrJgFWeOE9ch18hawi07V7/5krKMRKsYv2xDWGgRKn0ZJpoVxePm4LYb
1o8cf6KV/Bo7vtB2uX6ZD9+na2c22miT6oA5P8vLHmdIN/MLrjor65U8ODW507Iy
2njaibZtCVZvYpm81zonHC2pz/WrHVSIOlGwHjdGSFJywtRLw5JuKyqq3mKqN9Eu
aDy4FUSZ8SO86Hx1DIP2IrytoBGgUWBngx7cxwpc3r/hTInKhJwgRHOd+VujJpmI
q4uwpAx8gGn2nNUuREGUY9WKhLeCu6OeM1Jx21c1APERPVKQKNn8lkU/dJX4zK1t
7fKa5mv12d+eEVmjqMaNbuIEdlpbKVFpYvavoo0Se6Pfwarxk1HQ/lckzh3lWkMe
EDK933Dbgp53nErjG34UXjyBLSy3Usbtuvim14KLCOhKKTx5neLi6Q0NFJx+BZxx
cWVn29yvAnLXmCS3YBCWrC+eo5yKAOsnFa50mcykQYgg6qHu1XFnLmwD9k1ZuNdp
qBbLIRZMDTnNyZj2ao1v5bVoicpEvh2KnpZjWZRFkQl3eNrzWko/Fa2Hz40fezl1
gZPm3B4Ix8wCpMgKdJrfmoG+go5Nir2d8ykvADEjh9wbWZgoPpTtOwsS3ygn+hNS
l2YicUoCOc8CedicApxZhvwbAEpE3p3SZ23PvFSQuwtmxB6ZwFURBtgqo4aBpKPO
NrkyeTeDV2iQl9O/BtDJgXUKLEBNXvD8+rhK2u29qepILQpLuTa3NfL2pDwriw/Z
Pw1vrXgh+aMqrrRmhnl56NWNqZUx854IxpMnIBciOD81+lePUjBSqxo0/Ha7cHY9
nXDiDUFbayh3U0T3A08FuPyjytanmUYy51FTf550/wzY7+BAXROOVvR9kRMyFlC+
Y/UQp0cmLoJhs1lS0YjTIvm2guJIEmmpk0Zb9o1PZo8wXohEsE/DWggvk/PsUjmf
YDVRWCeITnQoXfiR/f7OKrv6Wj9Rto48U/vmlnLD1QW5x+BaJkAeJv3UOP56ckjU
UIbAQTGxW51FnKYnO7mXxjru+bRjjw6XMXvPbcV2xYzzAu/MG94p960j1dCq/3tU
ACCVY9YJdF5ZbWGDWUe16pJ+/25E4dz9oymTlMKvRv/YbQ2EK/CYTvwnJqhxo39C
tkgVquMSCrwtM1wOWKwwqMHJZnxjFsZMHp4KBwdLhjvOVoce8/CJqossYC1HGjIO
7rNZfZkypCS3Aw9zlj16uWSclfGhlPRW7e1uYVR8jW9DLwRV8yYzumGbRcGH3WLy
8Qv5UloZZXaNRDN48O2wTWYt/vhMX1gf3eVZdqILrPtI8qKadyNlAVSWebl4+0ge
dc9LkHmtJhx8TodHDMCBtWcuDvEdSNW1mygM8VhTP1IW8xC/wWtlLWBvq52120ms
w0gHRkllNSIdigHjs/q4hWaS+z6vJMfBM5+BqP9ltIOrBln8hwjAp+vAInq/N1u4
H6LtigPQ99BTW9kT/Oh3H00DKZvTbHI7A3FMidYA7mReDU+vv+VtFZJjYOT5V1dd
pbXEd8IM8fcF8JK49/4XjfR2z+zQ8NdYuYAm1lneHmljiXwq6XacaRUBJqoX5U3/
Jvi5Ch8PxRteG1v6q5x2J1F+ILsgsaKeeJ+yVF1Xj36C5QsgIPEr2Ae2hsS3n2rS
RomT21zAWg1xw6N2W9Xz5tokCxtBfdt/ntlAM5L3VlhP4n8qnMhIzBMGEqFOQnWQ
9OKqDrr7c9qwAnMzJpYRbIOuoLlTbMWMCuJzXDSWL+GDHlpZ2D9VpWAbfcrHCP2D
JXUFDc2Jb8PucIgffS/POvRGUbEa81Jz/G8yN/wFW1deL+ti8Ii+aH8+EpIL+LdZ
BJhyNN7tmMf5WA/2lWuDZE77VfwJS0B9cnAhCZLv8F2DCzmAl7IDKBYAnmoQJF+v
OD7FbaPUnehpNu8Qkk8T6n0aNVUbxV0JlU/XQnkoxVwUM0zhKoxNCb1OKLYTggjB
8Qvba8qvsvPbWG1VA2aj+x7YoxdeJL16400qljDpeTGc/Hy3yzVXP1cfKRji6Dec
HxKIwJtdaqyBe1BctbipLmpvDivNEB2nzrF31ow+m/CuV/YZsg9c2FNy6T3cLX9v
yVDb/ASmiqWS0vi7J45AYpOwNSmXgjTt40vXe6l1zZHnaeP+bAEu6DdInQK8Z2k7
Utusl3m28Ast0fj4ItrTIcM5er7HZo6Szo+wBj/uv31OMYR4oY4X9GfE9qDfspVC
d49qizbSIIpP+y5qiX/bo9aUQpYEUjLpYVLA7Eo5bvyMM9ZTYfjaI89oeVL+qsuk
optCtCKf05m5ijxeqZxDXzexinkYJEYtZL+Kq+KOVDcsTBGOBsJBuTLdtzkR189Y
pneB6DQtNMB4JGWaaeQXcdnpD0fNlynpFIYvhxDyW77H1FTxMWvYoVC+RhHibTEK
7vm78Ujf4IaDRv595QpGPZaH6effIiB+k73ex7vF4yuwVluPu03N+AM7fXolCriu
rSZJk2UGlPfzAJKRapgZxMtGOVbg87y029kRh9KmuSM3ewRSpaGp+7oHQCRYIGo6
ucQJ8vaWS1vk2brNQjIWRzWDkwaKhdMkokdRkjzsjoKiXSiR+7HX4D30qkhPcv0Z
PrDVjbsgXpzy7YHvQvYa6BdoAb/F/ue73PwzpUeruYUOGIONJiaJyGzV2xVdKG40
oDHxZHoXFBaBiN/16SzNeyZpXoL55azul2fiIf4KQNwQXxaVs2mTRyxpL65LvjV7
zb0KDp/H+9rltui9FZ2S9L1b1LYDvlt3pDjWgv5lfO3LqpJb4Nc+88wWWAT7Co6p
67xDv0BCmRWXp4fN8bZOqhDFOn12myY7YN2M0vaBbOGEjaVA/WLnbPFpghrEd1yC
CHI/rdwkrKxmKnUg0ua7xR5GV/DYEPH2SMMNP+zeMBpN2Yc2PLq7Mg9CCAloFCS0
qh8NXUCA5qcMzq3e43WYyK9VV0vufsGBtWjZ3Yh8pC21zT6D4DzwZbaiFpfk1xDz
E0qL3JpsYAonfaLD4GY9gFR2FP4HgtJQZRZ3B1BE82jldYyIJowEybGL85UOH5sf
t28hFlRNF4kAB4uSvAiRiwvFpRrCNCz5gboAOguajXHAWp1Rwc0GaYdEzH0TD88k
Hma6xUuCzSK3Kht6dbsHyKXtXlRHsVR6Wt6kjKlJ/tZCh7At8QzZJHaHGxiGkeMw
8o9GOj8C1OAcuo032MFZ2g==
`pragma protect end_protected
