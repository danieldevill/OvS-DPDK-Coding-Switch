// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:34:47 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kSpiff7LE+e49oDqGEbFCNc0PcSiQwR7aLGRi408FVmv3WBdCIVC9uJ0SmMwDwKU
EmdXWiHJrXWziYgBhE8y5iEnFCQrqVjmKFg9s5AK3i1VrwnjtjBBhs2mtuybQ9Fn
1Ve6QpdtyFn96E7zdnk5HJEcyPkWU2YzWNuJXSXT324=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21904)
lcnqwVuDteiqzlDBQ5oXAB6Wwz1s/jt2ixBmncN1ihYkktLHq4Ch1Y0xSM7wLeBu
VcRtNQy8CC2kgpKTCHDlQgtSLuUvvcViBlX9BICxUNjTMmAk5OrEDG2q8YlLuHUw
9bHgtyJi2h/dDs/qhse8xrePJeSeKbxDPfErIFXVMuAVBWBbjp2/mdWXve7VbgIZ
4vuJJbmQY33/G24jIvzWcwZxQIhzPedFrsgXapETKDY6KK6rzPD81bB8qY3fchv+
KUYok20N5VN2tAHZ3F/muzeXGZ9szbtvYldA88sDxNLXjf84AZLZpm1APKG9G4/e
yZI68aGr+l7BWkTyZs12Ezh8gfq+WBulrvUxEfuCcHhRv/JWbV8OoPETks6DzzNo
GllWr/XhyAUL/xtPO10ZaCYoLz57EoxjSfMJ+eDRID3lgE+39qm6ioDXyOs6m+sR
gfoRiBEkWmI8zL5bUWZiq+Mt8koF/ckbhb36k0b48x9SStgnYenPr3bVjVCWkpEs
+319Bz2VEUQtIRa8L1qmYJgHY3sIP0lRz/FrSP83GMz34EZnLz4tUWSGB5cCsj3A
0cK64CMZ5Y87PSMaTjOmYVymIHAuXM8m37kYOP55jjB0Td4KTFhzf26Wqkzter+4
myy9/JBtT5+GxMxqC1TZLaw23n6m38jmrnA7pBj3Bgo/PENj1Tu+ouAbjk6HOXJ2
605sBxc2+CNWFh9+1PqHpZ5uJ3wAHRzJ9gz29RZDdLm0CTAsAlXTe+8y1KoKx2Le
HkU52ZzgJoCR6tLGq0du2ivLdBSbXgLwD5TXoNlD3/QxUQwHI1M9kLz780L4+2Yk
Q0QVVq9GdJdTVjozlpUxUnLw++/Rc/W3EtTk6+74F6SXywCTDaF3yFXXfvY0lyaU
GRyorQn9Bn0uOhPUnl228XLMHk0wPt7LcnRcJXEZ7MnNggFa4JXlmcg79C4PfNYu
RNi3GO/iSIXQNlQONKKIXIE9UdI0JYD3g3LdvhwbOa4H2zZdoB5OOC2e/QweYCtg
NX/Y+yovHaJWExEEQGemrHfjTAPA8vYWSbjW5UCba2cNnBNf8/ruZ7MH26byxDTz
n9zFGNU4l7YgXwYvrzAecUvOdl61VYZsn4u2OeSm8Ok+hQc98xIxuB+EY08fPQZg
Kz1YN7FCLjUpYAY6fTUisRwx4BfZ+0K8Ti89K91IwBHzHDS9l5Opljb1IRhONEud
m1PShWOQqB2lLlXvcUZ2e5HGY/5GfZ0WmccpbZhOtZb1Uqx8kYZQ2CUEtfIQqOAb
i+kA4DEtyiQuqdCsxCMCJsWDTHvpim7Kbi6k1O+Z0iFBd6lu6Swk+kSK6BxZBuS5
LKHjYCaYNMehprvxG3ikZWOKTJj5tx6n7Ay9OhvrqFmNUR5/QmkOqXr+Fqvlx5/Z
+tM7nThNx5Jo+Y+YP6jgDltWu6j+wWQMFLqHIpdgkvzMsH6vaWUO1z99H/E5yGjk
Y8TFzimpkLafeLzJvlJflSXXJPR2G6PWLIOLxFps01qZUwORaUDajARGSu0nQplx
6kFe3AFttVOApdTsmE9ygMQB/j2rM/JzR42Ho7BDu5t5U4tCkVweN6FuCpipBCaQ
QBOPDwpjioy4jJ0Q8QIZyKMU1WHkaKd+HhE/XOx6Iua60p0JyHDmoQeJpwbCP+A0
m909Z2L+cWjZHXmtPjP32C8Rq9gGoxzi+5O1Hc3nfDEH62LV/GjsQVWzfSsTjHgH
32jZ5Ou0mR5QG0VxAbGISdg9zeKUZHwZjC5r4+aAuRxTBcoSi790NjGhU6kim0kC
+hzW5TccGrTW4L4ijrFU4S+hq765+WNKS8XbmC7IBAMtaCjaZsnONeJbDv/PHd40
6wJnJx2SMEeNa1vx14AW6R3UBierVXTuVNRrfnymDE2ybF7Dc3gD/TWt1tYDIz/4
UH+VB7icNNU+Yqf8Q6UcyyfV+c5ISeZSvaSX5o4PXhE5qlMxldNKGRCw8oRI9zXZ
wesW+Kxswkal4XhOiQJ1bQbMU2b6RNCvXQoSJGPKA2pjPKMUBTna4wqPFl7SCu1G
mRhxPEPxBYH4JnnojxcBNUI+MiqRnX8FSecijrijSrkHwMw061adTQkOOpNNwgjW
EEuz7bojqFw09OwP/mkb+NDrmiLHvXIpP8ryqeqDDQNhX6hQu5MUk7cUfhcykdKN
vfw7w2qUQZNC4pj3K6Czh1iGYvFkzvNvZohPdxhjvcNP7XqeITBh41EdeuDPu/e1
fKK5IJHhorODCXofLsZdPzJpsIDWaxRC1Qx2ek0lfy0WU57PXo2K4r/yUNFSaYj9
Nm9OBUVqD7jMq/bDhgOTb9lLmRo9UQzX8WE7IYQC1AVELlxFUl1H2RA2fYeBOBc3
trhEg4seDt1+9mtkZ0x3ezo+WORMlWd1ZWvabsCTZQwxyjHx39OlL573YzLOwLSq
CgJ7j1ninl708bb1zcd6HYEI1SI49oP2QdubGqnZP9w8PLATXZ64zIUzScOEO0py
IJ12+mj80XfuMJ6VRig+Zz6fKYrlzIA1FoNA6ZRkJM7VHpO4WdaWwXGlTNO9LNTQ
xjIOwfByggUe4GUeI47K6m2kdGydURmREyhRpbdKmyeUytaukJ6YZJzniV1/O7nr
KSKAoTZR88qTYUXOCRAKLAf15AVeNFj9+0rSpk92PW+nfzUR0EvPiEESo7SWr4pL
Eqm/ss1SV3Hh3phOUvAQEUM+MvLY7UYP2+ECw++xx2P4Gi4lL0p7ojYSAssZOYJ3
d8L+E0pT8b4rWTZoYkiN55parN1XpdgkKwuZQG1R669y+CcbteOEgoVVBFhicHqs
n3gXgFVo2oQ20qR23EjKC5pS/jzcoXjWmPI8WmvFWjgJ3XgTpZ8kpEsUeK5VXWip
s0ARbVfYKr7tBARbr5ONiQjAbGdWseI8HbyxqqsG05g8yCGDV+N8NDLGUGDT2x/c
cfp36M/lJMDa4SrNxi1+TPzx8USh99kUUIBlHerdOKKKnoYL0ytN7KNABEtxhwzQ
kD4AgZQqhFK4zmJrh2H0LEu2sozz6+ItAJmFHhj4AiHUqTGThU7TPCpsN21zhQBj
GrML4xRX8v2FUwfGIsGFKO1T6ilMMBPShvC8YXnMnQzbLpMxCFFYo7svZ37yCb/V
l4F7by0XDwum+7ALN2ZVK9XW4+CFjHrz5526eAP2/qJNs2fbLfNnn9i6gsvdFWbs
hjhntjEdussiDWdJw0MshtgxV6+4+cVJrofUZgH7lFrewYGzwxQCBRvWk7DSEgJg
Apf1w/0tMJCmXbVjLB7xqglRUeHqUonj/T0Pb1/Z0W/KCpfmgap29IAIkSEJYSWj
6GbismFUvJu0FgMuWALjfzW+E3YG+HIbSPZ+07QJVEGr1Cv8ncnIITOJO5vQNFk8
N6k4K7ryUulVRt6JI+olR2QWK3p21is5/wkvSF2WoSmXePjdTBDwhGtQeNw1iqTU
14bbLmWOkVECtKlckXiWhnkx5m/mvGePnVgXAZBStEVNeU+dLq5sCnJHDsRgJUKt
vazYDKp14KeUJS6wCyCOsh0IfL7KJVl5pTu73i3oGjoxV7ruXI0ySnHjX3HKSiX/
+4NFR1tm531YYBrHXqEpn99tjXDPVun8jHA58tYJQlI/uiRe2suIn9eSlT1lK6W5
On70QON5dsZ8+SbN/LLirBTwCOzO955zb/WIoSLyhX8Oq9OhsP2EAqYW4vwMEc6v
coHcrM2TKCbbL9/88w1CgHYQJd2Vtn3m96gI6v9apCzEZPrkWlgIyXwlIZF8NdBP
xC1j0PvXegJBtKi5mVDpCV2IQJPQTRUa+aIG4m/oUAZUGoGYy9RnXp9Yg/TVFOft
aGBAND7VuDy4yNH4R397GNpxbjLNZ1ZMVoMsBQFtFlxKjTUH4q4Qp94A8CSeluLT
bFtDCTVljD3vlXmDHs2xSH/169mWXgI+h2nlAhd9Eki0+Ond54ookiKquwGa0Cks
L/B3hzNC8wDeeaqgd/N9ha2fpLvkD33wfiNlWwcmkoJi9KnPzWQMdCiFBtE2o7GC
PfRV+JVdbLJef4uoBcyHFI7NGRXGNVUjXs2lhiHqm9DEOp158cB+9ooGj+kk9Ls6
7lxpEkJosXzT9QAFpvWnPdc2OIzWHsPdoXzVTj941PbtGNvRf7NwwtFOSHgS4ca6
F85wwOtw5EV7YL7GR6damEcaftvQjKGeFm86yDfWXhTgQRU9IB30iSJDiJR3bnWL
rBCR2E28ye/2fSiqxoi0XSdR97MgVeegFg6O8GievHsK8rjCuHFssACmIey6LU0a
1r5k2geUJP+6bGqB8GHt+feFfZVe8oW2KB4MnUvR+Yha5ReyiRbfp2nsA2kwbSR4
8xCUHXzSayUvx0GHq2SF4ktggEfozveyesoaiMyrcaUurY4/haaE3xKHhKM3XeD+
AVGtiFeyT+VLAyk1jilylYZuBnc8KNhQY9BolTzGUAgG9zEc2cmeJPOe3abEKfrz
MmKJhIAOByKvC317B1T63GnAHI268LeKiDszcEUEMJN8bXii4VCi1qV/NNFF4Fd4
1gaWRiLD8EO4JUPYRoI6vuA6AN8ylB2jWZvQ8O9VFrHq8gpvSFUYZyN6/eWNPhhG
NLfKcoMXITd80tB6x+RSnVy6tr+I44K/fAmV3+qqfnHOm+VrrDIDGzq1eGJa5mQV
XwZvUTV2JYaHg1jgv2DTvIQbys8F2LeY5ZjtitaUDx7YGc4ACwNuW84SUighC3pO
LFX+75FkQiQMh9iVfCb5yANg5HS3lapo9xHojemYI8VPYvvZ2jjtNbLDRfmfvxlV
KMumoJpc2rSi903ATKNYUK2N3UFQtXOWTG5M6x0XBdIUMnvbgbW0oCq52PHTuhES
gmmGDcG2+nSPVQh9AldOB3JaTMEB5mg/TOCwBPdBmmhUV4pGIwIb7BaVSZi0oFe5
x68tzVgDcZB+oWGpkZA7PESLLVa1YxA0kBkNJEk5EVXSnDtiMR8NtQpQHJT9B4Zh
SlSJiB4QFoMxNcJm+dcCAoUt9q/gZEgXmiOoB8u17h+hoRyJl7+YJXz+OZ+/gru6
tOEDOFqlim+MKHmn4VX05SQo8Zf6qmdDB1TCRjKTWge6mqQw9kzFZAR+j35H/VZY
kZwXv3tPaTS/WRC2TU5zUCOatD4jc2iLgnJNBXfCt5fCSucpNYBMUnIxQEC7bFA2
VkEE6xTL00mThPPG2a60daWNw+2FV2HPYBJz+pY9lULJFovK2N4NKm4z98ME/WQV
/RJZGnasmadMNiW00jsSWrc7IeWI3BbA7kl1Nx4Kk/R0pUbtlMydjRna2sGYNWAp
WMhTfOuvUk002RQLc7QCELgIa6Ac8urRIBML1BIe+1BaNPMfKYXvE8hvIlBQRDhy
aCGHy86/3MeImzTtdljM4rr931NhpT+qbbuQq7xTXIHM7MfcdVLmqQT6w8MpJlJi
kjO8D2FYtkYbFWF55YFQHUv8iNw0JtUFKpVb+I53Ao23jT3LDqGy7QxQJqR+rlfk
mOwbzrX7zfhmIuXpKpIUh7TIGyQqhz7jiGHBX9O+5iqmIemVZr0W/16epaUWy2o9
+5PzkmfEsDRSKGvrVyfS9U5hYj5jE3P+xc6FZHrFoqduHZM1s6DYJesh8KFLs+x4
n9AYUFUPdrxS1x1JisfbxQcH8PWzRT8G61KDXD5ttG29ow9dZ7KmwyFZj0zBr1o7
l46hq8jFAsCVypZ70Ekp9WLTWpuBu5Z/7RRz2VZ5FjKBNruicNJkiVtHEmwykQkO
oy3dDWtHIHI0nN/r5J3yh8wbZQx/nF2iLY5IwZYMGJeno1jvwWkDrpO1xNsEw9fo
tHMunAe517ztf484waY5XFesN92PitoVqrq0l4QXIUptSaAw42pVvTh2yf88YVgU
zZOGcPFDS05aQUphZJfvikx3kNNDmrL9nx/BbNe3bX7kycOxi1ZUtchhhlGXEPKd
6+MwC87ClKfv7lvUuz+cU6ozbvDTP5EaozvtwlVTQz8T1xzHp9+iKY9IaP28V+0M
AvnUQ5fvT1zy3FqQsnKYVCWe5Od1PvgOA7TPQaNBrejamvcZlxxAyuYDsSlqNRE1
FMseaP7ism84WCwyqmGGhKRAtA9wCA4oGKKpqkpdpct0FIf8Ii8qAwbF9QyIDZhB
L8kqeUPpo/VOzm6y1zHaIEwM6bJMDIYKpdzOk3ZyUz/KuGvFFeQK7+NMaeHdLfEj
68OQJSb3/Q/zfCaoCpD4drZeN8nYExF0VEGLDqYX9VEvOhu3ixiVwB7I4lFAvAgd
4/st13K2qdBGCsAYZTQJRnqY+d4AXdhihPbiRA3/39T3VE/e+/ka2zAhCjLCL8nR
yfgmaO+UEe6mdlrgBtpdnrnh7QTdRjKvLlUfPXYx3zMjMGV9KfU0o6S9e7qm0H/v
kB+/wVrbHD5ItdxhnTJilQjLYGOS36UThDQNw6zgYjcstXbrk2D/9OgmOhnEuc1N
fyMCBT9hrfjlOl6tU9AwREBGtazik4EDPkqXHre/P6WanMTUISLiYbJgSv1bjIbX
skI5BANQp4d2umQQCMa1txFjYmPLrCrF+Q+4TIvH//ZKFGYbHa6B+HjNuEUVXg3b
Z6UntCruYjuJi3HwraSPOpYzqlxBSVvfTMAuXacqQu11VCyUB/uM4PpRH2z+t3Ee
EcITz0bRkkouPgxgg2V7pHiYKCmXWWqc0b96Hr/6oyE2ufzAoFbgXgOjXPgRpqZu
6kltGKjCM2bEWDF9gztmXUFjq6qgaPj2Je4AscZ3fTpEhEDYQLrXsz96IG/Qp4oj
priEka1bwVHRxeLmKsWHedwma0I5svKk/rXEYL1Ht1tnnQNqihZc3FNDbGhQqVdQ
qUX9zgnFTi01D62bvCPQlKpf573IQ/yTBk1ElW5kDO346V5rXAYUD4BhwfDu3/m3
2cAkiGZfwQVpB1Z4zJi6yln1ANdGoe3s3/tDvCI8XWXIl2H2xS3Fz7Kk9lUB6D1O
+nL2MWm1sBwDWSjGR5+Qh4QGhWCbCrY8EqbFDWxC7gQKFLep3TE0JR+04Hdamze/
nbHlwubgSCNNZz7H8vhEMktiC36WRcDZE/dE2UzDeXGx3ixz3wKqAytXHz2NX3ig
J8fPQJNU9wrsVP0xB8zajKGJyaaIgDvZUWRerLcpnBT6gbszuMZS82NMC5Nwupr0
7DH8HUjMGuix13j1kZOMrgsGbxE/uLulUS32NSb9Dx5ZtCiUFLNaHdEbnmzs5YCB
V2VzNqOGc2LxfedF2EpI5RE4sdkE/lI6ZXBAdZv9oLCytPbxhi896+VWlV70Q1je
wFcf2/Bt71XOE2m1V8fy5RXYY37goLAP0/Ht9OQ/jSBDWtGV8/LQ2R3m8LIMC3sf
Dm2RWBxHNO5Ub7vlki8P7Uvm7xlKCYUIg+8B3MxOcEjyK36Uynmgy34gQT8qMKQO
Nik2f6oJyvRCHAVorcmn1GmK6Mze2OSrZF6LIR4ZJTW550ZAU500wq0h5SSSHXq/
ISakaeq+6UPbkEK837uBFWojU4JpI1YQJw6NjSw8Or4a2VnMEFso8qZPUwFmbCKq
BhVrvJoJerPXCSiS8WHUvkqLBXnCGRVsNFCAozbJP6HzPUW/q9HI/45rF+bKBEQ6
2HGnUtbGcnsK9Nodu9aXTfOblW0yOjdBNi2ena8gPJwq5HzIFLmDmJzQypO/Cj63
UAPvju58iDPilxLgwDmU+HgDpf4i08HbneIZ8Se9wIh3P7SjWZOzFeaJsMaAXKdQ
af9BsvgddqIGBsXPrYcSsTsskebsUhFKvmDS8Psu3GA38OZDWUaMOpWayTjnHQiX
GN7XcE2ZZUtgqg4CN1SKtDKV2A4tAkrDhdiTxZf7bnc+ezElKw5RAhvvejIoov+w
aPqgVq1EgwpqE0i3SsE2mKbVG3zDHEecsObWRypFcgI13rTcYnUAxqprPkzR1x9q
fi4Y1CAkgLa5kpXpzGmQFDqVNrX5nGeZ5FolmvvklClJVhHS6NI00R0im84rBPo+
zJvfwZOWWi3Rfj2Bta1PmH34Fk27QjfM4OvFqsF9lixSgGSmIoIbBi+BVJcyo7/v
XwAi2Kn7nsZzr6m91X3SnZxVfPzeDjqxI9iDKsT4xiPVPk9taL0mxGPMDOaGM5pa
fa3dcQHMxs4XdGu7eTXtY+wqkf6KLvststt2m+P//iYop8h88yBSS0/Ru++SsD4W
saLFkuNTlTm60nUztr1pU5m1HwWEGhRhAucZaZGA38OM6c5lZEkNMElGlB7ni8q1
F8/7jsphHzBP5pn1WPomTCQPF4/rDsB+hsVtf5J29wkZzM/dJcegdmnhNxYKoVfl
i8tmolQXNWz1IMcP7CR/gpiu4PV3y25dQaNn6FkJ2MiH8I0L+9ygyJ7OOls1DLGF
iIfxpAsF2Q6QvuuhRkvP2iL9xnddQ6M3fvbutgVQ7uHmdmRhfLWuNAY6I5/xn1pu
aWVw4BasFWb9zC2ms5eiet/8s800g7lG3rr8vUg+5BACe4xuYVaOQiMt4zZC2fRX
KCby1EyMe6J8nTDYeQLd3UMrIaUa7LLbfa/5OpG5QePYAUlQt4zbtpLAddDa2fWZ
dIWlYWILNpNAMA00eWxI65s40FjXNwiNkuQN5jKpEwWHKmMV/s5O5oBqYofdhGGr
lB6SdYZSS3UjbLy54QLBefrEiCeLgxO4eZ9zIYO5BwB7UziG9mhJUlC8FFvdHCMP
gQgz1Im1VK82grK10XpXD9mI7bKb+PnIvCQLIzuiahig71uX5w/0w8dT27SxcfbR
AvHwdlQbA38eWlFySf5za7QSgnm3S0oYOcpNqxrRNhz+ckIiklU3G0FRmvyNMIKr
uhmT8TuDUAPltYxh3+b20Q7jySHv4uQgH4xI1vvmNmV1gX6v2Aatld81nog4eE/u
aZWg104WcGl+KmcoLzXhPTL9Y1h2alfj2ZZrTK2gNi+4KF0/ymMQJmtuA1D8A9XJ
q9nDLaqVlRpGyEHugGGWsYqnSDz6L3U78btQj9LaDOqWzxKxsA9YRbcemdom2feS
B8I8trGsBLVH/QiWDThCBTAOd2KVqIDPVXKuYQaCOn6O6JIwif1n0SJ+3PhpcaQo
ba7U5ohjOpHcV1SfDjCEvW06mj8QWNpr+3acAd928tiBAXLv5j4p2I+/8GOzak4I
Wg8ludjKRrjAhCMJ78lxgKnmlXW6C4aWm4JahPCaGCFiq1qCZAtRK46022SSWocp
wovTtjwokWWzStPKT9KFkNy3yg5P1g5kS6sGvfG5/dk6kVz6ZlXG5WG5C/MpC+Vk
6UabTqoCeipLoE50Zjmd3wKrq7XHEWWuoosdM29b9SPC+qiPAhzfZ8BlGMK/0Gsp
pTjBGoDY6zZuUgus43yhHqpePZ3YpBu8m3OmED5uSqKdaJli29BhE5wqWSMbekX8
gfGv9Shkx6WiXDCTppDz5o4mB0UomFBUdJNAF39pzY+1ulN8JGPZdof+0xaGFJVK
do5dUaTUoxC9F07D15OnoX6kq9ocZJzdevu9fQunfwD9GlmqZI6k3HMzPNyXvYdP
rJ6A7AN8fAT/6a/0EpzB70lJJMryWlNxj/bqNzjbs8NFIKUgqWBwtih6LzVnv7Al
5P15TkmnqkjGMxQy3BFS1vKjiwIrigvdRlynT56ajTOl8vAbGxtU55FGRb6F4JKp
soTtgn97828osc926tiAMJESfFZVFElxtQMELH4lOeWJVfsyRQaeyhCCjSoY0s15
tJu7zDGHTY0b1qbC6e+I1XuOEOlG9TIAhteBea3L0ydnDw0XdYdUwqtoIWTG7gru
VoJ8yrLhUw89DHBPqwy/6NDNYlUPA5L4ajir1+SxI9Fzd+ZhmWFwcntl9phSpYwV
9T6dl4158I3z6W0vtBsmu2cR+PZf/JhCw9nxgHcO7lX1qXhaxQ8XabFptSM09nJk
KN/thzPX3q2bdyVSfiyd8Flo1XH/UT8o1eTbfnxH/SepgGClRyxiNRwa+pvqJ22x
QbYm9YzxXVBGyPdpPwpWbX8cH8uKfpCQOJuB/ykLDLXJg4u5OSzrfXwUPy/BXcul
hKt6LuTBiN+NLBm1FWfALkZDVtCo7AdAYARHvHMNNxNMqx9PixaYwFCMMXmYJvnB
PKWN3T5jpY2oHRCKi31N/8stiyDUbwJhLfjSH1TLpxpYjWaS3BekHmsQUfSnU6Bo
/Sqxluve6P0nAc0HZ5p8fw2jLb/SfIPRF0rkty1imNfFzACntGi42z33S0l3Lyy8
zd/365m1AzFmoRZ1m8KmTNEvUHb4xxCIVerJJcPgVX35JOsgCrX42ey/1q+IeVD0
GBzLrrjMBMTAMh+G1Y6TTrM2iQcE/5RORwf/1kGfYo4xDZXfRQY/IepRointQB0K
MIAoWK+k6/1IjT3leQ3mIugC2NM9SilkgBfy8+3qP8Ljc36Hu8HCLkB+Z+yYD3ip
wJo1j4HqOYHtkE3S+EB0cI3jrJKlxCHATEYUAwqxi74d8LosZIZCPljdwjwS+976
7+VNM5QrVzqJyBm8tKvQR5mivM9WZAN48DyFaJn3RNvoGJ/5oqTaH5heZzMbYbaw
gWQHZnNOZm94eO8FZAicKcHipWyUO6ubzh65LOHHdrvLmTVk5m/E5q6uKeJB2Sgh
1eNmLP6Inicw8oxI31tQCXnch5pFrKOsRrN0AACZLUroWD0teS5sapo877siS+63
HuWGdSXIMIwxIaAQjgZpjWNZ7jvII5u2+6EbpuEOaK6GN+7xh/7sqahMarzxS9u0
gNPmp7hDJFD6XDOIaqrto90bebU07KtkgYRwJ2QR8FmeQUyTDlMVyGF3hy83DDDb
0tks2ZkOxxGHbQxTnVB7GbufZf/kQkwsfn714vbD+oPwYfnui0qAPDZhKxDhJDn7
zprPyz8DyzxBbyI5S8FV5W1xhpC9vQoSN82X8C15EmNUJp5142lV89N9KRO74J4y
R4MUZdC+dGzNxeNX0PtgFI8iJMpHYtZF1X2bR+5JZUJoHBx03OcEguOAbP/vdWSr
Erw8ELvWG3wxzYiTpT3Es+8nheSumrgnlRMbJQJBBUauJ9cfXLRuEXeSB1yYEuix
GZdIOkT7QU1KG7QadTnuwMk72hfe2pSO6YCmDNEAXVnJkT5v6cKjd4+YgrxEomKg
HK6g/nI2wwgNsGGXNmmgHDRqMJUPmCIDN9KK3aRq9cabl7Us2pY5ANHSZtTCaBjZ
GNReGqRL+HsHJ1Q7xIdXONml937w70UB0vZnpDBG2ixDH3IkRyylx1eCVXIZHAnM
CC2tAXHOmwpNi0Y+CHBp/DIzaUaME5oWDOI/hrWxPpSQdNZcRoiQRQJcVsxzGzvC
kjX9JrBrLmxT6QK8KjNvgiXFDlnd5QB0eYC6DuhJiyuTPQls1XPzzHng+wtyd1mx
vsJweQ6eUlHVh/rzUfmrlAFAU0wHBuHvCbhQM0c61U4mqETp02LbHNsvcVXg/m7K
PyVP5tgzC9ZozQOZCKZMdWfg4D2Kdft1FJ0j3KNHmXNPQCskyxel1nLAKObUg4O1
FweYLQJ42e8j338vAhAj6fP5bdk2ybntx18v0L+wWasZXGOCuE3+/s5g/7LBZtP1
OONPm3lcQ271H4HYeesrXaWihGaNpGQmUfZna2EyMNLW8k9+yKGavNikESXwjfNS
+2s/UhoSyaiM4qFi0tXRopIEZuYpRhb5/PLeylXCcI/4Pu0rrazu+Z8DdGiZN7d6
QMrnDq1wxfyybzv512nXm66rjuEPOlDxBlokoS/XInXsST/2pOzJ5fLU9YCEPt+X
g1sPuOP1yKAHWgJpjFLjvSw3ZEeMb+vCv+9j/NeCQr9RbQHq4SFzGtPxTzj88m4u
GZzAu1W5Oe3BWQovhOmt6NHOksxIMI9Uj5+P54xrIzInd6mIyEusrSMQr03MjyH9
+WdR0XI0mR2yRku4pjE0F4z6az2ehE3uKZN+gJpLD7h4QmgY5+IGWkcx0Dt2KX10
W1hT469AAVbWA47mooonxKM5QWmChruc7Ul82ojzzt60HdGCm3Ebei+UI4JVrlVt
r51tsW/yUvbdvQpIbyR5Bzl1TmKgzDUPu0lpMGXNu+yhkK9Xaf7uqBEZY2gVk+Ix
eOcXBm3nWU4+5vfk0D0fTNHIFZAgPWL8A+6S7xzLG9zv2ghx7Udv1mCfCSHIsih6
NkLmVI4Pl41x/Jrze4/DFGmRR/e6xPt9XapfzSY63ny6tPn4WeS9WaYzaI0MSdBJ
YIGv54x8lEwyj7RoZAkpfZZJ/uVqRsgKjaw/RPVmoRXdJ+MT7DMxM5t7dOXxvlPz
6khplQuY1OoWrp7VKZh4HZ9dkWp+P4zb/vZlnAPKHcIH3bvMoVKeE4tSUP9cXxqH
WElyqXTW6Zx6RBI1q8KfEsho3lQpw0kgfoFxuRpTMRqWf8CZS3SCIvEW0T10Wh6j
fDJZgew0GYsUsqYV6o8Q6L92g4paLyVIT+4AZx4kPp8qWTFM9aZ4KDYX/WbbsQKE
tGhhsmYxTTEV99/HbciT6u+mYs4ojEVT2nWSTl4mbaj9sH2boGi3B43xGWxIUBIG
6OPM4kgViNRvPc3uVmOxe65JTgzG//MC/EYaJkxr6d8KZTKcpAndc9XguumoAmgV
81HwhT2ZQgpVcdsFcHanotxaU6ptqEpW2yElLcwmZsiP6M64649VyTU1OnjESvbv
JhILrZpq4fGN1t30lwirIbo4Y1QqmbmVJOMc5eEoJujqns+FA+JLCBh2IAdyYRUN
94rz1UA5b4aaCTPwN2NvQHbmqIqcbGmZ72g8qF9qNyO0eo5PfXzlP5tNh5HoUzEL
cHwtB6HA94TsEAtdR1dzH1VbxdcCw83MhpMkHyXk6BFOeZibrhVTwU3uxjsXoeLq
MzH+aG+EfvMOhToqm1v0y0uN87l32SCKCY+L6lvz+nA8GF+Cre/lB+0r8ZTHshOh
AjNynVk/8LXPcfxNQwy4jueFQ9MHdY4Klr4IIUHsql6BJGzF9Vdp17JnIUiWUdPC
Mc+5Y63zxA44fQst9arF/3TXpa51WyNinB9uMI1BafT2l8sifpeKX2zQYcZmCMWD
vnRExSu9pm7QRcmn90XNuQPdWexlZBLMOJ4zsVtoiYcMWEcPrLfde3sYmI57XCPM
5ntgfw0vwP9Jz5SaHrZIiv23zELMCJwku+rxPdNrBYGW7f16Wj5usVtzsZkqi3LS
GBoFg2xwG1AI0oyC/E7WlJXLBeuLloaIqqE/+Mb78Vg3foPANrcGFLpHsTBQqLYx
Ud9+oHleizkYJQO6XeosafrzvgGJZh+Gdc10W2BbahruvC0sGH0OHD2fnlC6b0Dw
hsAunw91T1CxUx//g1+I3Y37HPpWYbczys//DqGMBbrOn0vaH9iGCFu8qXWFHTlV
jSV0lkWyQEDCAFgXat2PlYQ1VsSm3s5vhjTSm7bNsKRmx5X8tWtSModI5Am1Xw/F
QhXuC/dG1GX6siLa6B5PS8z7bdWAuRuex/hnOvJjQBT/OnYWlzzDeGr5Jom9gIrP
FADeyXOE5xJmCC/O/73IRKXSgkbDau6tMEXmowc03+KlSxewG1XKjg3znyLNT0qr
To5lXOidGmpkBG8HBPrxw9i6DAHYNzGgotMRvYJRvQPAD1xt1C6xJEi0ORLNNtPu
RF+w/cP42lSEbMQRgi283r1NzZP0c373yDCcVI8nLo0WtCVJRBVOfhiHd01X4PmP
WOJRCCOytVedTgSaaa+XIHrG7rRmaurVidLuIhERRNV68lxnrYCFdzkvrT68g0f+
DFnUTq0Fmfe/ApqZge5p/DG1m8GW/ytNj0GxOS5lBjSlBA8LJpGQADwYlFTw8vlI
NH9ERwfhZQvHMOL9i+EFeIf7GFYbTiBNRCiQAsGaeaG0OebQfLwAT3cOdb4r/MTg
LuMvxv0ZyKgji/lzYgpjaQB+rfGB2FCEbUXheieXr0udbQZHRYcu2MgNo371vRKv
RrjhYoFUrvdZOmK4Z1c76GKshn3Ky5CW6CWc7ZTPrAUv4TA8whIX39Lqx96JiSEs
MqCNdccSaJ72Pa9/tNoBQpwiYgG2+x+Rybi1GunN6yTcoB6sfcHjuPZsm1joZ5lS
tzCMqYw68chtt5f/GCdlZ99bdsOPG0R0F8FLnxFcmXdxWAo5Lr5g1pk/UjIZNYFl
u/I7vMfE1/NatUqFb5qjlOOzKNj4NPaJ/R6sr+Jvuu+RN9zPyJ2VSK/XInf9g+yk
gbOnIcLpfr68aY0rgLwPQML6ohi01E5qs536UPDL6EjipztCT1nhyoP1x0mJdFNR
DIaz5VeMOvKkxTi+LS17EySMDYsuJtCOsVLsfAAvkusHXiDdpZPGI36KfudLEPHA
LebPdb+rvnakWvucM6/oFJOJEFjk0joJGQWNxbxXsrv2/o5ZokTjRKpwD56WKnkR
Xe6rcp4dpkk/4RsU/LzU3pdHRsW4w3UydL8c5TGa52i7o3mCUq+GIy5m1CnBt1NE
yTL7u/mQYkejnJjGSsiqV6LzZ84Y3lJ2QRY6FUPrldCh0VRHflGLHIE538IzTuOi
rJW/cNbKP+m2UIke4oAXHIEqULUkbOJWkmsYhu3KLisu+25UJzdCm38CsnK+h+Vg
9MuOf/uXx5tXUyDqSclpsb63OsaodD+EqhKiLpVJEAIsrJZHufkJfBXLXyXHrRRS
EFQwPNqLkowII5ih+OofFGnprvDnNYz5uPk8NU0P30bzJ3im++oJHiYSP+aja05E
wt65ffdsXs6HrxGTw+4apKDrMs6aHzWVqQ9Zwy0lhLVCqMbTa15DTERXHkLCnf+V
YIU+OlnKTtU8CrWmdtrBQKPUJUx1hn0VchntUhmMEqHzJxT5uoK8BGnJCY//DCJi
ggTfRVAr+TqlIVCIE6Lvs2s9MVJL284kT1HD86MmlfEN5PggwTYt81/9oWLN/hzm
z+MpKu5pNGauvv4HjY5u9JS+3PJZt+oWDluPJifjekdwb+dq57Zkw5ayEbrREZX9
PbRpK/toEuf9W5s8GrFpGNap4HtSZFjK2TtY+wZ/kQAw1zLE3TvX2VbcBtYsJx9Y
G1RQDXuOVzYoMg4QnJwR38VI2TPK11jvD79I4t1hFwYgBNwlZu5eGajYQzbSV8an
rm7zrJnH0wcWaSfDL5DSGeOuzVMpR1d3DH9MqcK65Q/qvg/a3Y1hgJPQKygkjbIH
pjKps7f9mPPwezMFPjAb7RlkQ3m5KW54JemLSm0rvIieSFfV0l0rL4iNIX0DsJbo
N2xH38fAyiLqmK0CEcIvx37NXlH1zcUAlhUeEW6b6ZRWxAOBaWl/7N0TGAA2PTcg
U+fEmxDcB10GP7DS/mQ8iDgW7W9RWsFLnbCKgxsNG6XhWzn+CAzWZNZTJgcAS8Si
wUpam97pX4Mq4Exe7Tk6+nWEj7tzGD/j3llSHpfE8CuBS1sHCHZudLrXMaYHPc8S
m5l9Ps9JTM+PgnSvTNEpBqSlAaKZv2sfRP96TQjabgvR0aHANJ25DQJPzmwDc9Xb
is1k7ON/PRt5h3JpoUrqLobEdvCH+KRMlsVdQZzlad0FYr4M2MiScNWtKUsyel3p
LZTfKrpdFfMLyfBafJoUP1gJMISxHfioof4LWZIyzZKiRlbSQ52jNM1Oj904kGSN
mBkAOUye4rGlSL7bQIYtwwR6TzPnh2STrxnwGZ115k8G5fETKY9pXntPijWD0ZMt
LlXL/zjNytBcnwQP6jhhbMDgmONiVzXJPW1bV4sHxPyPYAMOETCgvXQrIJjkk19E
it3RnsAu3JhsEPWJXioxloiGJzkOMnCGyffDAQ5ns1UhK0Hxe29RvgfHaYT5Yp0a
9YP9cMImHKlT+bIGU6qu9ZL/aQzOg+7cgg2o0WwBxyc73CtsuJ5cRbI/5dpWyvzT
VQV+bs4eP2BxZi3r128nv4USwy47/oapXdvPKnCkYV4CVsqb0Gp7c/1EnEerq3Gj
sDCOlOoW4farAgqoFDT8pRvvAJJR8/T8c9O1RU+ASul43EhDRmFnV2Rc78Nyet/p
7WScSwC675XTVrSIus21toobB/bNbefc2/iFI70wJ2lT3nPmSxEvVriXv/jU6Cj4
Q3DEMJVFGxGBLr5K6o7V9CUbq2rqhyJE5Xkv5JxvCQdHtrNhpCI/DzE/fNXvPHlf
kDeqwnATBSh3axBEQgqVlVMCteCY7d79142GYDnlp/hTUW77xyoqgNBlrNp4UsR7
qEX/TR6XhDEHDYOkVlTgz1vY8Z0GPq7LcLA4EwvBfJZ1ZQdumT1atI2wL8qXmQoF
cn82v4u65cZaBw7/A0RnmLMEc4Wt3WuAoiN1xCUqfjcHXXXw83wRwuX9MXKOwZR/
h/LyTr8oYxjRaDAqanKGKnjKXYwf7j6AbEJC1qfKV6RgNcb1a+M2fw6ZD3PIqNjg
w/jG+E/EnqY/3skzCxWTpJmmIQxq7Egz2Wujda28xzZP0xklFrdHlnGurmsvqRiy
Hmj9IQBBiUkGvocgy5zK7ASEFraEwozmhR0+DSfzmW1XHrQyQNZh1Ay9TGhihGSP
Ho4QxfxgmRvChqRjs1uDQD4CV74dwuXKrgTbSz1JKAXadk21lFauUsFw/Ak4loYs
cnDwNOl2eaM5yuQ+nWbc1EryF5wpqbJRAjktnxOqr83CnyrXueHUQIcd+Qr6/nBy
pg/q7+TWR7peTLQu9j26JyFNznMlqhylD03/HfQin1VMgm3qoFpvFSJYHdSKOxk1
zqTD3wBXWvDTHuXGMLMcyks4gz7uC3HiYpHSFcj8hi1wWFfb8roETkgY3DgRIHM5
M6j/HGaj7TM1VLXeafYkBqOANAfZqJX6kW1u+cw1WaEAugxoU0uVt/Y3ne83VGn1
8y6yefpSKwQZzOXIf0Hs47zwX0B3nY5oGDxmXc80z2uAx/NK3lPNEI2sn++kd5m+
7u4Bv8YfqZYDU99+mPjhxLwFddJFvhK54zK/AKL7gZ6kloQyoKI/HHFyVYPoojzG
/g5Kitj4C+26+z7HPoJsQCxbvWKZtpzlAMn2WGItXKge4T00uYncP/BVBDJrkz5M
5PmRV54zdPq9NC0P1oAYyOfa/UuisZJTZyUtjFJj02eGBgrrl6MqDSNFSweLA8Ey
QXG2tb4Li1ISYhULwiF33DxX4X6tfhJC/TZZnm5Jd8Hdju1DTz8d+FS6yvDgo8sf
k5G4geZ6eZrBVNn6emlWh/CbRJYIsrDXjJvRlxwoc4sv8JN9vZABGzt1WIiIabbw
HEsJCEhYmyYiytLYh5qz54Pyd7ucxPsG9G/D5qmt8OYKyS3TptOrBX4+hRGhug1X
Cu1FCrypV3/2C3CN2vW8eLLNzOq4Ao/x2wf7Ks2z82i84Y92SscvR4H413g4QdOF
MOOQS6MLwRdmkxmCY20zTjHEiBLr5jlNmuCylBbSDGZMC6TRDWcr3wJYYihfjHdo
JXV13cKVzq6wjXvUp9hvN4vLP6jCAw7ECLq7/0YhE0CoN5NarLWxe4ysW+JTISUO
wbxO1badYv9Jkf6a7tsnMvHgiGncq4KV2R892md68AwAWsaCQCfZfsAs8floypO7
SyFUAP1yo1b54XeBS6WjzCj18/mLi80izLbZRNQUHDIkUo6Pf7nzEYl7UbBXPbuM
XdRSfUkw+LKUKxgjn91kBchkl0TN2SIjSVvbzT62zG2qexdbRvWo3H8Sp7+OOKVv
UCS+cZct1eMdrPkrCFBh6fpNsswu0LIc/y5JFnnvCYNNHx1lARiXdudvL6MP6fg0
FXBLc9LmJsDGTkH1XgzOK9v539i/YzxcwKF99z4w/oBdFgxzmIIyunfkogiqGyiE
ZvKjxGi9HvyR+P+VE+W6Hr9Zd5GvF9wG9g2hh7JGsV21fy1g1aMzpZe9pR7/Ghv1
3HB9DKOonDj1x6LJyM+jjCCInEkWgrfZKAyajn3HKvZJhFZXRhV5cZCnCZ5bMrBc
fKB0R1y5De0JGg9MSoGaDRIoU4X9MyZsV2TtXnSuLQd5IaeoeVYokBph3gpU3EXm
6+c7ihdfEV8OCZVAyEPqs7N1MRXaEZz8KkhPZ00a1AFKcFYjcQLIO3/wtfOIzwSY
j/vazOXu22JVm6lcKaWCaLDGs6lpHVpQUACNGPNYHwLmbL9g81AgmWYF3ws4QMUn
Nv9n5EJ9l25IlUtlHkppbsIz32U3nggHyxTPYnBQO9mvz7L6iZKBGUjlYUJpx/m3
TIxnF9P3pPQGFSuEEeE8j0HUwC95FnqWUQQ3O918MLuIC32kqYexjdzm7ahqn8BX
D7P/PtOpqsnMs43ldM2swSPUwwU+gUwR+FWOJHnucPYmIuiNOvpfQhJsKA2stjU/
Kb/8aoCGWXNww7ns7xfydKKRAaFS2nad/BaqV85ufKahaGdRs6Zpp8Druj1Ooc/J
rqOKXq/42lFqR8VYCvUlYZbmYYHEBgOuF0BzQMUhaYaE/5NINrWwYeoUJl1SFVY6
eJRVFNQvsfiWeMZ0Bc2mckBvHQ3PmdDd71LDAzDz/9WxyAa80/Wc9sDW6ALvx6yw
bmA1no+4iILe66BFPucbk0mca4nxDc3LhL7KNPujYsCWxEYgnZjpEYR8GfRD7Vin
2jINlSMPJlYMZkOfbpH9H/JIaIvir+BoZ4lrt0wqersfZB93Ao8eyLlLlkuqGq/8
l/OU5KfIgsBLTBiVpDZl12ytl00ZfjWqARLW9Y4dWHY+MQl/plv9SEFLRcpum89p
HL7/IBmCbxETN67MKNp3GzglXGnlWMYdLUedhLaigXJ6JIkLPeAZdpQH7+goIr2w
uqBrCNnOjnEMSSG/QpikGMT9orYl0RHZVixP+2FWKerq6jgkEfsS0TgZ6VNRe6jl
8xoK7RfwfkQgkGtgVJPQbPnsIbBZizZe46w6TBZMzDn5SVVbrxxq/SoXr6P9Bi7C
+8jsBrz/8hUsc6R0ab1Wz7Xc9yFyzBlFNaxjlQszeu+OdIJog76MYjb+v12IkfHX
TdONlev+y142Vfxhe4Ytvue6/bLjGmXmM3cPwkLYGllsbnkjGqtnFg6y9fRrVviJ
3VtO49dmlmiKLBJprfh1Tl0xpw1RTA/6qtuRvobdPMi3uiemYDL8oSlOhukIbqr1
XIkV2ZhGJPEdAwZlLiAUriq+gFysOha3rrLWygO+Wtbr8Lnar9Qg190GTcY5YleS
FsXO/OugpkIrmLLno7syKrWcQS/R/NxOt4Oqen7CTzw2aZ36JEIviKieY0DqerWO
kscSqkiWr/ddz1UE2qnfm17Roe1H6RIbdJxPWguRQazJ2l2I4pwwbeE4ZNOONohY
0/SUPNl3Y6ryCNPH404KwZkBH2NHh0ZnJ4y1KcbUbWiQvtgbrmrI7Glhi+nGw5Ek
pfvePzPtoqWo3sIhPijOh4pqAQdpzOwrcnmr512PMwefU2dYfKvaaHCX9skvxjXO
YW2goe1kQVitFSDXqlJv/JjjTFv+w9ghaTHdwlJ8ybQ0P0Cnw18CVYc03qUcU07V
mtW18tye/lmvn+topomQo5eFvrVTmtuAxoe8YDN6zEw0eLfGIP3sxRB8AxdccMuz
8fKnNryiWTyS93jt8QU+j5/DYiDsUfMqVBApGVWCeRUJkCjtQaoL3aOZJrKIz4Wo
xfhmEGkDSY0KoO0i/rmeB4g9Gql1bGzmtYSXHVs+KjUTss9nPEx8gundXCNFdJSj
lrIxVeVYr6+cgUum1Vdr1v8SACnZllnVdWG2yavv3tiB6gz8nvHeNneBiAoP3CrA
x2/7EOjFxVYVQm6tbamfXdiwC5TBgcA47lL3UNIBkeAgrSS09qu/gM9m5jQ+gOvD
t1P9Irn6gZGQwWjdhHxmu7H3BgIhkHrdL6vpqJqE/RRtvcFoCY0nHYkDrBnpf0RA
KzphKUrIixZ40627GHb6YqgX4mPKVk+QXrzSU7Xc6CE0NddWpRYuxJENSntsuUq5
2WZix8jD4ODSxn1YlgKB4sUC9pMTi3Cf/ihAQGZIA4oVuLMVCarvqViu5IMQihWW
P6BSi4+66EogeFVs3hFUfTGLsFtZkF8WQzvU+mRhOUeiKvoyRgnkmp18Fv25D2QJ
+hHeE0d5Lc02DBnr1AUbcLSZjLfiw9nr7Ezg4+9fsAoCGJSK4pzwgSJ5adrMFm2I
3rvOmDRbS4eEM7wIP3SHTm2JtlFndpfZlNXHYtxJ1AQoqzB9fzbuGKpYPIMIBUQV
oG18NOQ7kzZ+AH8tzGCVxeScUV665B03jEmnI/zuv+q8JldJnwbfRMF4V//+gEvy
Hn+2LC/zgBOTC+vlqk4KlV8q8xfyHTfGYgWXkN9DSUVIZLahE7ud+yEJGUh5Df9s
czuVwmKMdFssMkFS9CP8XPx7URh6G6gCgb5pmutbTkIVm/rWr47Eaj5jmRRekJ83
KKY1xUHgh2r9AmfFP+eTOsi3HqWifnmeV1AzkvmCJD7dYWKYj6jYwv5dnxIp0iY4
Wae7wo+37G98GBtQmzvU7sfvvKZY2dsrt8e3wjkDkpU2iwwzeuv9qC2DE99/J9pu
qZx4tEIli9fumFldTbBcZZno7hmAO3OluCIdsJbfctwgcU3+kYgm5i8my4ZIWlL4
/HA/jsJVYeI+CuK0iWMZ+DE6yNUUASKqwWAXL2gX/k0VKxWc+vchILaDRb58h2ay
bd7pydons1ZC3CfFFJ54f15ZxjsUo2ZMvQoA8gqHFkkio9gG8JMCGAmnI7UeIXHi
l4rmWd6F9sz0DS9TUrpwnzCRzvGWKWOjwk8pqOoIn930ERhFYrfFlgI1mX8L5fhc
qa0Ob8RCLNPkOJCu9a4qGc1cyt6HgGi+DWHmuri79r54wBV1AfUtR7bx0pHOfrCC
Xaqqn7vpnOo0rss7EnmofOSrQ+5bym4VIrqNnJPlk0ShgNzglhpGHOwTYWvTSCBO
avRK1aLf6bR+GNoX4PN7Ay0tFh4lM4zE9dHCQ4eh4XILgESQ5JSBFxMbSoIs36Eg
NsUC4hEWecPzl4Y1rlNDUeOQ/cSx0eHO3FOI/fzj/tYw0IYHbaZvkz3mXzZr69e8
cAicsYvZ3ZLZaZizYajnE6Rz4h1qHR2U4pwZllHgQr3V2Asn45eoju+cov0guLTl
6uueoqG1dvZI8XUFzjDREs0gwMxTwxHz5u2XsJDi6b1PPuXS0NvpTJpOaU+2Lw0C
BRYAE6m12xlom8bj26JkGxrCIDib7U4NiLSs0TicyEunwYJFxcbnQEwke/zIBsjh
Ig6N5lr7r84tudxMmObxRdKX8JMHc8nAnWl+A0yqpRltUEvZg96Yu3JYobSidZgs
IrV3j8r8dIgIeJbsJCNYEv6B3FVjcIuITkVkZ0wJdduH0/YDc7RFyo61A9ipVfHi
QVFnanhIcEW0I+l6pa+nlJeMyBXwIE+yNrLnlmUH00xI6kw5lUz1TN2/JLUV1uHg
qH5pZoaIgZZtOMhDnl8CD7/tbt4rHpX1CaTc1nDgEeVgxmd15pguweCwGwOU5zNJ
ps+x+FfOsAclMy81pElHxdktFTdVQKowJpiPLiuH5a4BEMQO4dvG7/0udrovCgKN
pwx9KjGTCHV/Vf7QtcHQzhz+/QSLppwfnJYuu629jsZ96ent/MrsrMx72rVIqF1S
YOVgoxDAgY9Hirv/pBDfbTLffR7y6ey8HHvOyTdqER7/XFd66PZEkrQe8znvfNJO
KAmTPVxtiRHw41CMOVZK5+xGaeLXyLMxpEFp2YJ6EecaWwlNbDuCWumzoBERrrUx
bm4VXyTxM1FSbQmyW4a/mGj+VzyR8mXeS8mnka0nhJJHcxNIfYTYBT23BUHn6EcS
UsSHE9QGajtiPQBgksIlFvkEJOC4GTzBG2/grv4JCVfw3npSjVqbkckh33p6ASvh
Z2+8HA5hup2nl5VUMoE5Dmc6q33P+UFjX0jMnHSrTEDhm/qlvpzfas2LIqGgapBU
YMLMSbrb4gAKI4Xvz/kZq29cf/arVqlaKccUoa9LJEKU3Y+IH2GbJzj8p8w1dMFW
+H5m4CmGVqsWX/Hwa4GpSRqzfk4p7NRIO3kjgDskKFs7GicO7TK+fHObrkA46by/
dXyBHVR8yXon4PSqU2N3mOSE7Xb7hPl9h1Of/6a+iqSMBS4DHCO+jePZu0O4VK/C
JgLCBZnb6kA4li98feOlJknOLc7Y0RNjOQJdznMlSeq6EJc7yyX/yqMtOhFeImr+
M4Wr1jiXuHL6hOQE67mDPHfLdzjc3q4vSkxLrn1wAC9TYKZcpQAnn+1hFVd23AfU
1ofxJqkMGt9LAS5b6a4fRzeO9dkGhur8QiCHRkIbAXS8y8hyIMM8Tu8CY6SaykGt
NaXN/UJSKUsYIdB+OqxXeLQiYVi398VwHehXTaVa1A3NZJv8zNigxkMc3Y8z0aUt
1x9B5WspAXf06YW+EO46Eoxkbhx96kNSpqXzmyJ+MjBqvPpHogJB9b7iq3MVwusb
5n3SCvtQotZ9JXwLQ2ok5nymdqNM8PJpHUn76xhWoI6KDDuA1uW4EC/sW45g7CUp
vRyT0Q3MArtNMZyGuEIeli/gDAesZ/fE19h/23TNAd+xiaiY0kVpvlvVOsLCRMcT
77Dd2jvIepJ8x9thhuagvir3umEYa68BxwMKxczAPNDO4Mjrw9OzDV9QG8dBvmQL
45waWtXOFM79aHnZxU73sJpOmB1vEmvkFwV9M6dOdok+s9xB6rFQSvu1n3QMzUT9
20JojKHjcANkUoL6Rs+JpEIw9xLF24wQXCsnHcCgRMgYMHs/+KTZZljp0e1fsgoH
onx4uLZ+WNlci4kZI9v1adMM7lrj8fIMHM+0Cir77fVxMZYL44RO0RmxeoTmXfpc
6vE2U7aeWoPGylkj6Wm+uaGqlmIfU0f1rwJ008+ynyTpzv13P5AHHRHxMEZsBhFY
G/DozFthKS/HR77l1mZlETkLHflCAGDFSJNQW3+sXB4gYN+gmU2S06whq/BvjuJe
/YKsLH8S+P7FoSo3Q4tF9PL0hlJX+z8ALvTM+BwH9wxucJXQV3ezVlyef/0lPuHl
k85gd0nx9BW+vgP+NrS5ihq8DLpAN0VKTOr5KTYBVdMYfQqFcnryC6hB9UNZwSXW
g0eYGn8xLlK2NJsswi/tS2NnnqCZaZlT0VDYU3LHFqQgYXsrW5oP72xDdboLEo5H
Tk/QqIYhyt2pViwX8zyLnE8sJExWKP0U6kx2NT28aFEb8fuR7GAPnDepAr6FkYxF
g/6wmm+eabJ/hgkok1LEdn4VSxUUw+HflEH/R6YR8HsAbVN/Bfe/6vnQB9nIYAPf
w/Tmtq38kDzN3AzhrflQy07kJ/wAFN4gGsv+sFHZUJMLGg810PqD60qw2SHrIPHg
L9WCf4rPPBDHwNt3odG9qb0iYwRXHOljxZ0/v6JP7ilBYUVkRKBhpIrkOyU9zLVM
szt9ISMss7RDltORveURcNAsCvfrSi6F2oBOBixytP27UWydadte2tOUf4Op/oKA
2hYx+WgRpMzX39jFtnI/0mAuYbO/s5BkwDNwZdLgAd2GGwXgxdUGHtNgEullFOhK
hMIagvGlUNA4pOYEY8eNJFxJktAsxOcxFCf3a8zI9Tmt6Q7C3PQRee/OasNsk5kM
oNKm5baZUglbm8OfXGkZrFNMZHwAC3u6CA192otyL7+6enmP75HPcYva7yvMoNrQ
JAkzy6jE7HbWJIfbrX58D6zXaPM6a76O5GLVsNcSUXHcU7S0GftfLXpMSjGVQ6ny
fnvxEnSyS+nj0eBkg8hbcZkt6xZhgjB0Wm0wValG76FMatiGcvQqy156y0KtkORE
o9mt3vhnZjvcItqjNj3j1RKEmua79zMw0FwW6GrDM6ngiLRpHPSlTGzl+Dy9FMLx
LtYVFYAcP3Y/w7KqUYZaYXUd4rv54OZTzexK/SlK0lmwvfwUglyGSnSGQxuKF3J5
M6LtSLoP1GmapSLtalLBAnUWxN7aWUsEJuSkXDEpBEoYtyC6ZJMqXZalhoJvaJOL
7o24xsddDeYGLfqojZwMJfsITs6WdQZw2xIOqFPHYzhpMmkZI5WnzWHer00RALWQ
I88lLvYZfthnHS5i/sdsH4vEzFU2SZpY1ZO+NEX7EI76okmac7B/ayTsK1Hj95s5
lwTNGl9Z6Ujk4WE91iZ63vIVQoaMMxfwBkCx+DDijRhpd6jf7Pv2QTWmJwf3tA1z
14RdZOPMX6ds41cCY1y8HXKapr63GB81s+z3r+MtmSSrpfKyfX6FAruwuJnPpb2y
ssEnMu+rTj5m4BmOb3IpVDNXbfygCE0OvF1l7GNBWD8Ie8V5Iz5q2jIeaNSFlQt7
BtGNOHcU9bzxMks1hLJw62gUAdFbGdPP7cy/RFvbmijvYque53jyHdCWUHnuYwQM
P4l1/z+TmjaV5W/0c0qGk6Judl08DZx/vDSdJKAS9EKtuVsezhVyXNxu48C9Afn8
rtTm98v8m4BAp97UvOZcxRDpERdMBjhuq0vI2nqA05SdOccWItff4+bdQTsUNqhu
iJScw1chPg12oYOulbylq4uHrAh3WLV7ljc6pI0p7ombly8sULuB6i4WL3GC15en
kzCVITS2UmxTQQErxbOnZRQsWS0gTnmBvb7JDLid1WcccufbreahTo7HcgpuTUZV
f+VGxhmtLZmeILIwACbfrOfEP5iSmAOSVa0IqkdLgyDloJOIkk1uY6iVAUApPgQS
NUJvgmSYt7LfftUMK65GrOAL8+QlGp2ERuJSav05YUbIZVvJbtXU9v9zhluPE64F
2Ng2izQhihnSiVPdy+HNiJdnDoBs5/l66AS3sKfEZypeVPxFGkl9PXBH1tIXZgwE
pn00+B7P6blqe46FRgC++loFw0oQc1UyqI7OwsnPaAIsC/+45xcjgNyN2EHJVkVw
0mA8Ozd8jHOaX6Svzeyo/DFev+bs2YGBidzMLt0vq0aFtuy+nxX0PlRNfix/J/Om
/CIeC60ZlVz613UH85swJsLzuI57lbSHTvVv6XskCzXgNMct05pq92qIRDa1ErMz
qaU6IkZS6NNL7T7O17Db2aaEOWUpO2E7MoT3k+V7DjXnsVTosoYVZQJXlmEyg988
e2sqVmm8QxvEVNR1hsBqu1IfFlhhuJqe8u0Rm7raVG4ACTgeRaUIDWSryg5Cdu5W
RbwBLWWzqb+FeIqs09zTNovcpQG0TnUAekmokfdNsLdH30gfZeuJIp82AEtVKyzX
RfdzQnCxIuCMvIGETD5OpCMb6HpommHDXShc1AJ7EiN5+qaAIj4V5/f42nW2KShi
kSX3OPlYylGYebOPX7ls3CEdGtyvz9LV0KOmPW2faqu5ClCMcTifWfpVRb0yrTi5
NGH430KXkBiSD1DN82Vv/yPJiwefwhgiEFSYi5AMB1lLO6tsOPFEs2DAaKqS2hXA
fKf8oMmn4ZbS+QmWVKktsLe1o3AdoWo18HomCVFgnoeMq5Ddk/qDEsS+BbRpCYYx
EMpScQ8CdgLgzw2tRabE59ORk9nVt/lGvtgRB7AVwSsLlBeIXE+cc5h4S6yorj00
wFxUZ3oUCXhBd7lxh/1IXVUaph4KtrXx3SNf9/bh5z0Ci5cAGAMn17mwYnGRZLjm
mYtLK4/haHl/V+CrMDv87JVqMHbcY5YZbpswBGYiEV4IFgVq51CY9Z3e9tkSsTl7
h9Wcyk+1CmGuMHuubLheK7MycX1Hley1FMZyfD6/iEH+zhbfazmA4QP/l898x2Eo
2+ol2fVyPDTYqirUJpMBYFwUQtJwNP24Nz9v3NM/Xu/zErj0ye3X+pnlvujD7X25
6vLH5zyf6BL4IFfUlRIxRsa4MCuWhY2WpCD8YhDf3FLHyRJAcgpAU3ncpj1vao8j
wm5ng+oXFiPpoI51lCrwBJgLhXx67Ymbbbh5nBt9wiMDpQSNi8XL/CXax++D/1JQ
BaV5F/Zm/+LNkYEzsqsJE5Pb9JzvSxvpEkdZR1MrvEft4S8UnFdbtIgke2QCoQvc
RDABHjZCmvXh5EdEHeg0hD49y6C0W8u8YSKXUxhypvf/PzxhKhn4K0ozaNiAccyj
EhrGop1ADT6IAjRHMsY1nwSlx/c/eUFn46cGkizrFuHEePSfKp9uR5SqaeoEabGX
zMQCKFTf3SwxBaZk27NoR2KA1KC+z2KKI6N3s+GcM1AyIux52nafy2ikMvoHiWC0
MDR029pTtN8sSul8ZJe5r+h818zTolgjkQ0Cjq47/yqZ7oXRftOvjMhiEUulGuCz
1iP0qiAuJ1qenuNtwHmx717tm2TS4sIZsuWrLjTlxBpP47vv744ku5HoYK+1kVtf
VFi7KIEGjthcdoDDfavcKDPWeAvQF22hGjsFwi8PQyo2crjyp3N60D8eAjCkjD9J
cleLF6AWrAOVaOMGrOdz1AxXEK+akM3866PpKAs318lOZZ059X9WKPXXNYdCS4zm
JECYUhlnpF12WkDVs8SqRky90aM1S0M4lHk4h+tZP/KupqtwPOCsy2H332QK3y6u
r0lPDFUWlX0SIlr6J39I4Y++MMSbm0AkvF8QuTtAqnZh4We17Xr65FeIisKUYqoA
LGsKtykYa/oTldqoHdFUq5+3GIZWZMLP+fYFreSFTe6RkJd+c0gVRkw6Ag/GBJIB
hK8FgBddtxv4e30+pAchWh5fASAS6VuZhes41s0hW/RD+Wpxzj5SjaLozCXEh5/t
gYJGWT8ZVWGCeu/i37GtvGK2mAvLtJikVnQcYU95lG8KXrTSCCfwhEx1ScfZ1FRW
KhGCOoz7vwlPun23788t653e0mlR3x0FB+8hGhE9lXFuS+JwCFWlfKeMBUtEvook
a1pgMTCzp7QO89evoQWFpWK1kHFJ+sCa71pBdqnuU08/8ssW7XVnLmRtMaJBq8We
i2ewP3dUg21Q+VRa8Gw3bciAmWKDOhWpi4sv2+GZeFIcbIzxmc4T9759ECxpEajN
zRDRr3LViJzi/JIY33JGe+k+b07mTTfZ+t/Yr2DFgSGMmqzAhK/kAKpWpELOyay4
gGOYiinFHHsCj3GOwTAOhWvelRbN9BvE0/3j3o9lJLmFLJr4nwjaqTuP4U0hYxh8
ISE+00xLbCAB5aDOa+0LO5/Gp9oRBbvxuBlzEBxs6g22HKU015eVLle+OeY6vNhf
5cP6A/htb3rq9bRTXf77s6cAibQVoBBLMtKCUi2SHB3AtGpYFdRbR5x42mlfRKA+
CdJWuy0oy1K0QG/iNBOPY7Q1+9M3ILYM8wVm6bYy15dr6559SsCr4oHWp1qcAtsi
GdtCp91SpfaJ1ZfcD7vnFntUiqo70/NdLwmGCnwzK6ualxkyjZjEc7CvmI9W8lzN
TE6eu+D5hftLmkvKXpywuN0uCG7pYfR42n5lIg0D8EVv8HLGFzKc0mhynhdYGYOF
/PKGv856Ivy5zHz6pkBMSnIrN5O4zIpcqS7xKAuwxC/MQVjcFJzAKjiix0XOXf2K
5cQxjpwqdReSHb8V4bpGcaSHxW9Bt1dxeitoyxrHGUTMi//sMBHk7fM3AP06yiJA
/7tG3cFK0MyFfIj3UH0chukIXLRjf5nu3/NJxSwe6KlJnYF0N8H85pG83O+lbdZm
YmK59iGtDaN62MtCsKVo6MbpfrOPYoWUMWmXbtqXX5a0avE5MaY9fzPIo2mXTdtY
G/IeS/aTMxODXTphrbUdYVjTcy/vzBf/QxLg3n4xV/J6gNWN3OlKwh+igJm6NX4N
cl7V74TCmQFhcNg/FLeOcyMLEy+9Gq/52TUtAlj0ZMxTtqWwXnyJyRihZqpZIvjj
fdHc+dQoM5LHk07aV7R+nkPTpIqreWFYsUS7KE88IZILg0IbrDTn6T4RN1JQLgur
Ycd3pIrV4EuUmOE/t3bR9pmkiSWa92UH8qXM/02TznddhSipGogI383i0UbJJ7yY
GEXcNl4Qkb4YntiwrrVAj6w7rP9lXX1joT3qm5aH1kW1YsL/0/03iRvBuBLhxFzE
L7MM3nyXEbm7onvR9qziU3nbB/P1o6WqLaWKfYxw3OTX0GCTKytLc0Z1M8HQbQgr
oraHzP0Eedn3kK8q7nosTepGqsC1u4p/DLFhUSDxTL8a8u5CmCa2plk3EWQRnJr7
CCVRU5E+3zs3mtgWsvRzqotH9SxA74pOkYz2RbPL8BcuuMtWCvhEpKexGxph0oPc
d0KRw8n85wsvwbKHArkFlR/Bp2pj3W+SfyQd3zNTS0ARgqxnF+2ohbMWTB138kiq
yHncxoEFxhWiR1VB0sxwaeTGd6K0V/v+WtsQ1WFo/aRcXGUdKxExbV5ju7gePqRc
Rto3HhGwGZAIhxfzctiJJ4oub0LeHEfC2DvgTUQho/gNvFBT1rciusvrwLcawREY
3Z42CqH83vpDYVZEXWsfxeRVmlJyBATAzTkxl63M2YxUcSOC/Jri0HR41CaBlxqc
IkFPwGlULPaHlLChZVo0/WPdqO6R4tC+gGMYN0SVwl9SfF0rJHm1s1Q+DY/3Ojex
h6gD91HzqZtzQ8OOH6rQZx0AzuPl0a+SkEjY9qJUWJ2vOKSKhL45kpEprBb6sltj
n+WuW9i29zPqklkTk1Y6qNXeTp9LaqdFVxqj++i3+tDjCtH6ddfc/7tvg+Zr5EJa
UPwHWUz+aG7gpEafM4JBnKY1Uw78lGHaUJrj4vDGTRjSkHVw9kS2+OPYrVEwCjbP
MLDW+GCP8Phpk7qWpAabqPsuR4QbLMMIO22+oQmpYMvHA+fcaQeakg70QQRnXLxm
8barbjYpe7yb1aFbEI809GfX0+OPi0SuRTopv85QbdC/gOrXYlMwkcgtht72eH2w
pDB012De3hJrIP5m9xboosQxZAFv+Fs/k+vQZX3no1eOCqAGfzOzz6omOZIfObO1
eZFg2/u37Fi8xoOY4+qlH8vZrHcw1utmFUt7A4vf/JlaFk9MeGqKtXDEbMEY1T9R
GIoVmJj7BHSSG0o5Ltger9MBemh+vvBd3RWJijGxmNXSLt+eM/iYHgxnAsehf1LW
i1sowjD3MxyDkOXQFC8t8oK0pEKCw6+UmNHoYHeNg1gK3WsuvpNNpUy92J7MtoZH
viu4cwYrQDnCfoO3jE2GO960JjvpX9EucYPdv5GkpWRzT+lLQynkLqZf56fRsyGj
uQbmfJxU+d/MUC9A9fCyIIemcoXqs54EjXik/1sOeOKR+0in3Xl/ulW14UKUU13t
7SjbrJsA2ArVwnrKNM6kXXhySTQElMYf7xehZDpRujo0ocoHeVQCadL2uyFmbbmq
Od5KAuu1Pgp8lvHRQk8EqA==
`pragma protect end_protected
