// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rUpAJ2LxO8Cy0Ufxq9SsboSJLNUS5Ih4652/c2OX4XARpOAdBNuKzpIqHOkpmz7Z
2jJj8twTVixj3eX0TwPcfjIcj+YuqwJaJK0eEVSqatspQc68YgK3W0ZslfY0VqRS
L+bQTr9brkRlOmSurqAfA7Uuw2R/oN1K/5ntey3eqFw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7536)
5wymdYfB6ujyMQ04he5hJUEmjsyZhwJaKcuMwTHmqvHZj6xF9gaoPghTuCZ6yGSR
ku44S39wIPvhVHLvhdTtyeGb/aIS1s6seBY6gZkzD0W8cN4nw3C7DMuhMaCgB716
JxTkJ1qoAUA3E5C7Q7K44HoiCJR7Nn4dR/VATQ3gsGSb3OQi4s4DcfM4OqdZI28z
/F+xZOqpIimITuQxq4WQwRbRpXUfBOOiNLPb6YWhqRjlTVjru6fxu0LGvlb4RxiL
lptf+Uj5HT8YWdHEn0fqm7WWixvNPoy2cchBxNHGvtK5c/rg8mD39zkVz7CMadJd
3pafI2n2rMMfvdTiSz2PIDi21QO2pWxuF668h9gRw1nGN06xUjDX8b54KXTRnxGT
9lZDwut0vM//fOaGglKP0sL3w2nzyoqTWeILmQLoFqbsNvslgOIHio2VTqFmZ1v7
tVRn2KjFtTg5u1GA5JVTQLXsulscXnKCkCgdzTEjZgRADOQC1xQo9rDSTs9KDiw5
46iMR/MGhM1GaoIkFwq3/IWAl5MK3ZXnMOiEBIDk0QzCl4bUenFroo/wRNnO/4UK
QW1VMCW/7kKif2my0U7m6OMYwLIecilKAmOX5O3xio6vOnLXpb4Sk9Lc4fr4xGPq
TPedtQs+8vgFXNAmw0ZJUFRNxbs3V8fEGIMG2dpUMZBwmFPu1Ui45xW/L4DUNIUz
JyqEQQ+PDcag1R2uH1mXFHb+bg10cJhisBQqKhp3kuXOA9kXqBcqZ2KCJ/r68eih
hUHteYL5ogafeU29KJ5MB6RiIUfjXVEX2x/Q7GavaPmz6cc+8d0ylmc/2Vfqe3x/
VZgqXBmTtSwX9awsK6GHOfTm5nT/1qjEt5l8K3RZlpkwRscE+2+s2SCWucm6+pFT
X9w+Pw9/bEwumorVXBBjnOgve9Hw4WKNPNIXMcgYqwhuoPbrCTu+2mggZikUVvS1
sM9nVxd7uBhtBJTJqtO1fT89T6hVGSBNluPQ6gtL/pG5o/uGB0b39iXF+rwVxH3R
u/xjZ//KMAWK25gpdjhOzJgNbn6cmcfB4G3DnxEHs5Omcujy/Pbesl2vkRJ+bqdb
lnjaA88NLgaUSXw9uvWBvgcnx4l0upQrHFUZrbgEdqifvQ5Iz2vuzUzgKI8PGEdS
JtOPBXfyq3re1faCML+GGam67Hv7z7yHPHTeYjT5sSHYlSrj8yEuBWIwcUCZrqDx
qe2Fc1dwa+ox8U/RmkgwWW9g5lOeluHrLK9ZG1od/0q4aCL+tVIhL7vopJjh/Cng
nZs8kWMI6QdFFQVMzwO25Tx5CD+BB3zBNnkpE9oWaRxUtxKrCgxhlOG+trrGEVJl
WaDgD58zuD5qzc82iLSN/4SBubQIHFVINa72ePVF9CTVPdc7+JNwbr0GjiCl0/6s
9dVCV9o4Edo+02oj8TpdtEQGyu5AB6kgJs2CSoHipc2ldkmYKYec0f4CPrAQYoTA
IYZ6b/mH32stj0Av3rxVDWJLoBhB5ve75BIQ366TV1v2HrUMrreBfIqxurT4S2Gf
pg52oopABQKnjy+Qd8ewCg92M9FfS9nS797LeBw5IrPoglX2IPWO/YQeuU6BEFUY
m846s0D1pP1/SnsGAJbeh9pU90XMW0aMk4Y1wn0Ap0v5EVinoWRXKJlh9lvx3m9s
IXmIqUb/TMZAhPQy05gMHaNFjkAFq/pKfWYkUkGFz9SWn0YHcr4JfdGWYElfSfZA
iDA7Wd9D/0Y6itrA+etXRpyo0ugg/rWnVIeIx1m5lo5ZR/NEocIptgFIYI3lIjnM
pdv13R8oj+okg0jUMaTa/6V9geONetjt4aGnwv0F0BhUzqT5cCbuAmN818P2RIRA
dNIM7x3rrqu1a70n+CHp1uV0iYAKRt+baWzWGzSgXVB7V5gBjuEvyh0R9ypGX8V7
/ngCL9iR1g8wUxxxQ2NWY0ftLveAX9Q5ryFTwQkg4jsYf2yKZILKTLb8SqvSTZC6
1Q9reAfrb3qOcsnlUgfY1c9+hvzsCfzckc+KMLn63Y9bOMmKsSzRrcR7VO8lB55t
QSOx7v9zucUDKD00auXkWxGFVcToW+SbPlUGs8f5CUezPNfVBmuctpbwfLqsBWAV
4lj0UZFeudVNb4ZgxERsAFKodYxKlsn9uRsU+Ut9Cv5FqTRFsirb54aHF3MnQEhZ
mtlBeIOr2drjQs/C0Glx9pPiU6wPFzokwXJHLhpp8ZsRgIBJHLn+xl4l0A8dgYmM
jPfuUiTU4cg3UEuFBFu9Rus8q012TQgDTHozIi6dFKstzK5o0H7I28rulFJt7VKz
mq3B5K3Vs6UWBFUufTkM4C/sozPn3IfHXh8lH8ICQEsxcj2X2B3BKpRdiYxggMvP
1w++AvgVkCB03yMh1AL0vFwXanU6VpbT0jAB1CvqF2MpI+9QBMf7KqWlLA74Z0jG
yZWoJdA0Mp3fgnu2AjASb+qxzl7cXA+RjB5l7puAXgz/n0zNqMDYhNR59r0Oln9m
2h+qU5gDdHDDytRfYcdeiRbcljGyvqdxln1ca+P9wP7mnBzBgoemTXCkMlNIpIIF
BGdar1jT+CX4A6lpYDqpP6nYGXoPyRKPLbqUDv/t6WIKOZPB6z1CRv8xugwQwGO3
V+yIO1+MP1786Lx7PXv42Pq9FmgM69qJXeej/9025F1SFSi4Pb6eJJ/SnTy7dhqg
vPPx8kDs10qjIO2lCjj2zeVpj1UtW6XVvXFEbuk5jGvtPvkPFBePVta/5HoTOgVp
vZnbRbN1HAZRF2yvNxS1tzr//qV0cGyibWipb0APbvTHfScI4EWwz9mtunVDnAPZ
O264Q4x1WquJ3BTsI5uwHBiSX4H6XHGPoEBEcTrGI39Hp0MIC6tRyTxwaYLz3Ued
fodua6W/yzSSwgR8waUPHi/TG5t4qCuRg2dud0YXwNLJ4YHDeR5NWy54wDRKnzau
Wc2AaSr8ohe9GzarxYGEJuglwXPNp8GhU4YX4xsWyVQm69H3ORL05Cuery1x/yhn
haa2uNl72RTbmMuoLOldxKf1uY9/np3TqYRUkNWHpNuPSw+4YQLoSfE/hju4Xt0s
H+74exPDfhYw4f2f2iJrO98MkFVEuHtmXUmUfzcwTOA/coKmYr++NCEugqnLHhmd
VZkcW88ZdJNAmU1lWDYi7673kJj9ZNAh2V3FoeEJ+1C1jbeMBJyY5sy/v52PZwkS
tpcgfcQ7NWsUxfcgxRhKLu6YxZX6XReSdj8Uw+bMBphwwbUSt8ZvXImdLddGlsoJ
W42MOwgP693f9TTT1cWbVb4je91WRGcwx6CWz4TlMdW4mTsAfOXlKX9qAk+prjM3
qZ9h2KPu7kQd2uNQpxDLPhwkcgiir6Di8xR9iHyIgD3+sTH9hpLVW6eumuwPFATY
DSYtB3qqGA0Gj+N22mFDuXS2C1fjDJ5wmFIUTffwj1mmrVIKjvFkyZx2R5cBVGlN
u5dndkHO6UlGR4IYp3xnbp2eNbgk1/+0QWSFSbz4L5t0lsrghEfWiPw1yvFmyO41
+cCRzVEuaEbmrfEb+1vtvCYEh20OQ4yzzfZNnD8TF1y0bofs0egCp2NjLavog54R
wNDMNLgxqWYnVWRPNuLMdP68UWNlzsYznbu7Mwk/3oNdQkMBvuMzTIuHokQjwmzP
giXprLAARRLBV+Y/LSGJsGQJe2KOOS1BASYIY2vmyeoyc2qhLXAhzxVLk8vNd+z8
LMBJ5x8V2LNI1dv6X2QJI4LTr/23YdDPOX/S1PPBDI35rtdpubF1RibIeh0IFaGQ
JdhuovR6Ld5zdj+Hir1Hnk7jl9/Kbb64a0UbEUegU76nvu5ol0R33BduufVE0LNd
ZESIMuS2jtszmLlUWPSt9xYM3AUD6e1aB3uBFSuk8IzleZ5H4+t8bBpwKDrL8zMI
WZSTmPT6H8UessmNZa8X/JodqlDXUqD9fbI5r+/88NlFMhe7T5yaxLt79iTthY47
u+yutIeT8rQSmBO+qV89mmL8SWAgIvofHqI/RDuIO6i8QsbUFZ3k2jhqIzHsBW0Y
Z/eFzp7iC2TuxIWfuX7BLb1QJ1CFCd2e4ZXQ/A2R/glrAtAV/g8anDNRjVoB7ibQ
UyoOtnvwZz84UbTvqJjOsEq5a7Id+wpvDt/nZzGZTLi2h4dqNRsZGSqtwtKjsvsx
iTzj9WMeqXhx7ML6zxVQw8SpgYficlFvLe0LnPaiRm6UjnaOpFpU+V2pLjZ1H7dy
JTlJPNhjrafp7wGDK55xfxdsVI2rFOntqAgyA8TRtKnLgNwwJvDfMo13a/AbGNK1
0LVKbxIDEzBd4hV8Bf8vhxAgU0NSBe4Eg4syPvDMu4E/rrbxlx45hk4QAGgsNrUJ
o94a5hs1a8KmJptwSGOkyzyddAKyY9Pl7PHFnI27FjODyGYJ171npLiGV/7yDdvl
WbznaMgCGLd0kSMnPF0LW4tpA2ciScgkYdpimCF+WJ2QYNAoNdiqZ+yby6TKoqGR
EbEbWHTJV96nFcaG/zIAu/mV7gPgKZGMssVPw3nDtGd7KsH6tJSfh6MP6teNQvHn
cI6C8Q0NU2biykglfXNu7UBL57EMvI+5SQvQB+60Z8ihj5Roh36BxgixGq/VPS41
KdsbADyXY3UFXICwTd83o9CiS2pb6RUpXs1nztZe0UG1OvZdRoYoG048lMTBN1aK
D8rbBDS/yFz6prhRQEFfxmsJAk5h4l6zkh9jVBujnpDSdkSMOs5k/aL9COKFGFnW
aVioJN/PgXT/N9Qrnv5FMtPUmIh1fN/0fFv4PACjKQ3F18AgpFZrFC3XQYihyND5
GL7JkiFSx2gcCgLFh43zGY0tUEjaPgwo+8YQRU7tIc3jJi3BLGoihHzVdzkTlnTo
ZXNX3md8XnSpxBmiGBykS3/ROFzou5G3fckRDcYSup/vHMUd/Mka3Zmy3cdw+3zB
fhVLKVPvP0Q/LfyuaXaMjk9GenyF34iJz0ykVThtMhf5JSfnQuC3/IqwwNOeBM1I
CiqaoqErnWC+TBdukOvP33tuHwlkhR0sG4EcOaMlBmNCR7EZdusYQ0cZWMQzNCzZ
cmXE+nlQKq0cMkedZ8nC7EBY5pr9s2xJ7zul6H/6cWXP8Qo8c2fNk/AHnpzEo4uR
J0V8jHu1CcL05Gh2wxvmTKv1i3qaYPz/0VKHlw8mqQFGLrG0I/YueHRF4k/XLANG
S8OUXey79AYcHmmKaA6YNTVcEabzYtv86dycqX7zwrjr4Uane3Z20NvUwAXrWsNy
ihEccjJXIP6/FtIh3Jg9WJ28fBHngA0EHZA/US4ykD+2orm+CYKBL5NK7yvV0p+S
F0IDWstTGKGRIS9C//lvPTe1iTxhTHGD/ImIvjURPpzaFFKjLBegm/rpo06YTW/4
T+9CpcM5gLrjVqS4SHdlDqVRwuhYjfuCGODakubxx5jemnRFguI7Ojaj0eia0mtQ
C7WqJRtik8+hRMTf3Ojm1+/EyiTvdL3OA/47Bm3Exmo/tww9D+XYtTYzmoMY/+lG
wVM5W+bqeUtkfz1oS1mWrlrkwoN2GllfXeH0LO3fFmbOEJh4wVrWQkbianeiAwOY
2OgYGtlqqARKU2cf5PGwGPO1iPf+iPaHiATGnzRjypzhodgxA6C1Vw6PCsT9PPAf
HOVWdD6VrMVYJjmbhG8R/+WT6bOVx+43akL+AGxzpXGyveJV76Bp2OyRg0m5B9QE
DONCN+Ojh1VWtcskkbLfofqtdHqrq6FltA9bLgGy/Ap3FqWYnOaCw4/B/gsSrqKu
F3DePtvHTkG346I7TMSFQJ9rPkRujGdV2ubHBTJ+iqJhLTF5RAO2ouzd71gAuRSH
VrU7S4nhq74gzVLJlGbeXsFWo96MU5mpDHIEsidFrvZtCsN1zIJvvorkjba1T9Ev
oSzDI+RIrEwevm6golv3zluLdgzCimFLaQBYCYTgJ+rv/H8WI3MujmxCPIidTGYr
FT1UxTIgtnquKe03pHOgX4G1FeHkk2M55Af0/fzoshD+ePOc/tEHnMM2oefenB3c
QM3G+u1YBDZb1pL9YmHNT4mIqgWq4lbeFAh0Vz6sPszOgumlIy3xAZESZh8GaCLc
ZXjjcqfoSaWuVewXiLLQnfUPc/Eh8y0ZL5O+ND+RlKazJXrUOFz+tdqm0Ts+SMW8
dSa3bOK5GelgpDSUfu/LZShw7gHzdduOAFgV9BwhqP9D8Sf+mqLYCpXl94giVNdK
rjmTTKoyMZpjyXse0kiXk7cDPAPvRLG3mEL2/Y/tB4P2c1NYT7XglsT2fHkPvbW2
hosCDrRDbySFrWpxVRQodvH8JLQ4YBiFho6LHIkAdo4XMSp807Xcl60f907Z9ei/
q0jLX9YVnI8NiEXSrPZmNxwxpGD7wTCnOMcdm746xNWvAHYb7dEDxUcRcRRdH9jE
c3lxTIl+fPJf4BxMHoB9TzPHhKgtEcumFkIFDfIHWZAkvjt/n0mgcb0oXxorbYkc
ishRfK2ivqDZHX17JKxdKXZezmhAt8M2FhJ8S+fXACZSujNKvynmjdQg8XqEZpQX
2NDWGdfTWFmPucBvgqc/g2TbwrmscDtUwxgeGiiJPayf9rvElAVNTWy/P16+72eV
/gfNIyzQUThuuxgMJ8ED+HPvRlfkFObmJkRmevbAwULZFs8jQYrlpbuyr9Dy2scw
0+nFcc/RSpKKjrctNDqg4Y8tAFXmbWeWzavA3IbigTfDJMGpQRYZyC/uAEKu7q1D
+8mX8hhJMSI+SfRnvkAPN6qCzXEIXCyQrnFw/JlD/XRzvv+lIszg3jTSDnmgUMnO
aScQR7HlLMQf72U8F/B9AYAXgJpQdJXQ4t8+qV2GkLJvntHnq5VLf7BLMSLxfNpW
AYDzrxRNKmQnCuzvHb8syRyRvmGmTKAORd3mmMOwi7faYZnw4MEziiYp1r89c1PR
owHQ8JRtmD4G1ZfIhlgWQ0WmBpNsE2Yhe7UwiK1JQY5PVPdiv3LOY6uR3Jk7ltJ4
Kl4hRYyFY2GluR6dx6zAFY1g9IBlg9gGRZjDqeBuanBsismN9iUfUyF1Wx7wys31
cHBAoxNzUepykhneff29NY8xsfH5shcaafufeIaUE4BLvlQNIG3XQv9LeamjII/x
4xdnYSuJJPIDvzOLihsk/MHlfHyklnYylNX9n06kS1/xW/f8Ef3ypomrr3KWonnS
Bi47C/PAPb4LIwW2eHO+lcHc1cidSKWAfmqbheRlHyDrZCqE0aOLKT8xWmmrQudo
z5sEyEiJJharphQXqz6uyGGleqo/9rLRqOyaGWrlJWzaTEN9o5NKGg+fwX6YTY3i
8gzlaMwOtA9fmuDAx9EIrs5VdOuyirB0clZeolTt6Pp+JRSKyt47387uAzQV3xRD
WUPZbT0b9W4EoSZp5JvjVkgIviXnx+MylOZ5HmpTdZwi5m5Ibzrs0sdJDyRRC/PG
JBHoSKk3hfWjV0j7IU2V8MXfgyJsxMSiNNz9YOc19Szxf9KxfURwjhtdo3uNULqU
1f9x5aB2qB9ntJeGai0QAsvqSMeT6q9D/N3Qh37j7KtO+RLPdvM2OkWmk9lu+Ed0
5OfkZFIyh46vVbT07B9N2DWqXlJVbaZn2VMKQfttWDsL/nc3K4P0JCVpCGwZyFHS
vXnSQ5incWsBdXZxibYSGBjVOEaBw8u3uDlnS1kljwh4JhipjBEyK2bY8mAzCf2b
BJ1CPQ3nq/4S33bvM/2EycVDqzUep/fcNMilmXC37s4rGWFOrJuiuYDAAg4/aFQ5
TP1bPdEgIYz/EmQTrF/vfr0TWVd1DHDR5GoUVyc5p7r6HTwZo/IEDSA8DqdyLQqH
gG3KTIIE909weqB3w6Ysj9HqyQC5gfCDND/e/7KxPE84Csou262iOwEzBHkR9Scm
dmThTLSRY0HsVQQ4YUAfrQC7BUZuWtU2jUmFA22lIqPHf3BR9BMx6Plk3aE6cZ5j
9zMsrUt5feK/FnK/DbN+RhpSDiZG9Rcz8bARGmuxluMLBR1DTirTp8BenX/ayAW0
It+GXxRfgsDJQdLPG5E3YqafUcaypym2pApEAnAMAjlHCco7aiKS5m/LvclRRqNC
GrnDmoH4CxEkrjp94L1/MdR9BpOx9BgH9kuDfoeae/V0CAXu9ukIuuhPjOwF81E4
yrRHgU9Jgb/bLa4nI1NCGLtb5PCLAxTgpFLu987EDiRJ0m0AX577tnz5y7SmCrR+
F05P++yptcgaFpe16IBoVOGXHW/hNhKdt2VRV+5XbVXu7Ycih2jZio3iQXoRmcAX
bb0aHhGVBtmSwaNd+2hmPHJmeBMz2M9AkZXFQla6sWHGbxaqs49ydd3iw2lW7DAJ
k+lKVah940nxLZFyrf4yU/uEZLSp91SHwwlZyzuC36qDCA64EyXLJWr8pJyO1yTt
R8+FRv90c92fVzdD3BPaIiqBS1a3HOcENp5s4uEJmmLjcmSKD6KuGMDQTx3Mkfa2
ijUyWbkvoAiwLvuD4U/weNRB2Y+ZcvVFrpYnQ/lGA7GQOIHPMTcWpqceVsKfbKZp
8+vdB5YnQr1fK836T1Uz7HNhht4CQ8x0VJotjjbChKc+SPOl0pFzfLvjPLw9lSSM
a6daz0ywbcDVgHsbHlvpSkw3w/XLPZuibqK2nRERdazPdL6IAIIV5Q5mppegr45i
SobKapcORVSTfFCcBU9VqDF3d8Sm64fQVkIGVNL7awN5Qd7nQcNlfMxvNCZsR4RN
SqSJViL8xnjLcIi6WTv9YwtHvgHywbm5bpdAeLTOjgS95b4QkI6WWU+DluNRxxwC
6DqE4ujfCdstJ8ZK0Bws6y991BQ3Ebo3uMHLgqQRn4GM0mRTlPJkfAp48NCpWnBY
37Bla2iFPD/1kb54hdHz9Z7ae3CBvS3cgREcLePnStEKx87zU1zFDaf6aQ4RnRdB
/uVTlrhje/IjXKZYH2qZ+6GZlq/dX7xgmGRSLUZXjG7rWUqBZOFM4jYa0uU8OlCA
/SaYszXRuLPg+20dCbtVNoANiUTkSoCtKT+MpXXZYuBraHlUu/pU9BdXQdmV7AJb
HBsVdMMfI23HQbf4uu4D71OIfR0Kr48ayapzU3zcZYrbqP0lxAYI+Gobill+kXtI
xReuFAI6abzt+aFLIyEY7lM/VtUuY0GBHSL9KK43BkO1vlarbCQabWqW4+H8sO30
Oe638otOPn14pSRp/ER45bfYnwGvt3oGHbKQKv+i1gru9pBAHNa/mtWN0j4sDybk
h+mbVmEDCFodBq937dFmQNYzbjOcxa4xT0Ali0m2HS7NSgMhSHmKV5d4sqNulSz/
ffUge6HdyvLOKciEj8Q+DQp5Ez3JbsAblCsq5fUH1/udZE9cqsXa2G1qmIFxqh2I
0d/CC3/Ak19ZK5cDWQ1/iUy+oeK2z/xCelv1YIYEwRK90JLyBFvRk/bvVvIjyugx
Hkn6p9pdEUF55B9+IMt64ItH6ytns4l+s03fwVh1l5XBfEN8VPOGqsq0s9AzZdSs
s/DluDb6/SoEA8Pimjl6vDuEB0kfMqcF6qCGRT/kJUVMeDljBqurUyol8weRI7j0
T1FsBC7yl94OLmgAff+NnO6Mi9Al97GUub4xABDfhleEN3Ze8KAoVG78k8UGkw8w
OF06Z1KDr18UPFr7deSMuYqL42Z4yIVwoV3BqvH8RBIl6abwCfieJxCH/cebVXMW
SXhK/gVIu8FlTVIkfeUBR1+Eqon00IJlYofXUUIYhjuJn0Nzj5G5Uyb1aH8AT0Fl
CG3AMiQpVT5GYW5CbW3qxoe31IB+V6XfRq5dQYU5ilGTuXj01XM7M+mk8MdtxVZL
2npGvAqaz/WymHhF4EQOq1TyTcHuGeXf5Hplbjh71vWKXWH74TiI0vcOq97utPqS
xwGjmS/C7dzhDmmymBMFzQZnt3Cq4wg1yxfxEBbWuxttT3eMLdt3Jt1m7FCt3vU2
gnqO10Z7vRFL7dffFZARhfD7SpbuVBoVycuzbPB/RUpqdi85Lbl7dTpVTXbLHp+W
ddR6b9T4Ieix7hPZ2y+/mHWJ+nB18jCx+mBrAhnjTjO1r6OGiRi0SCmqSseBUqQk
`pragma protect end_protected
